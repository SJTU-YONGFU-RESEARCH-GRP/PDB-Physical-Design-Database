module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire net17762;
 wire net17731;
 wire net17735;
 wire net17737;
 wire net17732;
 wire net17777;
 wire net17792;
 wire net17793;
 wire net17727;
 wire _00394_;
 wire net17726;
 wire net17761;
 wire net17723;
 wire net17729;
 wire _00399_;
 wire net17794;
 wire net17758;
 wire net17739;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00910_;
 wire _00911_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00981_;
 wire _00984_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01083_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01665_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01687_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01727_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01733_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01783_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01793_;
 wire _01794_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02386_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02406_;
 wire _02407_;
 wire _02409_;
 wire _02410_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02442_;
 wire _02443_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02484_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire net258;
 wire _02492_;
 wire _02493_;
 wire net257;
 wire _02495_;
 wire _02496_;
 wire net256;
 wire net255;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire net254;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire net253;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire net252;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire net251;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire net250;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire net249;
 wire net248;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire net247;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire net246;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire net245;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire net243;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire net241;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire net240;
 wire _03145_;
 wire net239;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire net238;
 wire net237;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire net236;
 wire _03165_;
 wire _03166_;
 wire net235;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire net234;
 wire net233;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire net232;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire net231;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire net230;
 wire _03203_;
 wire _03204_;
 wire net229;
 wire _03206_;
 wire net228;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire net227;
 wire net226;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire net225;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire net224;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire net223;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire net222;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire net221;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire net220;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire net219;
 wire _03279_;
 wire net218;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire net217;
 wire _03290_;
 wire _03291_;
 wire net216;
 wire _03293_;
 wire _03294_;
 wire net215;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire net214;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire net213;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire net212;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire net211;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire net210;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire net209;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire net208;
 wire net207;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire net204;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire net203;
 wire net202;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire net201;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire net200;
 wire net199;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire net198;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire net197;
 wire _03928_;
 wire _03929_;
 wire net196;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire net195;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire net194;
 wire net193;
 wire net192;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire net191;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire net190;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire net189;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire net188;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire net187;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire net186;
 wire _04001_;
 wire net185;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire net184;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire net183;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire net182;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire net181;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire net180;
 wire _04033_;
 wire _04034_;
 wire net179;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire net178;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire net177;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire net176;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire net175;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire net174;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire net173;
 wire _04153_;
 wire _04154_;
 wire net172;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire net171;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire net167;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire net166;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire net165;
 wire net164;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire net163;
 wire _04622_;
 wire net162;
 wire net161;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire net160;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire net159;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire net158;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire net157;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire net156;
 wire _04676_;
 wire net155;
 wire net154;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire net153;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire net152;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire net151;
 wire _04721_;
 wire net150;
 wire _04723_;
 wire _04724_;
 wire net149;
 wire _04726_;
 wire net148;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire net147;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire net146;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire net145;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire net144;
 wire _04759_;
 wire _04760_;
 wire net143;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire net142;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire net141;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire net140;
 wire _04808_;
 wire net139;
 wire _04810_;
 wire _04811_;
 wire net138;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire net137;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire net136;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire net135;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire net134;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire net133;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire net131;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire net129;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire net128;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire net127;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire net126;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire net125;
 wire net124;
 wire _05370_;
 wire _05371_;
 wire net123;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire net122;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire net121;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire net120;
 wire net119;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire net118;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire net117;
 wire _05410_;
 wire net116;
 wire net115;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire net114;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire net113;
 wire _05447_;
 wire net112;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire net111;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire net110;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire net109;
 wire _05474_;
 wire _05475_;
 wire net108;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire net107;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire net106;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire net105;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire net104;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire net103;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire net102;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire net101;
 wire _05543_;
 wire _05544_;
 wire net100;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire net99;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire net98;
 wire _05563_;
 wire net97;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire net96;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire net95;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire net93;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire net91;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire net89;
 wire net88;
 wire _06074_;
 wire _06075_;
 wire net87;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire net86;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire net85;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire net84;
 wire net83;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire net82;
 wire _06111_;
 wire net81;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire net80;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire net79;
 wire _06125_;
 wire _06126_;
 wire net78;
 wire _06128_;
 wire _06129_;
 wire net77;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire net76;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire net75;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire net74;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire net73;
 wire _06182_;
 wire net72;
 wire _06184_;
 wire net71;
 wire _06186_;
 wire _06187_;
 wire net70;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire net69;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire net68;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire net67;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire net66;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire net65;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire net64;
 wire _06238_;
 wire _06239_;
 wire net63;
 wire _06241_;
 wire _06242_;
 wire net62;
 wire _06244_;
 wire net61;
 wire _06246_;
 wire net60;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire net59;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire net58;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire net57;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire net56;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire net55;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire net54;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire net50;
 wire _06784_;
 wire net49;
 wire _06786_;
 wire _06787_;
 wire net48;
 wire net47;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire net46;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire net45;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire net44;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire net43;
 wire net42;
 wire _06842_;
 wire net41;
 wire _06844_;
 wire _06845_;
 wire net40;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire net39;
 wire _06851_;
 wire _06852_;
 wire net38;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire net37;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire net36;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire net35;
 wire _06881_;
 wire net34;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire net33;
 wire net32;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire net31;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire net30;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire net29;
 wire net28;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire net27;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire net26;
 wire net25;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire net24;
 wire _06931_;
 wire net23;
 wire _06933_;
 wire _06934_;
 wire net22;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire net21;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire net20;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire net19;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire net18;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire net17;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire net16;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire net15;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire net14;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire net13;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire net17768;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire net17800;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire net17769;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire net17803;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire net17775;
 wire net17785;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire net12;
 wire _07475_;
 wire net11;
 wire _07477_;
 wire net10;
 wire _07479_;
 wire net9;
 wire _07481_;
 wire _07482_;
 wire net8;
 wire _07484_;
 wire net7;
 wire net17790;
 wire net6;
 wire net5;
 wire _07489_;
 wire net4;
 wire _07491_;
 wire net3;
 wire _07493_;
 wire net2;
 wire _07495_;
 wire net1;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire net17748;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire net17751;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire net17744;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire net17747;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire net17757;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire net17754;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire net17734;
 wire _07639_;
 wire net17733;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire net17721;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire net17717;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire net17730;
 wire net17759;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire net17760;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire net17749;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire net17716;
 wire net17718;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire net17741;
 wire _07784_;
 wire _07785_;
 wire net17714;
 wire _07787_;
 wire _07788_;
 wire net17740;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire net17724;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire net17725;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire net17706;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire net17713;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire net17719;
 wire _07941_;
 wire net17703;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire net17702;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire net17704;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire net17709;
 wire net17710;
 wire _07987_;
 wire _07988_;
 wire net17707;
 wire _07990_;
 wire net17693;
 wire net17697;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire net17746;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire net17700;
 wire net17701;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire net17690;
 wire net17689;
 wire _08019_;
 wire _08020_;
 wire net17818;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire net17686;
 wire _08029_;
 wire _08030_;
 wire net17711;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire net17684;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire net17683;
 wire _08048_;
 wire net17682;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire net17681;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire net17685;
 wire _08070_;
 wire _08071_;
 wire net17679;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire net17691;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire net17743;
 wire _08081_;
 wire net17687;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire net17675;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire net17674;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire net17669;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire net17666;
 wire net17673;
 wire _08126_;
 wire net17665;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire net17664;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire net17667;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire net17672;
 wire net17680;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire net17661;
 wire _08581_;
 wire _08582_;
 wire net17670;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire net17668;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire net17660;
 wire net17676;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire net17656;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire net17663;
 wire net17677;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire net17708;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire net17650;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire net17648;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire net17820;
 wire _08650_;
 wire net17822;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire net17649;
 wire net17821;
 wire _08658_;
 wire net17643;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire net17642;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire net17671;
 wire _08669_;
 wire _08670_;
 wire net17819;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire net17653;
 wire _08694_;
 wire _08695_;
 wire net17644;
 wire _08697_;
 wire net17637;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire net17635;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire net17658;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire net17627;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire net17628;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire net17626;
 wire _09155_;
 wire _09156_;
 wire net17659;
 wire net17622;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire net17620;
 wire _09164_;
 wire _09165_;
 wire net17619;
 wire net17618;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire net17617;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire net17824;
 wire net17623;
 wire _09185_;
 wire _09186_;
 wire net17614;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire net17657;
 wire _09206_;
 wire net17613;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire net17624;
 wire _09212_;
 wire _09213_;
 wire net17610;
 wire _09215_;
 wire _09216_;
 wire net17621;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire net17611;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire net17612;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire net18241;
 wire _09236_;
 wire net17606;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire net18242;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire net17605;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire net17604;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire net17607;
 wire _09282_;
 wire net17678;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire net17609;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire net17600;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire net17756;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire net17601;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire net17603;
 wire _09749_;
 wire net17593;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire net17599;
 wire _09757_;
 wire _09758_;
 wire net17602;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire net17825;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire net17592;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire net17596;
 wire _09774_;
 wire _09775_;
 wire net17597;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire net17585;
 wire net17590;
 wire _09788_;
 wire net17584;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire net17582;
 wire _09796_;
 wire net17580;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire net17579;
 wire _09808_;
 wire _09809_;
 wire net17578;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire net17577;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire net17581;
 wire _09830_;
 wire _09831_;
 wire net17575;
 wire _09833_;
 wire net17574;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire net17583;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire net17576;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire net17586;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire net17591;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire net17567;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire net17568;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire net17572;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire net17573;
 wire _09939_;
 wire net17616;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire net17589;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire net17564;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire net17561;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire net17608;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire net17588;
 wire _10380_;
 wire net17559;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire net17565;
 wire net17625;
 wire _10404_;
 wire net17552;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire net17560;
 wire net17555;
 wire net17548;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire net17546;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire net17823;
 wire _10480_;
 wire _10481_;
 wire net17570;
 wire net17539;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire net17536;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire net17571;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire net17598;
 wire net17920;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire net17535;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire net17534;
 wire net17857;
 wire _10524_;
 wire net17849;
 wire net17531;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire net17848;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire net17529;
 wire _10539_;
 wire net17846;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire net17844;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire net17527;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire net17530;
 wire _10565_;
 wire net17528;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire net17525;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire net17830;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire net17832;
 wire net17522;
 wire net17521;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire net18392;
 wire _10592_;
 wire net18535;
 wire net17523;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire net17520;
 wire _10601_;
 wire _10602_;
 wire net18518;
 wire _10604_;
 wire net17524;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire net17532;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire net17519;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire net17517;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire net17508;
 wire _10633_;
 wire net17505;
 wire net17509;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire net17515;
 wire _10640_;
 wire _10641_;
 wire net17540;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire net17492;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire net17545;
 wire _10660_;
 wire net17497;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire net17488;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire net17489;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire net17490;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire net17544;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire net17484;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire net17547;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire net17491;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire net17483;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire net17538;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire net17516;
 wire net17526;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire net17493;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire net17485;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire net17482;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire net17512;
 wire net17533;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire net17475;
 wire net17469;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire net17468;
 wire _11326_;
 wire _11327_;
 wire net17465;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire net17473;
 wire net17464;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire net17463;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire net17470;
 wire net17457;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire net17460;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire net17467;
 wire _11373_;
 wire net17459;
 wire _11375_;
 wire _11376_;
 wire net17518;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire net18536;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire net17453;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire net17451;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire net17445;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire net18278;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire net18252;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire net18388;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire net18378;
 wire _11434_;
 wire _11435_;
 wire net18729;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire net17449;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire net18633;
 wire net17443;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire net18615;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire net17456;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire net17450;
 wire _11525_;
 wire net17441;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire net17446;
 wire _11599_;
 wire net18614;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire net17448;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire net18613;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire net18728;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire net17434;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire net17430;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire net17436;
 wire net17424;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire net18611;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire net18588;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire net17417;
 wire net17415;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire net17418;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire net18610;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire net17413;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire net17411;
 wire net18695;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire net17421;
 wire _12174_;
 wire net17416;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire net17412;
 wire net17405;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire net17402;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire net17400;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire net17404;
 wire _12198_;
 wire net17454;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire net17395;
 wire net17406;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire net17422;
 wire net17392;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire net17399;
 wire net17389;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire net17397;
 wire _12243_;
 wire net17391;
 wire _12245_;
 wire net17386;
 wire _12247_;
 wire net17387;
 wire _12249_;
 wire net17382;
 wire net17380;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire net17379;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire net17383;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire net17375;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire net17396;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire net17388;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire net17370;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire net17398;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire net18700;
 wire net17378;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire net17371;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire net17542;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire net17366;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire net17361;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire net17374;
 wire net17372;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire net17358;
 wire net17377;
 wire _12946_;
 wire _12947_;
 wire net17385;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire net17356;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire net17384;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire net17373;
 wire net19076;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire net17354;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire net17351;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire net17348;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire net17353;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire net17349;
 wire net17347;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire net17381;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire net17355;
 wire _13038_;
 wire net17390;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire net17345;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire net17340;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire net17344;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire net17339;
 wire _13065_;
 wire _13066_;
 wire net17335;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire net17401;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire net17346;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire net17330;
 wire _13108_;
 wire _13109_;
 wire net17350;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire net17338;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire net17332;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire net17472;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire net17471;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire net17317;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire net17342;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire net17341;
 wire _13172_;
 wire net17352;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire net17343;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire net17329;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire net17306;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire net17312;
 wire net17308;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire net17307;
 wire net17300;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire net17299;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire net17311;
 wire net17309;
 wire _13724_;
 wire _13725_;
 wire net17296;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire net17303;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire net17301;
 wire net17290;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire net17291;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire net17305;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire net17292;
 wire _13770_;
 wire net17282;
 wire net17288;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire net17284;
 wire net17277;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire net17315;
 wire _13792_;
 wire _13793_;
 wire net17283;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire net19063;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire net19267;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire net19332;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire net17266;
 wire _13866_;
 wire _13867_;
 wire net19306;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire net17270;
 wire net17264;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire net17262;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire net17261;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire net17285;
 wire _13897_;
 wire _13898_;
 wire net17259;
 wire _13900_;
 wire net19305;
 wire net19177;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire net19282;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire net19513;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire net20459;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire net17248;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire net17246;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire net17250;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire net17253;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire net19450;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire net19492;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire net17236;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire net17238;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire net19491;
 wire _14485_;
 wire net17235;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire net17237;
 wire _14495_;
 wire _14496_;
 wire net17234;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire net17232;
 wire _14505_;
 wire net17233;
 wire _14507_;
 wire net17244;
 wire net17242;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire net17252;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire net17230;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire net19462;
 wire _14527_;
 wire net17228;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire net17227;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire net17255;
 wire _14538_;
 wire _14539_;
 wire net17229;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire net19456;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire net17239;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire net17219;
 wire _14573_;
 wire net19455;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire net19461;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire net17215;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire net17220;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire net17216;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire net20436;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire net19849;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire net20629;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire net20737;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire net20696;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire net17203;
 wire net17206;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire net20761;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire net17287;
 wire net17201;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire net17276;
 wire _15198_;
 wire net20913;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15213_;
 wire _15216_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15224_;
 wire _15225_;
 wire _15227_;
 wire _15228_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15260_;
 wire _15261_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15279_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15348_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire net17695;
 wire net17755;
 wire net17662;
 wire net17736;
 wire net17655;
 wire net17745;
 wire net17594;
 wire net17808;
 wire net17595;
 wire net17629;
 wire net17502;
 wire net17496;
 wire net17479;
 wire net17431;
 wire net18612;
 wire net17428;
 wire net17359;
 wire net17369;
 wire net17304;
 wire net17461;
 wire net17241;
 wire net17243;
 wire net20762;
 wire net17205;
 wire net242;
 wire net244;
 wire net205;
 wire net206;
 wire net169;
 wire net168;
 wire net170;
 wire net130;
 wire net132;
 wire net94;
 wire net90;
 wire net92;
 wire net53;
 wire net51;
 wire net52;
 wire \dcnt[0] ;
 wire \dcnt[1] ;
 wire \dcnt[2] ;
 wire \dcnt[3] ;
 wire net259;
 wire ld_r;
 wire \sa00_sr[0] ;
 wire \sa00_sr[1] ;
 wire \sa00_sr[2] ;
 wire \sa00_sr[3] ;
 wire \sa00_sr[4] ;
 wire \sa00_sr[5] ;
 wire \sa00_sr[6] ;
 wire \sa00_sr[7] ;
 wire \sa01_sr[0] ;
 wire \sa01_sr[1] ;
 wire \sa01_sr[2] ;
 wire \sa01_sr[3] ;
 wire \sa01_sr[4] ;
 wire \sa01_sr[5] ;
 wire \sa01_sr[6] ;
 wire \sa01_sr[7] ;
 wire \sa02_sr[0] ;
 wire \sa02_sr[1] ;
 wire \sa02_sr[2] ;
 wire \sa02_sr[3] ;
 wire \sa02_sr[4] ;
 wire \sa02_sr[5] ;
 wire \sa02_sr[6] ;
 wire \sa02_sr[7] ;
 wire \sa03_sr[0] ;
 wire \sa03_sr[1] ;
 wire \sa03_sr[2] ;
 wire \sa03_sr[3] ;
 wire \sa03_sr[4] ;
 wire \sa03_sr[5] ;
 wire \sa03_sr[6] ;
 wire \sa03_sr[7] ;
 wire \sa10_sr[0] ;
 wire \sa10_sr[1] ;
 wire \sa10_sr[2] ;
 wire \sa10_sr[3] ;
 wire \sa10_sr[4] ;
 wire \sa10_sr[5] ;
 wire \sa10_sr[6] ;
 wire \sa10_sr[7] ;
 wire \sa10_sub[0] ;
 wire \sa10_sub[1] ;
 wire \sa10_sub[2] ;
 wire \sa10_sub[3] ;
 wire \sa10_sub[4] ;
 wire \sa10_sub[5] ;
 wire \sa10_sub[6] ;
 wire \sa10_sub[7] ;
 wire \sa11_sr[0] ;
 wire \sa11_sr[1] ;
 wire \sa11_sr[2] ;
 wire \sa11_sr[3] ;
 wire \sa11_sr[4] ;
 wire \sa11_sr[5] ;
 wire \sa11_sr[6] ;
 wire \sa11_sr[7] ;
 wire \sa12_sr[0] ;
 wire \sa12_sr[1] ;
 wire \sa12_sr[2] ;
 wire \sa12_sr[3] ;
 wire \sa12_sr[4] ;
 wire \sa12_sr[5] ;
 wire \sa12_sr[6] ;
 wire \sa12_sr[7] ;
 wire \sa20_sr[0] ;
 wire \sa20_sr[1] ;
 wire \sa20_sr[2] ;
 wire \sa20_sr[3] ;
 wire \sa20_sr[4] ;
 wire \sa20_sr[5] ;
 wire \sa20_sr[6] ;
 wire \sa20_sr[7] ;
 wire \sa20_sub[0] ;
 wire \sa20_sub[1] ;
 wire \sa20_sub[2] ;
 wire \sa20_sub[3] ;
 wire \sa20_sub[4] ;
 wire \sa20_sub[5] ;
 wire \sa20_sub[6] ;
 wire \sa20_sub[7] ;
 wire \sa21_sr[0] ;
 wire \sa21_sr[1] ;
 wire \sa21_sr[2] ;
 wire \sa21_sr[3] ;
 wire \sa21_sr[4] ;
 wire \sa21_sr[5] ;
 wire \sa21_sr[6] ;
 wire \sa21_sr[7] ;
 wire \sa21_sub[0] ;
 wire \sa21_sub[1] ;
 wire \sa21_sub[2] ;
 wire \sa21_sub[3] ;
 wire \sa21_sub[4] ;
 wire \sa21_sub[5] ;
 wire \sa21_sub[6] ;
 wire \sa21_sub[7] ;
 wire \sa30_sr[0] ;
 wire \sa30_sr[1] ;
 wire \sa30_sr[2] ;
 wire \sa30_sr[3] ;
 wire \sa30_sr[4] ;
 wire \sa30_sr[5] ;
 wire \sa30_sr[6] ;
 wire \sa30_sr[7] ;
 wire \sa30_sub[0] ;
 wire \sa30_sub[1] ;
 wire \sa30_sub[2] ;
 wire \sa30_sub[3] ;
 wire \sa30_sub[4] ;
 wire \sa30_sub[5] ;
 wire \sa30_sub[6] ;
 wire \sa30_sub[7] ;
 wire \sa31_sub[0] ;
 wire \sa31_sub[1] ;
 wire \sa31_sub[2] ;
 wire \sa31_sub[3] ;
 wire \sa31_sub[4] ;
 wire \sa31_sub[5] ;
 wire \sa31_sub[6] ;
 wire \sa31_sub[7] ;
 wire \sa32_sub[0] ;
 wire \sa32_sub[1] ;
 wire \sa32_sub[2] ;
 wire \sa32_sub[3] ;
 wire \sa32_sub[4] ;
 wire \sa32_sub[5] ;
 wire \sa32_sub[6] ;
 wire \sa32_sub[7] ;
 wire \text_in_r[0] ;
 wire \text_in_r[100] ;
 wire \text_in_r[101] ;
 wire \text_in_r[102] ;
 wire \text_in_r[103] ;
 wire \text_in_r[104] ;
 wire \text_in_r[105] ;
 wire \text_in_r[106] ;
 wire \text_in_r[107] ;
 wire \text_in_r[108] ;
 wire \text_in_r[109] ;
 wire \text_in_r[10] ;
 wire \text_in_r[110] ;
 wire \text_in_r[111] ;
 wire \text_in_r[112] ;
 wire \text_in_r[113] ;
 wire \text_in_r[114] ;
 wire \text_in_r[115] ;
 wire \text_in_r[116] ;
 wire \text_in_r[117] ;
 wire \text_in_r[118] ;
 wire \text_in_r[119] ;
 wire \text_in_r[11] ;
 wire \text_in_r[120] ;
 wire \text_in_r[121] ;
 wire \text_in_r[122] ;
 wire \text_in_r[123] ;
 wire \text_in_r[124] ;
 wire \text_in_r[125] ;
 wire \text_in_r[126] ;
 wire \text_in_r[127] ;
 wire \text_in_r[12] ;
 wire \text_in_r[13] ;
 wire \text_in_r[14] ;
 wire \text_in_r[15] ;
 wire \text_in_r[16] ;
 wire \text_in_r[17] ;
 wire \text_in_r[18] ;
 wire \text_in_r[19] ;
 wire \text_in_r[1] ;
 wire \text_in_r[20] ;
 wire \text_in_r[21] ;
 wire \text_in_r[22] ;
 wire \text_in_r[23] ;
 wire \text_in_r[24] ;
 wire \text_in_r[25] ;
 wire \text_in_r[26] ;
 wire \text_in_r[27] ;
 wire \text_in_r[28] ;
 wire \text_in_r[29] ;
 wire \text_in_r[2] ;
 wire \text_in_r[30] ;
 wire \text_in_r[31] ;
 wire \text_in_r[32] ;
 wire \text_in_r[33] ;
 wire \text_in_r[34] ;
 wire \text_in_r[35] ;
 wire \text_in_r[36] ;
 wire \text_in_r[37] ;
 wire \text_in_r[38] ;
 wire \text_in_r[39] ;
 wire \text_in_r[3] ;
 wire \text_in_r[40] ;
 wire \text_in_r[41] ;
 wire \text_in_r[42] ;
 wire \text_in_r[43] ;
 wire \text_in_r[44] ;
 wire \text_in_r[45] ;
 wire \text_in_r[46] ;
 wire \text_in_r[47] ;
 wire \text_in_r[48] ;
 wire \text_in_r[49] ;
 wire \text_in_r[4] ;
 wire \text_in_r[50] ;
 wire \text_in_r[51] ;
 wire \text_in_r[52] ;
 wire \text_in_r[53] ;
 wire \text_in_r[54] ;
 wire \text_in_r[55] ;
 wire \text_in_r[56] ;
 wire \text_in_r[57] ;
 wire \text_in_r[58] ;
 wire \text_in_r[59] ;
 wire \text_in_r[5] ;
 wire \text_in_r[60] ;
 wire \text_in_r[61] ;
 wire \text_in_r[62] ;
 wire \text_in_r[63] ;
 wire \text_in_r[64] ;
 wire \text_in_r[65] ;
 wire \text_in_r[66] ;
 wire \text_in_r[67] ;
 wire \text_in_r[68] ;
 wire \text_in_r[69] ;
 wire \text_in_r[6] ;
 wire \text_in_r[70] ;
 wire \text_in_r[71] ;
 wire \text_in_r[72] ;
 wire \text_in_r[73] ;
 wire \text_in_r[74] ;
 wire \text_in_r[75] ;
 wire \text_in_r[76] ;
 wire \text_in_r[77] ;
 wire \text_in_r[78] ;
 wire \text_in_r[79] ;
 wire \text_in_r[7] ;
 wire \text_in_r[80] ;
 wire \text_in_r[81] ;
 wire \text_in_r[82] ;
 wire \text_in_r[83] ;
 wire \text_in_r[84] ;
 wire \text_in_r[85] ;
 wire \text_in_r[86] ;
 wire \text_in_r[87] ;
 wire \text_in_r[88] ;
 wire \text_in_r[89] ;
 wire \text_in_r[8] ;
 wire \text_in_r[90] ;
 wire \text_in_r[91] ;
 wire \text_in_r[92] ;
 wire \text_in_r[93] ;
 wire \text_in_r[94] ;
 wire \text_in_r[95] ;
 wire \text_in_r[96] ;
 wire \text_in_r[97] ;
 wire \text_in_r[98] ;
 wire \text_in_r[99] ;
 wire \text_in_r[9] ;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire \u0.r0.out[24] ;
 wire \u0.r0.out[25] ;
 wire \u0.r0.out[26] ;
 wire \u0.r0.out[27] ;
 wire \u0.r0.out[28] ;
 wire \u0.r0.out[29] ;
 wire \u0.r0.out[30] ;
 wire \u0.r0.out[31] ;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt[2] ;
 wire \u0.r0.rcnt[3] ;
 wire \u0.r0.rcnt_next[0] ;
 wire \u0.r0.rcnt_next[1] ;
 wire \u0.subword[0] ;
 wire \u0.subword[10] ;
 wire \u0.subword[11] ;
 wire \u0.subword[12] ;
 wire \u0.subword[13] ;
 wire \u0.subword[14] ;
 wire \u0.subword[15] ;
 wire \u0.subword[16] ;
 wire \u0.subword[17] ;
 wire \u0.subword[18] ;
 wire \u0.subword[19] ;
 wire \u0.subword[1] ;
 wire \u0.subword[20] ;
 wire \u0.subword[21] ;
 wire \u0.subword[22] ;
 wire \u0.subword[23] ;
 wire \u0.subword[24] ;
 wire \u0.subword[25] ;
 wire \u0.subword[26] ;
 wire \u0.subword[27] ;
 wire \u0.subword[28] ;
 wire \u0.subword[29] ;
 wire \u0.subword[2] ;
 wire \u0.subword[30] ;
 wire \u0.subword[31] ;
 wire \u0.subword[3] ;
 wire \u0.subword[4] ;
 wire \u0.subword[5] ;
 wire \u0.subword[6] ;
 wire \u0.subword[7] ;
 wire \u0.subword[8] ;
 wire \u0.subword[9] ;
 wire \u0.tmp_w[0] ;
 wire \u0.tmp_w[10] ;
 wire \u0.tmp_w[11] ;
 wire \u0.tmp_w[12] ;
 wire \u0.tmp_w[13] ;
 wire \u0.tmp_w[14] ;
 wire \u0.tmp_w[15] ;
 wire \u0.tmp_w[16] ;
 wire \u0.tmp_w[17] ;
 wire \u0.tmp_w[18] ;
 wire \u0.tmp_w[19] ;
 wire \u0.tmp_w[1] ;
 wire \u0.tmp_w[20] ;
 wire \u0.tmp_w[21] ;
 wire \u0.tmp_w[22] ;
 wire \u0.tmp_w[23] ;
 wire \u0.tmp_w[24] ;
 wire \u0.tmp_w[25] ;
 wire \u0.tmp_w[26] ;
 wire \u0.tmp_w[27] ;
 wire \u0.tmp_w[28] ;
 wire \u0.tmp_w[29] ;
 wire \u0.tmp_w[2] ;
 wire \u0.tmp_w[30] ;
 wire \u0.tmp_w[31] ;
 wire \u0.tmp_w[3] ;
 wire \u0.tmp_w[4] ;
 wire \u0.tmp_w[5] ;
 wire \u0.tmp_w[6] ;
 wire \u0.tmp_w[7] ;
 wire \u0.tmp_w[8] ;
 wire \u0.tmp_w[9] ;
 wire \u0.w[0][0] ;
 wire \u0.w[0][10] ;
 wire \u0.w[0][11] ;
 wire \u0.w[0][12] ;
 wire \u0.w[0][13] ;
 wire \u0.w[0][14] ;
 wire \u0.w[0][15] ;
 wire \u0.w[0][16] ;
 wire \u0.w[0][17] ;
 wire \u0.w[0][18] ;
 wire \u0.w[0][19] ;
 wire \u0.w[0][1] ;
 wire \u0.w[0][20] ;
 wire \u0.w[0][21] ;
 wire \u0.w[0][22] ;
 wire \u0.w[0][23] ;
 wire \u0.w[0][24] ;
 wire \u0.w[0][25] ;
 wire \u0.w[0][26] ;
 wire \u0.w[0][27] ;
 wire \u0.w[0][28] ;
 wire \u0.w[0][29] ;
 wire \u0.w[0][2] ;
 wire \u0.w[0][30] ;
 wire \u0.w[0][31] ;
 wire \u0.w[0][3] ;
 wire \u0.w[0][4] ;
 wire \u0.w[0][5] ;
 wire \u0.w[0][6] ;
 wire \u0.w[0][7] ;
 wire \u0.w[0][8] ;
 wire \u0.w[0][9] ;
 wire \u0.w[1][0] ;
 wire \u0.w[1][10] ;
 wire \u0.w[1][11] ;
 wire \u0.w[1][12] ;
 wire \u0.w[1][13] ;
 wire \u0.w[1][14] ;
 wire \u0.w[1][15] ;
 wire \u0.w[1][16] ;
 wire \u0.w[1][17] ;
 wire \u0.w[1][18] ;
 wire \u0.w[1][19] ;
 wire \u0.w[1][1] ;
 wire \u0.w[1][20] ;
 wire \u0.w[1][21] ;
 wire \u0.w[1][22] ;
 wire \u0.w[1][23] ;
 wire \u0.w[1][24] ;
 wire \u0.w[1][25] ;
 wire \u0.w[1][26] ;
 wire \u0.w[1][27] ;
 wire \u0.w[1][28] ;
 wire \u0.w[1][29] ;
 wire \u0.w[1][2] ;
 wire \u0.w[1][30] ;
 wire \u0.w[1][31] ;
 wire \u0.w[1][3] ;
 wire \u0.w[1][4] ;
 wire \u0.w[1][5] ;
 wire \u0.w[1][6] ;
 wire \u0.w[1][7] ;
 wire \u0.w[1][8] ;
 wire \u0.w[1][9] ;
 wire \u0.w[2][0] ;
 wire \u0.w[2][10] ;
 wire \u0.w[2][11] ;
 wire \u0.w[2][12] ;
 wire \u0.w[2][13] ;
 wire \u0.w[2][14] ;
 wire \u0.w[2][15] ;
 wire \u0.w[2][16] ;
 wire \u0.w[2][17] ;
 wire \u0.w[2][18] ;
 wire \u0.w[2][19] ;
 wire \u0.w[2][1] ;
 wire \u0.w[2][20] ;
 wire \u0.w[2][21] ;
 wire \u0.w[2][22] ;
 wire \u0.w[2][23] ;
 wire \u0.w[2][24] ;
 wire \u0.w[2][25] ;
 wire \u0.w[2][26] ;
 wire \u0.w[2][27] ;
 wire \u0.w[2][28] ;
 wire \u0.w[2][29] ;
 wire \u0.w[2][2] ;
 wire \u0.w[2][30] ;
 wire \u0.w[2][31] ;
 wire \u0.w[2][3] ;
 wire \u0.w[2][4] ;
 wire \u0.w[2][5] ;
 wire \u0.w[2][6] ;
 wire \u0.w[2][7] ;
 wire \u0.w[2][8] ;
 wire \u0.w[2][9] ;
 wire net17799;
 wire net17802;
 wire net17774;
 wire net17765;
 wire net17772;
 wire net17767;
 wire net17773;
 wire net17778;
 wire net17770;
 wire net17771;
 wire net17784;
 wire net17776;
 wire net17858;
 wire net17780;
 wire net17850;
 wire net18014;
 wire net17814;
 wire net17781;
 wire net17789;
 wire net17782;
 wire net18240;
 wire net18178;
 wire net17783;
 wire net17786;
 wire net17788;
 wire net17810;
 wire net17791;
 wire net17816;
 wire net17817;
 wire net17805;
 wire net17809;
 wire net17796;
 wire net17797;
 wire net17798;
 wire net17801;
 wire net17815;
 wire net17807;
 wire net17804;
 wire net18194;
 wire net17812;
 wire net17806;
 wire net17811;
 wire net17813;
 wire net18012;
 wire net18298;
 wire net17988;
 wire net18001;
 wire net17828;
 wire net18438;
 wire net18310;
 wire net18309;
 wire net17989;
 wire net18292;
 wire net18297;
 wire net19156;
 wire net17991;
 wire net17854;
 wire net17995;
 wire net17981;
 wire net17831;
 wire net17836;
 wire net17837;
 wire net17843;
 wire net17999;
 wire net17863;
 wire net17941;
 wire net17861;
 wire net17842;
 wire net18010;
 wire net17853;
 wire net18003;
 wire net17973;
 wire net17908;
 wire net17845;
 wire net17847;
 wire net17855;
 wire net17851;
 wire net17859;
 wire net17852;
 wire net17856;
 wire net17921;
 wire net17867;
 wire net17997;
 wire net17860;
 wire net17870;
 wire net17862;
 wire net17885;
 wire net17868;
 wire net17866;
 wire net17864;
 wire net17873;
 wire net17871;
 wire net17869;
 wire net17879;
 wire net17874;
 wire net18160;
 wire net17965;
 wire net17883;
 wire net17875;
 wire net17872;
 wire net17877;
 wire net17876;
 wire net17880;
 wire net17881;
 wire net17884;
 wire net17909;
 wire net17958;
 wire net17928;
 wire net17905;
 wire net17949;
 wire net17903;
 wire net17925;
 wire net17918;
 wire net17907;
 wire net17891;
 wire net17967;
 wire net17895;
 wire net17893;
 wire net17913;
 wire net17896;
 wire net17898;
 wire net17904;
 wire net17959;
 wire net17923;
 wire net17900;
 wire net17910;
 wire net17902;
 wire net17906;
 wire net17911;
 wire net17914;
 wire net17912;
 wire net17924;
 wire net17917;
 wire net17915;
 wire net17962;
 wire net17916;
 wire net17930;
 wire net17945;
 wire net17919;
 wire net17936;
 wire net17922;
 wire net17926;
 wire net17929;
 wire net17960;
 wire net17979;
 wire net17998;
 wire net17940;
 wire net17931;
 wire net17934;
 wire net17932;
 wire net17937;
 wire net17952;
 wire net17938;
 wire net17933;
 wire net17935;
 wire net17939;
 wire net17942;
 wire net17950;
 wire net17946;
 wire net17947;
 wire net17977;
 wire net17944;
 wire net17971;
 wire net17948;
 wire net17953;
 wire net17951;
 wire net17956;
 wire net17954;
 wire net17955;
 wire net17970;
 wire net17957;
 wire net17961;
 wire net17963;
 wire net17969;
 wire net17964;
 wire net17966;
 wire net17968;
 wire net17990;
 wire net18016;
 wire net17972;
 wire net18009;
 wire net18176;
 wire net17976;
 wire net17974;
 wire net17975;
 wire net17978;
 wire net17982;
 wire net17987;
 wire net17980;
 wire net17986;
 wire net17985;
 wire net17983;
 wire net18002;
 wire net17984;
 wire net18189;
 wire net17992;
 wire net17993;
 wire net18007;
 wire net18000;
 wire net17994;
 wire net17996;
 wire net18004;
 wire net18181;
 wire net18005;
 wire net18188;
 wire net18006;
 wire net18008;
 wire net18165;
 wire net18162;
 wire net18013;
 wire net18148;
 wire net18066;
 wire net18187;
 wire net18011;
 wire net18186;
 wire net18015;
 wire net18041;
 wire net18067;
 wire net18024;
 wire net18023;
 wire net18034;
 wire net18029;
 wire net18020;
 wire net18096;
 wire net18039;
 wire net18025;
 wire net18026;
 wire net18027;
 wire net18033;
 wire net18028;
 wire net18051;
 wire net18032;
 wire net18101;
 wire net18038;
 wire net18037;
 wire net18036;
 wire net18042;
 wire net18040;
 wire net18046;
 wire net18132;
 wire net18072;
 wire net18047;
 wire net18103;
 wire net18053;
 wire net18056;
 wire net18049;
 wire net18052;
 wire net18050;
 wire net18060;
 wire net18076;
 wire net18058;
 wire net18115;
 wire net18063;
 wire net18061;
 wire net18064;
 wire net18071;
 wire net18097;
 wire net18074;
 wire net18102;
 wire net18082;
 wire net18078;
 wire net18124;
 wire net18173;
 wire net18084;
 wire net18091;
 wire net18111;
 wire net18089;
 wire net18087;
 wire net18085;
 wire net18088;
 wire net18090;
 wire net18092;
 wire net18107;
 wire net18095;
 wire net18098;
 wire net18099;
 wire net18100;
 wire net18104;
 wire net18105;
 wire net18108;
 wire net18130;
 wire net18109;
 wire net18122;
 wire net18113;
 wire net18112;
 wire net18119;
 wire net18114;
 wire net18121;
 wire net18120;
 wire net18125;
 wire net18117;
 wire net18116;
 wire net18127;
 wire net18147;
 wire net18128;
 wire net18159;
 wire net18155;
 wire net18158;
 wire net18152;
 wire net18143;
 wire net18131;
 wire net18133;
 wire net18149;
 wire net18138;
 wire net18134;
 wire net18135;
 wire net18137;
 wire net18145;
 wire net18136;
 wire net18141;
 wire net18139;
 wire net18140;
 wire net18142;
 wire net18144;
 wire net18146;
 wire net18169;
 wire net18154;
 wire net18156;
 wire net18150;
 wire net18151;
 wire net18166;
 wire net18153;
 wire net18157;
 wire net18232;
 wire net18161;
 wire net18305;
 wire net18222;
 wire net18185;
 wire net18163;
 wire net18206;
 wire net18180;
 wire net18177;
 wire net18167;
 wire net18170;
 wire net18168;
 wire net18183;
 wire net18174;
 wire net18175;
 wire net18182;
 wire net18179;
 wire net18239;
 wire net18184;
 wire net18238;
 wire net18221;
 wire net18204;
 wire net18201;
 wire net18251;
 wire net18291;
 wire net18234;
 wire net18304;
 wire net18200;
 wire net18199;
 wire net18279;
 wire net18282;
 wire net18294;
 wire net18289;
 wire net18208;
 wire net18207;
 wire net18215;
 wire net18223;
 wire net18209;
 wire net18211;
 wire net19155;
 wire net18303;
 wire net18250;
 wire net18228;
 wire net18216;
 wire net18210;
 wire net18236;
 wire net18212;
 wire net18213;
 wire net18217;
 wire net18214;
 wire net18224;
 wire net18218;
 wire net18225;
 wire net18219;
 wire net18220;
 wire net18226;
 wire net18227;
 wire net18235;
 wire net18233;
 wire net18231;
 wire net18229;
 wire net19110;
 wire net19109;
 wire net18365;
 wire net18283;
 wire net18368;
 wire net18272;
 wire net18355;
 wire net18352;
 wire net18540;
 wire net18333;
 wire net18329;
 wire net18318;
 wire net18321;
 wire net18320;
 wire net18267;
 wire net18275;
 wire net18265;
 wire net18270;
 wire net18255;
 wire net18363;
 wire net18276;
 wire net18257;
 wire net18261;
 wire net18268;
 wire net18260;
 wire net18274;
 wire net18264;
 wire net18266;
 wire net18269;
 wire net18300;
 wire net18301;
 wire net18271;
 wire net18280;
 wire net18273;
 wire net18277;
 wire net18299;
 wire net18287;
 wire net18281;
 wire net18284;
 wire net18285;
 wire net18288;
 wire net18286;
 wire net18290;
 wire net18293;
 wire net18316;
 wire net18295;
 wire net18296;
 wire net18302;
 wire net18449;
 wire net18455;
 wire net18454;
 wire net18444;
 wire net18312;
 wire net18585;
 wire net18534;
 wire net18526;
 wire net18335;
 wire net18596;
 wire net18358;
 wire net18317;
 wire net18343;
 wire net18344;
 wire net18346;
 wire net18410;
 wire net18330;
 wire net18319;
 wire net18323;
 wire net18322;
 wire net18324;
 wire net18327;
 wire net18326;
 wire net18328;
 wire net18334;
 wire net18325;
 wire net18349;
 wire net18424;
 wire net18338;
 wire net18350;
 wire net18331;
 wire net18431;
 wire net18332;
 wire net18337;
 wire net18339;
 wire net18336;
 wire net18340;
 wire net18345;
 wire net18341;
 wire net18342;
 wire net18404;
 wire net18505;
 wire net18595;
 wire net18348;
 wire net18347;
 wire net18786;
 wire net18351;
 wire net18353;
 wire net18594;
 wire net18544;
 wire net18380;
 wire net18376;
 wire net18357;
 wire net18369;
 wire net18354;
 wire net18356;
 wire net18359;
 wire net18374;
 wire net18361;
 wire net18360;
 wire net18362;
 wire net18389;
 wire net18364;
 wire net18366;
 wire net18367;
 wire net18548;
 wire net18373;
 wire net18370;
 wire net18371;
 wire net18372;
 wire net18375;
 wire net18377;
 wire net18383;
 wire net18379;
 wire net18465;
 wire net18546;
 wire net18501;
 wire net18381;
 wire net18547;
 wire net18382;
 wire net18384;
 wire net18472;
 wire net18385;
 wire net18545;
 wire net18386;
 wire net18387;
 wire net18436;
 wire net18433;
 wire net18538;
 wire net18393;
 wire net18390;
 wire net18396;
 wire net18397;
 wire net18399;
 wire net18394;
 wire net18395;
 wire net18403;
 wire net18400;
 wire net18430;
 wire net18401;
 wire net18408;
 wire net18402;
 wire net18405;
 wire net18409;
 wire net18406;
 wire net18407;
 wire net18411;
 wire net18427;
 wire net18413;
 wire net18417;
 wire net18412;
 wire net18414;
 wire net18415;
 wire net18421;
 wire net18416;
 wire net18418;
 wire net18422;
 wire net18419;
 wire net18420;
 wire net18539;
 wire net18543;
 wire net18541;
 wire net18439;
 wire net18432;
 wire net18426;
 wire net18428;
 wire net18429;
 wire net18437;
 wire net18434;
 wire net18435;
 wire net18447;
 wire net18446;
 wire net18442;
 wire net18445;
 wire net18441;
 wire net18452;
 wire net18537;
 wire net18443;
 wire net18450;
 wire net18448;
 wire net18479;
 wire net18469;
 wire net18510;
 wire net18451;
 wire net18453;
 wire net18502;
 wire net18467;
 wire net18458;
 wire net18457;
 wire net18503;
 wire net18464;
 wire net18462;
 wire net18459;
 wire net18468;
 wire net18460;
 wire net18461;
 wire net18463;
 wire net18593;
 wire net18466;
 wire net18482;
 wire net18727;
 wire net18722;
 wire net18488;
 wire net18476;
 wire net18500;
 wire net18592;
 wire net18474;
 wire net18486;
 wire net18475;
 wire net18478;
 wire net18481;
 wire net18483;
 wire net18484;
 wire net18487;
 wire net18490;
 wire net18485;
 wire net18597;
 wire net18491;
 wire net18493;
 wire net18558;
 wire net18492;
 wire net18489;
 wire net18499;
 wire net18496;
 wire net18495;
 wire net18494;
 wire net18498;
 wire net18509;
 wire net18497;
 wire net18504;
 wire net18506;
 wire net18591;
 wire net18523;
 wire net18507;
 wire net18508;
 wire net18512;
 wire net18517;
 wire net18511;
 wire net18590;
 wire net18514;
 wire net18566;
 wire net18524;
 wire net18562;
 wire net18522;
 wire net18527;
 wire net18531;
 wire net18528;
 wire net18601;
 wire net18530;
 wire net18529;
 wire net18609;
 wire net18567;
 wire net18560;
 wire net18602;
 wire net18600;
 wire net18559;
 wire net18608;
 wire net18607;
 wire net18646;
 wire net18721;
 wire net18720;
 wire net18719;
 wire net18631;
 wire net18630;
 wire net18629;
 wire net18628;
 wire net18570;
 wire net18589;
 wire net18561;
 wire net18565;
 wire net18574;
 wire net18636;
 wire net18627;
 wire net18637;
 wire net18603;
 wire net18577;
 wire net18584;
 wire net18564;
 wire net18563;
 wire net18616;
 wire net18580;
 wire net18626;
 wire net18606;
 wire net18604;
 wire net18582;
 wire net18568;
 wire net18569;
 wire net18576;
 wire net18573;
 wire net18571;
 wire net18575;
 wire net18572;
 wire net18581;
 wire net18578;
 wire net18579;
 wire net18587;
 wire net18634;
 wire net18583;
 wire net18586;
 wire net18788;
 wire net18625;
 wire net18624;
 wire net18726;
 wire net18632;
 wire net18621;
 wire net18698;
 wire net18697;
 wire net18680;
 wire net18679;
 wire net18678;
 wire net18645;
 wire net18644;
 wire net18718;
 wire net18643;
 wire net18620;
 wire net18677;
 wire net20435;
 wire net18244;
 wire net18623;
 wire net18962;
 wire net18902;
 wire net18901;
 wire net18694;
 wire net18693;
 wire net18676;
 wire net18692;
 wire net18691;
 wire net18690;
 wire net18689;
 wire net18675;
 wire net18701;
 wire net18688;
 wire net18717;
 wire net18687;
 wire net18686;
 wire net18974;
 wire net18652;
 wire net465;
 wire net18716;
 wire net18973;
 wire net18656;
 wire net18715;
 wire net18972;
 wire net18746;
 wire net18742;
 wire net18714;
 wire net18243;
 wire net18751;
 wire net18785;
 wire net18663;
 wire net18655;
 wire net18668;
 wire net18671;
 wire net19029;
 wire net19027;
 wire net18753;
 wire net18762;
 wire net18725;
 wire net18763;
 wire net18672;
 wire net18737;
 wire net18723;
 wire net19120;
 wire net18993;
 wire net18683;
 wire net18665;
 wire net18736;
 wire net18734;
 wire net18657;
 wire net18654;
 wire net18733;
 wire net18730;
 wire net18658;
 wire net18662;
 wire net18670;
 wire net18667;
 wire net18659;
 wire net18660;
 wire net18669;
 wire net18661;
 wire net18664;
 wire net18666;
 wire net18713;
 wire net18682;
 wire net18732;
 wire net18696;
 wire net18731;
 wire net18705;
 wire net18712;
 wire net18704;
 wire net18710;
 wire net18761;
 wire net18754;
 wire net18706;
 wire net18744;
 wire net18724;
 wire net18760;
 wire net18758;
 wire net18757;
 wire net18756;
 wire net18755;
 wire net18759;
 wire net18740;
 wire net18784;
 wire net18749;
 wire net18783;
 wire net18782;
 wire net18764;
 wire net18739;
 wire net18709;
 wire net18707;
 wire net18770;
 wire net18769;
 wire net18768;
 wire net18752;
 wire net18992;
 wire net18988;
 wire net18738;
 wire net18708;
 wire net18735;
 wire net18767;
 wire net18766;
 wire net18987;
 wire net18741;
 wire net18825;
 wire net18796;
 wire net18780;
 wire net18781;
 wire net18779;
 wire net18778;
 wire net18777;
 wire net18776;
 wire net18775;
 wire net18774;
 wire net18773;
 wire net18792;
 wire net18748;
 wire net18772;
 wire net18824;
 wire net18810;
 wire net18765;
 wire net18801;
 wire net18797;
 wire net18823;
 wire net18986;
 wire net18822;
 wire net18985;
 wire net18771;
 wire net18743;
 wire net18745;
 wire net18747;
 wire net18750;
 wire net18991;
 wire net18787;
 wire net18990;
 wire net18791;
 wire net18989;
 wire net18952;
 wire net18950;
 wire net18911;
 wire net18819;
 wire net18949;
 wire net18964;
 wire net19051;
 wire net18818;
 wire net18904;
 wire net19090;
 wire net18813;
 wire net18817;
 wire net18816;
 wire net18794;
 wire net18815;
 wire net18814;
 wire net18800;
 wire net18798;
 wire net18793;
 wire net19054;
 wire net18866;
 wire net18865;
 wire net18864;
 wire net18820;
 wire net18802;
 wire net18795;
 wire net18809;
 wire net18799;
 wire net19053;
 wire net18977;
 wire net18867;
 wire net18976;
 wire net18804;
 wire net18975;
 wire net18803;
 wire net18899;
 wire net18898;
 wire net18971;
 wire net18897;
 wire net18863;
 wire net18896;
 wire net18808;
 wire net18807;
 wire net18806;
 wire net18805;
 wire net18862;
 wire net18861;
 wire net19092;
 wire net18848;
 wire net18860;
 wire net18834;
 wire net18833;
 wire net18894;
 wire net18893;
 wire net18892;
 wire net18891;
 wire net18878;
 wire net18890;
 wire net18884;
 wire net18871;
 wire net18870;
 wire net18881;
 wire net18853;
 wire net18838;
 wire net18845;
 wire net18882;
 wire net18248;
 wire net18970;
 wire net18969;
 wire net18839;
 wire net18836;
 wire net18918;
 wire net18917;
 wire net18851;
 wire net18847;
 wire net18880;
 wire net18837;
 wire net18888;
 wire net18883;
 wire net18841;
 wire net18842;
 wire net18843;
 wire net18840;
 wire net18879;
 wire net18844;
 wire net18846;
 wire net18875;
 wire net18877;
 wire net18849;
 wire net18869;
 wire net18850;
 wire net18852;
 wire net18868;
 wire net18854;
 wire net19091;
 wire net18900;
 wire net18872;
 wire net18953;
 wire net19184;
 wire net19107;
 wire net18945;
 wire net18932;
 wire net18906;
 wire net18944;
 wire net18247;
 wire net18246;
 wire net18978;
 wire net19037;
 wire net18876;
 wire net18873;
 wire net18889;
 wire net18886;
 wire net19036;
 wire net18885;
 wire net18874;
 wire net18895;
 wire net18903;
 wire net19035;
 wire net18943;
 wire net19034;
 wire net19033;
 wire net18934;
 wire net18916;
 wire net19032;
 wire net18887;
 wire net18930;
 wire net18910;
 wire net18905;
 wire net19031;
 wire net18968;
 wire net18967;
 wire net19030;
 wire net18914;
 wire net19088;
 wire net18913;
 wire net18907;
 wire net19089;
 wire net18998;
 wire net18919;
 wire net19001;
 wire net18965;
 wire net19026;
 wire net19173;
 wire net18908;
 wire net18909;
 wire net18915;
 wire net18912;
 wire net18984;
 wire net18920;
 wire net18983;
 wire net18928;
 wire net18923;
 wire net18966;
 wire net18927;
 wire net18924;
 wire net18982;
 wire net18925;
 wire net18935;
 wire net18931;
 wire net18929;
 wire net18926;
 wire net18979;
 wire net18933;
 wire net18995;
 wire net19172;
 wire net19025;
 wire net19024;
 wire net18947;
 wire net19528;
 wire net18940;
 wire net18936;
 wire net19087;
 wire net18960;
 wire net18937;
 wire net18938;
 wire net19086;
 wire net18939;
 wire net18941;
 wire net18942;
 wire net19019;
 wire net18946;
 wire net18981;
 wire net18957;
 wire net19052;
 wire net18948;
 wire net18980;
 wire net18951;
 wire net18963;
 wire net527;
 wire net18954;
 wire net18955;
 wire net18956;
 wire net18958;
 wire net18961;
 wire net18994;
 wire net19014;
 wire net18245;
 wire net18997;
 wire net18996;
 wire net19028;
 wire net19119;
 wire net17587;
 wire net19050;
 wire net19038;
 wire net19039;
 wire net19049;
 wire net19048;
 wire net19047;
 wire net19000;
 wire net18999;
 wire net17543;
 wire net19085;
 wire net19084;
 wire net19083;
 wire net19003;
 wire net19002;
 wire net19004;
 wire net19106;
 wire net19009;
 wire net19010;
 wire net19007;
 wire net19055;
 wire net19006;
 wire net19011;
 wire net19095;
 wire net19105;
 wire net19104;
 wire net19060;
 wire net19059;
 wire net19016;
 wire net19012;
 wire net19041;
 wire net20432;
 wire net19015;
 wire net19044;
 wire net19022;
 wire net19023;
 wire net19021;
 wire net19005;
 wire net19077;
 wire net19008;
 wire net19020;
 wire net19013;
 wire net19040;
 wire net19018;
 wire net19017;
 wire net19046;
 wire net19058;
 wire net19043;
 wire net19042;
 wire net19045;
 wire net19057;
 wire net19056;
 wire net19171;
 wire net19118;
 wire net19117;
 wire net19116;
 wire net19115;
 wire net19103;
 wire net19075;
 wire net19081;
 wire net19061;
 wire net19074;
 wire net19114;
 wire net19266;
 wire net19160;
 wire net19163;
 wire net19162;
 wire net19097;
 wire net19154;
 wire net19122;
 wire net19102;
 wire net19072;
 wire net19101;
 wire net19100;
 wire net19123;
 wire net19153;
 wire net19152;
 wire net19132;
 wire net19099;
 wire net19065;
 wire net19069;
 wire net19067;
 wire net19062;
 wire net19064;
 wire net19066;
 wire net19068;
 wire net19071;
 wire net19070;
 wire net19073;
 wire net19131;
 wire net19082;
 wire net19079;
 wire net19078;
 wire net19080;
 wire net19108;
 wire net19112;
 wire net19315;
 wire net19124;
 wire net19126;
 wire net19514;
 wire net19130;
 wire net19121;
 wire net19127;
 wire net19128;
 wire net19316;
 wire net19314;
 wire net19529;
 wire net19125;
 wire net19167;
 wire net19161;
 wire net19166;
 wire net19262;
 wire net19313;
 wire net19148;
 wire net19165;
 wire net19164;
 wire net19261;
 wire net19149;
 wire net19257;
 wire net19144;
 wire net19139;
 wire net19256;
 wire net19183;
 wire net19135;
 wire net19600;
 wire net19129;
 wire net19176;
 wire net19136;
 wire net19179;
 wire net19240;
 wire net19239;
 wire net19134;
 wire net19133;
 wire net19137;
 wire net19138;
 wire net19151;
 wire net19140;
 wire net19141;
 wire net19170;
 wire net19145;
 wire net19142;
 wire net19147;
 wire net19168;
 wire net19146;
 wire net19143;
 wire net19169;
 wire net19150;
 wire net19238;
 wire net19237;
 wire net19174;
 wire net19175;
 wire net19178;
 wire net19312;
 wire net19271;
 wire net19270;
 wire net19512;
 wire net19223;
 wire net19212;
 wire net19209;
 wire net19194;
 wire net19192;
 wire net19195;
 wire net19191;
 wire net19273;
 wire net19304;
 wire net19180;
 wire net19181;
 wire net19303;
 wire net19274;
 wire net19300;
 wire net19275;
 wire net19283;
 wire net19249;
 wire net19198;
 wire net19190;
 wire net19182;
 wire net19197;
 wire net19188;
 wire net19196;
 wire net19199;
 wire net19189;
 wire net19193;
 wire net19269;
 wire net19268;
 wire net19311;
 wire net19226;
 wire net19227;
 wire net19208;
 wire net19228;
 wire net19248;
 wire net19251;
 wire net19201;
 wire net19255;
 wire net19207;
 wire net19205;
 wire net19220;
 wire net19200;
 wire net19242;
 wire net19310;
 wire net19258;
 wire net19206;
 wire net19254;
 wire net19202;
 wire net19232;
 wire net19272;
 wire net19234;
 wire net19217;
 wire net19203;
 wire net19210;
 wire net19218;
 wire net19204;
 wire net19211;
 wire net19231;
 wire net19235;
 wire net19214;
 wire net19213;
 wire net19253;
 wire net19215;
 wire net19216;
 wire net19252;
 wire net19247;
 wire net19225;
 wire net19222;
 wire net19219;
 wire net19221;
 wire net19224;
 wire net19230;
 wire net19229;
 wire net19241;
 wire net19246;
 wire net19233;
 wire net19243;
 wire net19265;
 wire net19263;
 wire net19264;
 wire net19260;
 wire net19278;
 wire net19411;
 wire net19331;
 wire net19322;
 wire net19321;
 wire net19309;
 wire net19245;
 wire net19244;
 wire net19308;
 wire net19250;
 wire net19307;
 wire net19320;
 wire net19277;
 wire net19276;
 wire net19285;
 wire net19281;
 wire net19404;
 wire net19783;
 wire net19319;
 wire net19318;
 wire net19295;
 wire net19294;
 wire net19290;
 wire net19293;
 wire net19289;
 wire net19280;
 wire net19286;
 wire net19279;
 wire net19292;
 wire net19291;
 wire net19284;
 wire net19343;
 wire net19361;
 wire net19287;
 wire net19288;
 wire net19370;
 wire net19410;
 wire net19371;
 wire net19298;
 wire net19317;
 wire net19328;
 wire net19385;
 wire net19384;
 wire net19338;
 wire net19299;
 wire net19296;
 wire net19337;
 wire net19334;
 wire net19372;
 wire net19409;
 wire net19326;
 wire net19325;
 wire net19297;
 wire net19302;
 wire net19301;
 wire net19408;
 wire net19324;
 wire net19323;
 wire net19327;
 wire net19330;
 wire net19407;
 wire net19329;
 wire net19360;
 wire net19359;
 wire net19358;
 wire net19339;
 wire net19351;
 wire net19357;
 wire net19356;
 wire net19355;
 wire net19354;
 wire net20679;
 wire net21513;
 wire net21512;
 wire net19341;
 wire net21511;
 wire net19782;
 wire net19335;
 wire net19336;
 wire net19350;
 wire net19349;
 wire net19781;
 wire net19383;
 wire net19382;
 wire net19353;
 wire net19348;
 wire net19347;
 wire net19346;
 wire net19847;
 wire net19696;
 wire net19381;
 wire net19846;
 wire net19821;
 wire net19362;
 wire net19380;
 wire net19368;
 wire net19367;
 wire net19366;
 wire net19352;
 wire net19342;
 wire net19365;
 wire net19364;
 wire net19363;
 wire net19379;
 wire net19378;
 wire net19377;
 wire net19406;
 wire net19376;
 wire net19369;
 wire net19375;
 wire net19779;
 wire net19405;
 wire net19394;
 wire net19397;
 wire net19396;
 wire net19395;
 wire net19392;
 wire net19391;
 wire net19390;
 wire net19389;
 wire net19388;
 wire net19426;
 wire net19486;
 wire net19485;
 wire net19393;
 wire net19415;
 wire net19414;
 wire net19403;
 wire net19413;
 wire net19423;
 wire net19412;
 wire net20451;
 wire net19475;
 wire net19425;
 wire net19474;
 wire net19526;
 wire net19472;
 wire net19464;
 wire net19525;
 wire net19454;
 wire net19402;
 wire net19399;
 wire net19398;
 wire net19460;
 wire net19429;
 wire net19453;
 wire net19400;
 wire net19420;
 wire net19452;
 wire net19419;
 wire net19416;
 wire net19401;
 wire net19422;
 wire net19418;
 wire net19417;
 wire net19421;
 wire net19511;
 wire net19451;
 wire net19427;
 wire net19524;
 wire net498;
 wire net19473;
 wire net19490;
 wire net19428;
 wire net19523;
 wire net19695;
 wire net19489;
 wire net19471;
 wire net19470;
 wire net19694;
 wire net19559;
 wire net19693;
 wire net19853;
 wire net19449;
 wire net19668;
 wire net19459;
 wire net19448;
 wire net19431;
 wire net19430;
 wire net19654;
 wire net19447;
 wire net19432;
 wire net19522;
 wire net19505;
 wire net19488;
 wire net19510;
 wire net19484;
 wire net19467;
 wire net19483;
 wire net19436;
 wire net19434;
 wire net19444;
 wire net19433;
 wire net19458;
 wire net19446;
 wire net19469;
 wire net19468;
 wire net19439;
 wire net19442;
 wire net19438;
 wire net19437;
 wire net19435;
 wire net19457;
 wire net19440;
 wire net19441;
 wire net19443;
 wire net19445;
 wire net19465;
 wire net19463;
 wire net19487;
 wire net19508;
 wire net19504;
 wire net19507;
 wire net19506;
 wire net19509;
 wire net19482;
 wire net19481;
 wire net19480;
 wire net19466;
 wire net19479;
 wire net19478;
 wire net19477;
 wire net19476;
 wire net19521;
 wire net19503;
 wire net19502;
 wire net19496;
 wire net19495;
 wire net19494;
 wire net19493;
 wire net19501;
 wire net19500;
 wire net19497;
 wire net19499;
 wire net19498;
 wire net19520;
 wire net19519;
 wire net19653;
 wire net19518;
 wire net19517;
 wire net19516;
 wire net19515;
 wire net19527;
 wire net20416;
 wire net20450;
 wire net20442;
 wire net20441;
 wire net19558;
 wire net19557;
 wire net19556;
 wire net19555;
 wire net19530;
 wire net19984;
 wire net19554;
 wire net19533;
 wire net19532;
 wire net19599;
 wire net19531;
 wire net20460;
 wire net19553;
 wire net19550;
 wire net19552;
 wire net19551;
 wire net19541;
 wire net19628;
 wire net19540;
 wire net19537;
 wire net19534;
 wire net19539;
 wire net19598;
 wire net19597;
 wire net19538;
 wire net20695;
 wire net19580;
 wire net19581;
 wire net19579;
 wire net19578;
 wire net19577;
 wire net19569;
 wire net19549;
 wire net19542;
 wire net19536;
 wire net19535;
 wire net19545;
 wire net19566;
 wire net20765;
 wire net20602;
 wire net20764;
 wire net20614;
 wire net20613;
 wire net20612;
 wire net20611;
 wire net20588;
 wire net20578;
 wire net19548;
 wire net19544;
 wire net19543;
 wire net19560;
 wire net20490;
 wire net19565;
 wire net19563;
 wire net19546;
 wire net19547;
 wire net19562;
 wire net20439;
 wire net21082;
 wire net19927;
 wire net19639;
 wire net19595;
 wire net19564;
 wire net19582;
 wire net19587;
 wire net19638;
 wire net19576;
 wire net19575;
 wire net19637;
 wire net19570;
 wire net19567;
 wire net19568;
 wire net20262;
 wire net19616;
 wire net19607;
 wire net19594;
 wire net19593;
 wire net19592;
 wire net19586;
 wire net19585;
 wire net19574;
 wire net19573;
 wire net19926;
 wire net19571;
 wire net20261;
 wire net20254;
 wire net19627;
 wire net19617;
 wire net19982;
 wire net19981;
 wire net19584;
 wire net19572;
 wire net19591;
 wire net19583;
 wire net19596;
 wire net19980;
 wire net19590;
 wire net19589;
 wire net19979;
 wire net19640;
 wire net19588;
 wire net19606;
 wire net19605;
 wire net19604;
 wire net19602;
 wire net19601;
 wire net20418;
 wire net19978;
 wire net19636;
 wire net19648;
 wire net19647;
 wire net19603;
 wire net19646;
 wire net19645;
 wire net19767;
 wire net19613;
 wire net19612;
 wire net19634;
 wire net19615;
 wire net19614;
 wire net19609;
 wire net19610;
 wire net19608;
 wire net19611;
 wire net19936;
 wire net19914;
 wire net19895;
 wire net19917;
 wire net19951;
 wire net19859;
 wire net19619;
 wire net19644;
 wire net19621;
 wire net19633;
 wire net19626;
 wire net19629;
 wire net19623;
 wire net19652;
 wire net19823;
 wire net19632;
 wire net19631;
 wire net19625;
 wire net19618;
 wire net19630;
 wire net19620;
 wire net19622;
 wire net19983;
 wire net20942;
 wire net19624;
 wire net19857;
 wire net20678;
 wire net19685;
 wire net19674;
 wire net19662;
 wire net19660;
 wire net19659;
 wire net19655;
 wire net19658;
 wire net19635;
 wire net19657;
 wire net19656;
 wire net19651;
 wire net19643;
 wire net19642;
 wire net19641;
 wire net19977;
 wire net19650;
 wire net19692;
 wire net19649;
 wire net19661;
 wire net19820;
 wire net19691;
 wire net19345;
 wire net19344;
 wire net19684;
 wire net19683;
 wire net19669;
 wire net19852;
 wire net19667;
 wire net19666;
 wire net19675;
 wire net19665;
 wire net19664;
 wire net19663;
 wire net19333;
 wire net19766;
 wire net19851;
 wire net19677;
 wire net19670;
 wire net19676;
 wire net19671;
 wire net19778;
 wire net19682;
 wire net19681;
 wire net19673;
 wire net19680;
 wire net19672;
 wire net19819;
 wire net19690;
 wire net19710;
 wire net19689;
 wire net19688;
 wire net19687;
 wire net19679;
 wire net19678;
 wire net19764;
 wire net19763;
 wire net19756;
 wire net19755;
 wire net19709;
 wire net19698;
 wire net19686;
 wire net19850;
 wire net19848;
 wire net19697;
 wire net19717;
 wire net19716;
 wire net19715;
 wire net19706;
 wire net19705;
 wire net19701;
 wire net19700;
 wire net19699;
 wire net19708;
 wire net19340;
 wire net19373;
 wire net19386;
 wire net19762;
 wire net19761;
 wire net19760;
 wire net19704;
 wire net19703;
 wire net19751;
 wire net19707;
 wire net19702;
 wire net19387;
 wire net19374;
 wire net19718;
 wire net19259;
 wire net19561;
 wire net19730;
 wire net19236;
 wire net19185;
 wire net19721;
 wire net19729;
 wire net19785;
 wire net19711;
 wire net19738;
 wire net19714;
 wire net19712;
 wire net21096;
 wire net19713;
 wire net19726;
 wire net19737;
 wire net19753;
 wire net19728;
 wire net19723;
 wire net19727;
 wire net19720;
 wire net19719;
 wire net19187;
 wire net19734;
 wire net19186;
 wire net19113;
 wire net18648;
 wire net19733;
 wire net19098;
 wire net18650;
 wire net18649;
 wire net19111;
 wire net19096;
 wire net18711;
 wire net18703;
 wire net18702;
 wire net18685;
 wire net18684;
 wire net19754;
 wire net19722;
 wire net19736;
 wire net19725;
 wire net19752;
 wire net18681;
 wire net19724;
 wire net18674;
 wire net19732;
 wire net18673;
 wire net18653;
 wire net18647;
 wire net18642;
 wire net18641;
 wire net18640;
 wire net21510;
 wire net19759;
 wire net19749;
 wire net18699;
 wire net19731;
 wire net19744;
 wire net19735;
 wire net19739;
 wire net19740;
 wire net19746;
 wire net19741;
 wire net19743;
 wire net19817;
 wire net19742;
 wire net19745;
 wire net19795;
 wire net19777;
 wire net19748;
 wire net19747;
 wire net19750;
 wire net19773;
 wire net19758;
 wire net19757;
 wire net19765;
 wire net19772;
 wire net21509;
 wire net19768;
 wire net19784;
 wire net19816;
 wire net19769;
 wire net19771;
 wire net21508;
 wire net19770;
 wire net18639;
 wire net18638;
 wire net18619;
 wire net20677;
 wire net20676;
 wire net20675;
 wire net19776;
 wire net19818;
 wire net19775;
 wire net19774;
 wire net19856;
 wire net18622;
 wire net19813;
 wire net21507;
 wire net19794;
 wire net19786;
 wire net19793;
 wire net19792;
 wire net19791;
 wire net21506;
 wire net19843;
 wire net19809;
 wire net19832;
 wire net19831;
 wire net19787;
 wire net19780;
 wire net19812;
 wire net19804;
 wire net19799;
 wire net19815;
 wire net19788;
 wire net19790;
 wire net19789;
 wire net19798;
 wire net19800;
 wire net19797;
 wire net19796;
 wire net19830;
 wire net21134;
 wire net19814;
 wire net19803;
 wire net19829;
 wire net19828;
 wire net21505;
 wire net19801;
 wire net21504;
 wire net19845;
 wire net18617;
 wire net18618;
 wire net18605;
 wire net20694;
 wire net19855;
 wire net19805;
 wire net19810;
 wire net19802;
 wire net19807;
 wire net19824;
 wire net19854;
 wire net19806;
 wire net19811;
 wire net19822;
 wire net19808;
 wire net20760;
 wire net19844;
 wire net18470;
 wire net18473;
 wire net19918;
 wire net19858;
 wire net19826;
 wire net19825;
 wire net20733;
 wire net20736;
 wire net20674;
 wire net19839;
 wire net19838;
 wire net19916;
 wire net18440;
 wire net20232;
 wire net19947;
 wire net19864;
 wire net19863;
 wire net19862;
 wire net19861;
 wire net19949;
 wire net19868;
 wire net19835;
 wire net19837;
 wire net20574;
 wire net19827;
 wire net19833;
 wire net19834;
 wire net19836;
 wire net19939;
 wire net19867;
 wire net19938;
 wire net19866;
 wire net21081;
 wire net19842;
 wire net19841;
 wire net19948;
 wire net19919;
 wire net19950;
 wire net19840;
 wire net19860;
 wire net19937;
 wire net19865;
 wire net19920;
 wire net19976;
 wire net19957;
 wire net19961;
 wire net19953;
 wire net19970;
 wire net19966;
 wire net20253;
 wire net20252;
 wire net19900;
 wire net19877;
 wire net19935;
 wire net19930;
 wire net19869;
 wire net19870;
 wire net19886;
 wire net19888;
 wire net19885;
 wire net19876;
 wire net19929;
 wire net19928;
 wire net19871;
 wire net19907;
 wire net19875;
 wire net19874;
 wire net19872;
 wire net19896;
 wire net19878;
 wire net19965;
 wire net21080;
 wire net19873;
 wire net20250;
 wire net19923;
 wire net19922;
 wire net19880;
 wire net19884;
 wire net19889;
 wire net19879;
 wire net19881;
 wire net19882;
 wire net19883;
 wire net19915;
 wire net19887;
 wire net19894;
 wire net19890;
 wire net19891;
 wire net19903;
 wire net19893;
 wire net19892;
 wire net19902;
 wire net19898;
 wire net19897;
 wire net19899;
 wire net19901;
 wire net20249;
 wire net19921;
 wire net19904;
 wire net19912;
 wire net19905;
 wire net19906;
 wire net19908;
 wire net19911;
 wire net19910;
 wire net19909;
 wire net20243;
 wire net20210;
 wire net19969;
 wire net19913;
 wire net19964;
 wire net19925;
 wire net19990;
 wire net20061;
 wire net19924;
 wire net19989;
 wire net19956;
 wire net19946;
 wire net19932;
 wire net19988;
 wire net19941;
 wire net19940;
 wire net19934;
 wire net19955;
 wire net19954;
 wire net19931;
 wire net19933;
 wire net20073;
 wire net19975;
 wire net19974;
 wire net19944;
 wire net20075;
 wire net19958;
 wire net19960;
 wire net19952;
 wire net19942;
 wire net19943;
 wire net20069;
 wire net20064;
 wire net19987;
 wire net19962;
 wire net19963;
 wire net19959;
 wire net19968;
 wire net19967;
 wire net19945;
 wire net19986;
 wire net19973;
 wire net20124;
 wire net20136;
 wire net21079;
 wire net21078;
 wire net20033;
 wire net20032;
 wire net19996;
 wire net19995;
 wire net19972;
 wire net20114;
 wire net20022;
 wire net20389;
 wire net20269;
 wire net20236;
 wire net20012;
 wire net19971;
 wire net19994;
 wire net19991;
 wire net19985;
 wire net19993;
 wire net20390;
 wire net20251;
 wire net19992;
 wire net20005;
 wire net20003;
 wire net19999;
 wire net19997;
 wire net20004;
 wire net21077;
 wire net20241;
 wire net20226;
 wire net20192;
 wire net20183;
 wire net20173;
 wire net20225;
 wire net20167;
 wire net20016;
 wire net20157;
 wire net20002;
 wire net20001;
 wire net19998;
 wire net20011;
 wire net20006;
 wire net20020;
 wire net20208;
 wire net20350;
 wire net20030;
 wire net20277;
 wire net20273;
 wire net20019;
 wire net20018;
 wire net20000;
 wire net20029;
 wire net20028;
 wire net20027;
 wire net20010;
 wire net20060;
 wire net20015;
 wire net20014;
 wire net20007;
 wire net20013;
 wire net20008;
 wire net20017;
 wire net20156;
 wire net20059;
 wire net20049;
 wire net20009;
 wire net20048;
 wire net20021;
 wire net20031;
 wire net20802;
 wire net20190;
 wire net20268;
 wire net20263;
 wire net20026;
 wire net20037;
 wire net20054;
 wire net20025;
 wire net20034;
 wire net20139;
 wire net20207;
 wire net20023;
 wire net20053;
 wire net20169;
 wire net20055;
 wire net20050;
 wire net20046;
 wire net20042;
 wire net20040;
 wire net20041;
 wire net20024;
 wire net20036;
 wire net20035;
 wire net20181;
 wire net20172;
 wire net20171;
 wire net20044;
 wire net20043;
 wire net20058;
 wire net20039;
 wire net20038;
 wire net20083;
 wire net20066;
 wire net20047;
 wire net20057;
 wire net20062;
 wire net20164;
 wire net20163;
 wire net20045;
 wire net20063;
 wire net20056;
 wire net20051;
 wire net20363;
 wire net20166;
 wire net20138;
 wire net20077;
 wire net20103;
 wire net20100;
 wire net20052;
 wire net20125;
 wire net20085;
 wire net20143;
 wire net20209;
 wire net20135;
 wire net20222;
 wire net20130;
 wire net20065;
 wire net20067;
 wire net20165;
 wire net20068;
 wire net20086;
 wire net20070;
 wire net20162;
 wire net20071;
 wire net20072;
 wire net20161;
 wire net20082;
 wire net20074;
 wire net20076;
 wire net20079;
 wire net20078;
 wire net20080;
 wire net20081;
 wire net20084;
 wire net20094;
 wire net20145;
 wire net20089;
 wire net20126;
 wire net20087;
 wire net20092;
 wire net20088;
 wire net20091;
 wire net20129;
 wire net20090;
 wire net20096;
 wire net20098;
 wire net20095;
 wire net20097;
 wire net20093;
 wire net20099;
 wire net20113;
 wire net20106;
 wire net20105;
 wire net20102;
 wire net20101;
 wire net20111;
 wire net20104;
 wire net20108;
 wire net20116;
 wire net20107;
 wire net20110;
 wire net20109;
 wire net20112;
 wire net20122;
 wire net20117;
 wire net20115;
 wire net20118;
 wire net20119;
 wire net20120;
 wire net20121;
 wire net20123;
 wire net20127;
 wire net20224;
 wire net20128;
 wire net20131;
 wire net20133;
 wire net20485;
 wire net20479;
 wire net20132;
 wire net20154;
 wire net20150;
 wire net20134;
 wire net20137;
 wire net20149;
 wire net20140;
 wire net20141;
 wire net20142;
 wire net20146;
 wire net20144;
 wire net20147;
 wire net20168;
 wire net20153;
 wire net20148;
 wire net20151;
 wire net20158;
 wire net20481;
 wire net20152;
 wire net20155;
 wire net20475;
 wire net20170;
 wire net20159;
 wire net20160;
 wire net20175;
 wire net20177;
 wire net20193;
 wire net20191;
 wire net20174;
 wire net20176;
 wire net20474;
 wire net20214;
 wire net20413;
 wire net20182;
 wire net20178;
 wire net20405;
 wire net20206;
 wire net20502;
 wire net20473;
 wire net20179;
 wire net20188;
 wire net20184;
 wire net20180;
 wire net20189;
 wire net20491;
 wire net20488;
 wire net20186;
 wire net20550;
 wire net20185;
 wire net20471;
 wire net20503;
 wire net20577;
 wire net20204;
 wire net20187;
 wire net20194;
 wire net20195;
 wire net20199;
 wire net20196;
 wire net20212;
 wire net20399;
 wire net20198;
 wire net20203;
 wire net20202;
 wire net20197;
 wire net20201;
 wire net20213;
 wire net20200;
 wire net20211;
 wire net20205;
 wire net20242;
 wire net20227;
 wire net20422;
 wire net20573;
 wire net20220;
 wire net20215;
 wire net20395;
 wire net18425;
 wire net20267;
 wire net20266;
 wire net20265;
 wire net20500;
 wire net20223;
 wire net20499;
 wire net20388;
 wire net20216;
 wire net20372;
 wire net20217;
 wire net20415;
 wire net20259;
 wire net20343;
 wire net20351;
 wire net20360;
 wire net20228;
 wire net20219;
 wire net20218;
 wire net20374;
 wire net20221;
 wire net20229;
 wire net20248;
 wire net20233;
 wire net20235;
 wire net20237;
 wire net20238;
 wire net20230;
 wire net20231;
 wire net20234;
 wire net20240;
 wire net20239;
 wire net20255;
 wire net20244;
 wire net20245;
 wire net20246;
 wire net18423;
 wire net18542;
 wire net20593;
 wire net20271;
 wire net20247;
 wire net20258;
 wire net20260;
 wire net20256;
 wire net20766;
 wire net20272;
 wire net20601;
 wire net20572;
 wire net20276;
 wire net20362;
 wire net20270;
 wire net20257;
 wire net20264;
 wire net20275;
 wire net18398;
 wire net18391;
 wire net18259;
 wire net20274;
 wire net20311;
 wire net20319;
 wire net20342;
 wire net20278;
 wire net20335;
 wire net20349;
 wire net20344;
 wire net20301;
 wire net20334;
 wire net20291;
 wire net20279;
 wire net20409;
 wire net20407;
 wire net20394;
 wire net20411;
 wire net20381;
 wire net20315;
 wire net18258;
 wire net20292;
 wire net20288;
 wire net20285;
 wire net20283;
 wire net20298;
 wire net20280;
 wire net20281;
 wire net20286;
 wire net20282;
 wire net20289;
 wire net20284;
 wire net18262;
 wire net20313;
 wire net20287;
 wire net20290;
 wire net20331;
 wire net20293;
 wire net20296;
 wire net20299;
 wire net20294;
 wire net20295;
 wire net18256;
 wire net18254;
 wire net20307;
 wire net20312;
 wire net20297;
 wire net20300;
 wire net20309;
 wire net20302;
 wire net20303;
 wire net20304;
 wire net20305;
 wire net20306;
 wire net20308;
 wire net20310;
 wire net18253;
 wire net20314;
 wire net20318;
 wire net20316;
 wire net20317;
 wire net20325;
 wire net18315;
 wire net20322;
 wire net20321;
 wire net20320;
 wire net20340;
 wire net20323;
 wire net20333;
 wire net20324;
 wire net20326;
 wire net20361;
 wire net20327;
 wire net20329;
 wire net20328;
 wire net20337;
 wire net20332;
 wire net20330;
 wire net20336;
 wire net20375;
 wire net18314;
 wire net20338;
 wire net20346;
 wire net20348;
 wire net18313;
 wire net18311;
 wire net20339;
 wire net20341;
 wire net20345;
 wire net20347;
 wire net20358;
 wire net20356;
 wire net20353;
 wire net20354;
 wire net20352;
 wire net20357;
 wire net20355;
 wire net20359;
 wire net18263;
 wire net20369;
 wire net20383;
 wire net20385;
 wire net20364;
 wire net20365;
 wire net20367;
 wire net18308;
 wire net20376;
 wire net18205;
 wire net20366;
 wire net20368;
 wire net20370;
 wire net18198;
 wire net18197;
 wire net20386;
 wire net20371;
 wire net20384;
 wire net20373;
 wire net20377;
 wire net20378;
 wire net20379;
 wire net20380;
 wire net20382;
 wire net20393;
 wire net20391;
 wire net20387;
 wire net20587;
 wire net20392;
 wire net20410;
 wire net20498;
 wire net20487;
 wire net20401;
 wire net20496;
 wire net20406;
 wire net20586;
 wire net20397;
 wire net20396;
 wire net20571;
 wire net20400;
 wire net20398;
 wire net20425;
 wire net20402;
 wire net20403;
 wire net20404;
 wire net20570;
 wire net20424;
 wire net20421;
 wire net20417;
 wire net20412;
 wire net20408;
 wire net20414;
 wire net20446;
 wire net20438;
 wire net20419;
 wire net20445;
 wire net20420;
 wire net20497;
 wire net20428;
 wire net20434;
 wire net20427;
 wire net20423;
 wire net20510;
 wire net20426;
 wire net20472;
 wire net20430;
 wire net20429;
 wire net20440;
 wire net20431;
 wire net20433;
 wire net20437;
 wire net20452;
 wire net20551;
 wire net20457;
 wire net20456;
 wire net20470;
 wire net20549;
 wire net20447;
 wire net20448;
 wire net20443;
 wire net20444;
 wire net20534;
 wire net20564;
 wire net20576;
 wire net20501;
 wire net20458;
 wire net20568;
 wire net20569;
 wire net20493;
 wire net20492;
 wire net20449;
 wire net20453;
 wire net20553;
 wire net20454;
 wire net20455;
 wire net20552;
 wire net20567;
 wire net20548;
 wire net20563;
 wire net20559;
 wire net18171;
 wire net20480;
 wire net20478;
 wire net20476;
 wire net20477;
 wire net18172;
 wire net18164;
 wire net18086;
 wire net18083;
 wire net18129;
 wire net18118;
 wire net18123;
 wire net18126;
 wire net18110;
 wire net20484;
 wire net20511;
 wire net18081;
 wire net18080;
 wire net20482;
 wire net18079;
 wire net18077;
 wire net20483;
 wire net20546;
 wire net20486;
 wire net20538;
 wire net20489;
 wire net20495;
 wire net20504;
 wire net20494;
 wire net20537;
 wire net20547;
 wire net20518;
 wire net20505;
 wire net20536;
 wire net20506;
 wire net18075;
 wire net20535;
 wire net20507;
 wire net18070;
 wire net18069;
 wire net18062;
 wire net20610;
 wire net20596;
 wire net20595;
 wire net20515;
 wire net20508;
 wire net20509;
 wire net20528;
 wire net20512;
 wire net20516;
 wire net20562;
 wire net20527;
 wire net20513;
 wire net20558;
 wire net20514;
 wire net20517;
 wire net20557;
 wire net20544;
 wire net20554;
 wire net20543;
 wire net20526;
 wire net20524;
 wire net20519;
 wire net20520;
 wire net20531;
 wire net20521;
 wire net20523;
 wire net20529;
 wire net20522;
 wire net20525;
 wire net20530;
 wire net20561;
 wire net20545;
 wire net20533;
 wire net20532;
 wire net20540;
 wire net20539;
 wire net20560;
 wire net20541;
 wire net20594;
 wire net20600;
 wire net20556;
 wire net20555;
 wire net20599;
 wire net20585;
 wire net20542;
 wire net20565;
 wire net20575;
 wire net20566;
 wire net20584;
 wire net20609;
 wire net18065;
 wire net18059;
 wire net18057;
 wire net18068;
 wire net18055;
 wire net18054;
 wire net18048;
 wire net20621;
 wire net20583;
 wire net20582;
 wire net20581;
 wire net20579;
 wire net20580;
 wire net20616;
 wire net20673;
 wire net20672;
 wire net20597;
 wire net20598;
 wire net20636;
 wire net20693;
 wire net20608;
 wire net20607;
 wire net20656;
 wire net20692;
 wire net20604;
 wire net20603;
 wire net20606;
 wire net20605;
 wire net20691;
 wire net20690;
 wire net20658;
 wire net20615;
 wire net20662;
 wire net20661;
 wire net20660;
 wire net20657;
 wire net20659;
 wire net20649;
 wire net20633;
 wire net20732;
 wire net20625;
 wire net20731;
 wire net20735;
 wire net20689;
 wire net20648;
 wire net20618;
 wire net20635;
 wire net18073;
 wire net18045;
 wire net20686;
 wire net20626;
 wire net20685;
 wire net20684;
 wire net20683;
 wire net20682;
 wire net20681;
 wire net20671;
 wire net18044;
 wire net20670;
 wire net20666;
 wire net18043;
 wire net18035;
 wire net18031;
 wire net18030;
 wire net20619;
 wire net20617;
 wire net18022;
 wire net18021;
 wire net20631;
 wire net20627;
 wire net20620;
 wire net20622;
 wire net20680;
 wire net20623;
 wire net20624;
 wire net20628;
 wire net20663;
 wire net20630;
 wire net20653;
 wire net20632;
 wire net17897;
 wire net20651;
 wire net17894;
 wire net20634;
 wire net20647;
 wire net20644;
 wire net20650;
 wire net20641;
 wire net20637;
 wire net20655;
 wire net20638;
 wire net17892;
 wire net17899;
 wire net20643;
 wire net20639;
 wire net17889;
 wire net17887;
 wire net20640;
 wire net20642;
 wire net17901;
 wire net20645;
 wire net17886;
 wire net17882;
 wire net17943;
 wire net20646;
 wire net20654;
 wire net20652;
 wire net17835;
 wire net17841;
 wire net17927;
 wire net17840;
 wire net17839;
 wire net17834;
 wire net20730;
 wire net20702;
 wire net20734;
 wire net20697;
 wire net20668;
 wire net20669;
 wire net20665;
 wire net20664;
 wire net20688;
 wire net20701;
 wire net17829;
 wire net17742;
 wire net20667;
 wire net17827;
 wire net17752;
 wire net17750;
 wire net17787;
 wire net17753;
 wire net17795;
 wire net17766;
 wire net17764;
 wire net17779;
 wire net17763;
 wire net17738;
 wire net17728;
 wire net17722;
 wire net20699;
 wire net19094;
 wire net20698;
 wire net20687;
 wire net19093;
 wire net20938;
 wire net20759;
 wire net20758;
 wire net20700;
 wire net20756;
 wire net20726;
 wire net20725;
 wire net20711;
 wire net20717;
 wire net20729;
 wire net20763;
 wire net20755;
 wire net20719;
 wire net20706;
 wire net20754;
 wire net20727;
 wire net20720;
 wire net20705;
 wire net20716;
 wire net17720;
 wire net20724;
 wire net20753;
 wire net18094;
 wire net18093;
 wire net20713;
 wire net20709;
 wire net20708;
 wire net18019;
 wire net18018;
 wire net18635;
 wire net18831;
 wire net20712;
 wire net21070;
 wire net20728;
 wire net21069;
 wire net20932;
 wire net20891;
 wire net21068;
 wire net20722;
 wire net20723;
 wire net20718;
 wire net21037;
 wire net20721;
 wire net20752;
 wire net20740;
 wire net20739;
 wire net20738;
 wire net21030;
 wire net20751;
 wire net20744;
 wire net20743;
 wire net20742;
 wire net20741;
 wire net20747;
 wire net21029;
 wire net20774;
 wire net20773;
 wire net20787;
 wire net20955;
 wire net18830;
 wire net20780;
 wire net20775;
 wire net20786;
 wire net20771;
 wire net20770;
 wire net20746;
 wire net20745;
 wire net20804;
 wire net20785;
 wire net18017;
 wire net20750;
 wire net20769;
 wire net18193;
 wire net18230;
 wire net18203;
 wire net21075;
 wire net21074;
 wire net21073;
 wire net21072;
 wire net20830;
 wire net20792;
 wire net20748;
 wire net20749;
 wire net18192;
 wire net20772;
 wire net20829;
 wire net20768;
 wire net20767;
 wire net20757;
 wire net20784;
 wire net20861;
 wire net20798;
 wire net18829;
 wire net20828;
 wire net20826;
 wire net20776;
 wire net20779;
 wire net20778;
 wire net18202;
 wire net20855;
 wire net20801;
 wire net20800;
 wire net20799;
 wire net20790;
 wire net20854;
 wire net20808;
 wire net20777;
 wire net18237;
 wire net20850;
 wire net20841;
 wire net20793;
 wire net20783;
 wire net20781;
 wire net20782;
 wire net20791;
 wire net20789;
 wire net20788;
 wire net20807;
 wire net20797;
 wire net20803;
 wire net18828;
 wire net18196;
 wire net18195;
 wire net17838;
 wire net20796;
 wire net20795;
 wire net20853;
 wire net20794;
 wire net17833;
 wire net17826;
 wire net21076;
 wire net20812;
 wire net18191;
 wire net20805;
 wire net20825;
 wire net20809;
 wire net18106;
 wire net17712;
 wire net20819;
 wire net20816;
 wire net20806;
 wire net17715;
 wire net17692;
 wire net17688;
 wire net17654;
 wire net17647;
 wire net17640;
 wire net20837;
 wire net17646;
 wire net17652;
 wire net20815;
 wire net20810;
 wire net20840;
 wire net20813;
 wire net20814;
 wire net20852;
 wire net20818;
 wire net20811;
 wire net20817;
 wire net20851;
 wire net20839;
 wire net17699;
 wire net21103;
 wire net17696;
 wire net20827;
 wire net20821;
 wire net20820;
 wire net20822;
 wire net20824;
 wire net20823;
 wire net20832;
 wire net18190;
 wire net20836;
 wire net20831;
 wire net21503;
 wire net20925;
 wire net20908;
 wire net20881;
 wire net20835;
 wire net20834;
 wire net20879;
 wire net20833;
 wire net20860;
 wire net20878;
 wire net17890;
 wire net17705;
 wire net17694;
 wire net20877;
 wire net17633;
 wire net17645;
 wire net20875;
 wire net20864;
 wire net20838;
 wire net20856;
 wire net20842;
 wire net20848;
 wire net20843;
 wire net21099;
 wire net17638;
 wire net17537;
 wire net20844;
 wire net20931;
 wire net17541;
 wire net20858;
 wire net20845;
 wire net20847;
 wire net20846;
 wire net20849;
 wire net21071;
 wire net20857;
 wire net20907;
 wire net20862;
 wire net20900;
 wire net20899;
 wire net20910;
 wire net20897;
 wire net20870;
 wire net20866;
 wire net20863;
 wire net20887;
 wire net17878;
 wire net17888;
 wire net20859;
 wire net17698;
 wire net21522;
 wire net21521;
 wire net20949;
 wire net21502;
 wire net20873;
 wire net17865;
 wire net20880;
 wire net20865;
 wire net20930;
 wire net20872;
 wire net20869;
 wire net20867;
 wire net20868;
 wire net20871;
 wire net20915;
 wire net21514;
 wire net21520;
 wire net20876;
 wire net20895;
 wire net20874;
 wire net21098;
 wire net20884;
 wire net20890;
 wire net21097;
 wire net20882;
 wire net21519;
 wire net21517;
 wire net20885;
 wire net20883;
 wire net20892;
 wire net20886;
 wire net20888;
 wire net20889;
 wire net20901;
 wire net20893;
 wire net20894;
 wire net20896;
 wire net20904;
 wire net20898;
 wire net20905;
 wire net21119;
 wire net21516;
 wire net20902;
 wire net20903;
 wire net20906;
 wire net20923;
 wire net20928;
 wire net20924;
 wire net20922;
 wire net20909;
 wire net20920;
 wire net20911;
 wire net20917;
 wire net20912;
 wire net20914;
 wire net20916;
 wire net21530;
 wire net20929;
 wire net20919;
 wire net20918;
 wire net20921;
 wire net20926;
 wire net20927;
 wire net17514;
 wire net17511;
 wire net21128;
 wire net21425;
 wire net17507;
 wire net21524;
 wire net20933;
 wire net21523;
 wire net21501;
 wire net21500;
 wire net21275;
 wire net21529;
 wire net21499;
 wire net20934;
 wire net20937;
 wire net17504;
 wire net17499;
 wire net20935;
 wire net21409;
 wire net17498;
 wire net20936;
 wire net21527;
 wire net21526;
 wire net21424;
 wire net21498;
 wire net21497;
 wire net20940;
 wire net20939;
 wire net20941;
 wire net20943;
 wire net17510;
 wire net20944;
 wire net20945;
 wire net20946;
 wire net20947;
 wire net20964;
 wire net20948;
 wire net20951;
 wire net21496;
 wire net20970;
 wire net20950;
 wire net20952;
 wire net21495;
 wire net20953;
 wire net20954;
 wire net21542;
 wire net21538;
 wire net20956;
 wire net21494;
 wire net20957;
 wire net20958;
 wire net20959;
 wire net20960;
 wire net20962;
 wire net20961;
 wire net17495;
 wire net21518;
 wire net17494;
 wire net21515;
 wire net17480;
 wire net17478;
 wire net17486;
 wire net17466;
 wire net17442;
 wire net21051;
 wire net20965;
 wire net20995;
 wire net20963;
 wire net20969;
 wire net21525;
 wire net21026;
 wire net20966;
 wire net21528;
 wire net21414;
 wire net20968;
 wire net20973;
 wire net20967;
 wire net20971;
 wire net21015;
 wire net21306;
 wire net21012;
 wire net20987;
 wire net21021;
 wire net20972;
 wire net20976;
 wire net20974;
 wire clknet_leaf_35_clk;
 wire net21017;
 wire net20999;
 wire net20975;
 wire net20981;
 wire net20977;
 wire net20978;
 wire net20997;
 wire net20984;
 wire net20979;
 wire net21001;
 wire net20980;
 wire net21341;
 wire net20982;
 wire net20983;
 wire net21305;
 wire net20985;
 wire net20986;
 wire net20988;
 wire net20989;
 wire net20990;
 wire net20991;
 wire net20992;
 wire net20993;
 wire net21000;
 wire net20994;
 wire net20998;
 wire net20996;
 wire net21294;
 wire net21413;
 wire net21005;
 wire net21003;
 wire net21007;
 wire net21002;
 wire net21004;
 wire net21006;
 wire net21009;
 wire clknet_leaf_30_clk;
 wire net21008;
 wire net21014;
 wire net21543;
 wire net21010;
 wire net21011;
 wire net21013;
 wire net21458;
 wire net21439;
 wire net21323;
 wire net21018;
 wire net21016;
 wire net21036;
 wire net21019;
 wire net21050;
 wire net21042;
 wire net21060;
 wire net21020;
 wire net21022;
 wire net21023;
 wire net21025;
 wire net21024;
 wire net21027;
 wire net21028;
 wire net21031;
 wire net21049;
 wire net21032;
 wire net21033;
 wire net21040;
 wire net21034;
 wire net21039;
 wire net21038;
 wire net21035;
 wire net21043;
 wire net21041;
 wire net21067;
 wire net21061;
 wire net21044;
 wire net21308;
 wire net21456;
 wire net21045;
 wire net21046;
 wire net21047;
 wire net21048;
 wire net21488;
 wire net21056;
 wire net21065;
 wire net21052;
 wire net17437;
 wire net17462;
 wire net21053;
 wire net21054;
 wire net21055;
 wire net21057;
 wire net21058;
 wire net21313;
 wire net21064;
 wire net21059;
 wire net21063;
 wire net21062;
 wire net21066;
 wire net21309;
 wire net21487;
 wire net17452;
 wire net17651;
 wire net17425;
 wire net21105;
 wire net21100;
 wire net21123;
 wire net17641;
 wire net17639;
 wire net17636;
 wire net17426;
 wire net17634;
 wire net426;
 wire net17632;
 wire net17566;
 wire net17562;
 wire net17447;
 wire net17438;
 wire net17435;
 wire net17563;
 wire net17444;
 wire net17557;
 wire net17615;
 wire net17440;
 wire net17439;
 wire net17569;
 wire net17455;
 wire net17553;
 wire net17474;
 wire net17477;
 wire net17458;
 wire net17558;
 wire net17551;
 wire net17481;
 wire net17476;
 wire net17631;
 wire net17554;
 wire net17556;
 wire net17550;
 wire net17549;
 wire net21112;
 wire net21104;
 wire net21101;
 wire net21102;
 wire net17427;
 wire net21111;
 wire net21106;
 wire net21107;
 wire net21108;
 wire net21109;
 wire net21110;
 wire net17420;
 wire net17414;
 wire net21120;
 wire net21116;
 wire net21121;
 wire net21113;
 wire net21114;
 wire net21115;
 wire net21117;
 wire net21118;
 wire net21131;
 wire net21272;
 wire net17419;
 wire net21122;
 wire net21124;
 wire net21249;
 wire net21244;
 wire net21138;
 wire net21126;
 wire net21266;
 wire net21125;
 wire net21129;
 wire net21535;
 wire net21130;
 wire net21127;
 wire net21534;
 wire net21532;
 wire net21133;
 wire net21132;
 wire net21531;
 wire net21135;
 wire net21136;
 wire net21137;
 wire net21139;
 wire net21140;
 wire net21165;
 wire net21141;
 wire net21149;
 wire net21142;
 wire net21143;
 wire net21144;
 wire net21145;
 wire net21146;
 wire net21147;
 wire net21179;
 wire net21148;
 wire net21150;
 wire net21151;
 wire net21152;
 wire net21153;
 wire net21154;
 wire net21155;
 wire net21156;
 wire net21157;
 wire net21158;
 wire net21159;
 wire net21160;
 wire net21161;
 wire net21162;
 wire net21163;
 wire net21164;
 wire net21166;
 wire net21167;
 wire net21168;
 wire net21169;
 wire net21170;
 wire net21171;
 wire net21172;
 wire net21173;
 wire net21174;
 wire net21175;
 wire net21176;
 wire net21260;
 wire net21177;
 wire net21178;
 wire net21180;
 wire net21181;
 wire net21182;
 wire net21183;
 wire net21184;
 wire net21185;
 wire net21186;
 wire net21187;
 wire net21188;
 wire net21189;
 wire net21190;
 wire net21191;
 wire net21227;
 wire net21192;
 wire net21193;
 wire net21194;
 wire net21195;
 wire net21196;
 wire net21197;
 wire net21198;
 wire net21199;
 wire net21200;
 wire net21201;
 wire net21202;
 wire net21203;
 wire net21211;
 wire net21204;
 wire net21213;
 wire net21205;
 wire net21206;
 wire net21207;
 wire net21208;
 wire net21209;
 wire net21210;
 wire net21212;
 wire net21264;
 wire net21214;
 wire net21215;
 wire net21216;
 wire net21217;
 wire net21218;
 wire net21219;
 wire net21220;
 wire net21221;
 wire net21222;
 wire net21223;
 wire net21224;
 wire net21225;
 wire net21533;
 wire net21226;
 wire net21228;
 wire net21229;
 wire net21230;
 wire net21231;
 wire net21232;
 wire net21233;
 wire net21234;
 wire net21235;
 wire net21236;
 wire net21237;
 wire net21238;
 wire net21293;
 wire net21404;
 wire net21239;
 wire net21240;
 wire net21241;
 wire net21242;
 wire net21267;
 wire net21243;
 wire net21245;
 wire net21246;
 wire net21247;
 wire net21248;
 wire net21259;
 wire net21250;
 wire net21251;
 wire net21252;
 wire net21253;
 wire net17410;
 wire net21254;
 wire net21255;
 wire net21256;
 wire net21257;
 wire net17408;
 wire net21258;
 wire net21261;
 wire net21262;
 wire net17403;
 wire net17429;
 wire net17409;
 wire net17394;
 wire net17336;
 wire net17337;
 wire net17334;
 wire net17333;
 wire net17328;
 wire net17327;
 wire net17325;
 wire clknet_leaf_25_clk;
 wire net17357;
 wire net17310;
 wire net17302;
 wire clknet_leaf_28_clk;
 wire net17298;
 wire net17295;
 wire net21322;
 wire net17506;
 wire net21311;
 wire net21286;
 wire net21276;
 wire net21287;
 wire net21263;
 wire net21270;
 wire net21265;
 wire net21268;
 wire net21269;
 wire net21280;
 wire net21271;
 wire net21274;
 wire net21273;
 wire net17503;
 wire net21363;
 wire net21282;
 wire net21277;
 wire net21375;
 wire net21278;
 wire net21281;
 wire net21279;
 wire net21299;
 wire net21283;
 wire net21300;
 wire net21284;
 wire net21541;
 wire net21285;
 wire net21296;
 wire net21288;
 wire net21302;
 wire net21289;
 wire net21540;
 wire net21290;
 wire net21303;
 wire net21292;
 wire net21291;
 wire net21353;
 wire net21295;
 wire net21297;
 wire net21298;
 wire net21301;
 wire net17501;
 wire net21348;
 wire net21537;
 wire net21345;
 wire net21307;
 wire net21304;
 wire net21318;
 wire net21310;
 wire net21342;
 wire net21312;
 wire net21314;
 wire net21315;
 wire net21316;
 wire net21319;
 wire net21317;
 wire net21320;
 wire net21334;
 wire net21331;
 wire net21328;
 wire net17314;
 wire net21321;
 wire net17313;
 wire net21536;
 wire net21325;
 wire net21324;
 wire net21326;
 wire net21327;
 wire net21329;
 wire net21330;
 wire net21333;
 wire net21332;
 wire net21493;
 wire net21340;
 wire net21335;
 wire net21356;
 wire net21336;
 wire net649;
 wire net21337;
 wire net17500;
 wire net21338;
 wire net21339;
 wire net17320;
 wire net21343;
 wire net21347;
 wire net21344;
 wire net21346;
 wire net21365;
 wire net21492;
 wire net21351;
 wire net21349;
 wire net17294;
 wire net21350;
 wire net17293;
 wire net17281;
 wire net21366;
 wire net21355;
 wire net21352;
 wire net21360;
 wire net21354;
 wire net21358;
 wire net21357;
 wire net21394;
 wire net21359;
 wire net21361;
 wire net21362;
 wire net21372;
 wire net21371;
 wire net17289;
 wire net21401;
 wire net21364;
 wire net21389;
 wire clknet_leaf_22_clk;
 wire net21380;
 wire net21374;
 wire net21403;
 wire net21368;
 wire net21367;
 wire net21370;
 wire net21369;
 wire net21402;
 wire net21373;
 wire net21385;
 wire net21381;
 wire net21376;
 wire clknet_leaf_21_clk;
 wire net21386;
 wire net21377;
 wire clknet_leaf_19_clk;
 wire net21378;
 wire clknet_leaf_5_clk;
 wire net21379;
 wire clknet_leaf_15_clk;
 wire net21411;
 wire net21382;
 wire net21395;
 wire net21383;
 wire net21388;
 wire net21384;
 wire net21387;
 wire net21390;
 wire net21391;
 wire net21392;
 wire net21466;
 wire net21393;
 wire net21396;
 wire net21399;
 wire net21397;
 wire net21398;
 wire net21400;
 wire net21491;
 wire clknet_leaf_29_clk;
 wire net21429;
 wire net21405;
 wire net21408;
 wire net21427;
 wire net21406;
 wire net21423;
 wire net21417;
 wire net21416;
 wire net21407;
 wire net21428;
 wire net21412;
 wire net21410;
 wire clknet_leaf_1_clk;
 wire net21436;
 wire net21415;
 wire net21420;
 wire net21430;
 wire net21419;
 wire clknet_leaf_11_clk;
 wire net21418;
 wire net21435;
 wire net21432;
 wire net21422;
 wire net21421;
 wire net21426;
 wire net21431;
 wire net21433;
 wire net21434;
 wire net21450;
 wire net21490;
 wire net21489;
 wire net21446;
 wire net21437;
 wire clknet_leaf_0_clk;
 wire net21438;
 wire net21445;
 wire clknet_leaf_7_clk;
 wire net21442;
 wire net21440;
 wire net21441;
 wire net17362;
 wire net21443;
 wire net17433;
 wire net21444;
 wire net21447;
 wire net21486;
 wire net21457;
 wire net21449;
 wire net21448;
 wire net21464;
 wire net21452;
 wire net21485;
 wire net21451;
 wire net21455;
 wire net21453;
 wire net21454;
 wire net21484;
 wire net21459;
 wire net21465;
 wire net21460;
 wire net17363;
 wire net21469;
 wire net21480;
 wire net21461;
 wire net17280;
 wire net17278;
 wire net17360;
 wire net21471;
 wire net21462;
 wire net21463;
 wire net21468;
 wire net21467;
 wire net21476;
 wire net21470;
 wire net17423;
 wire net21479;
 wire net21472;
 wire net21478;
 wire net21473;
 wire net21475;
 wire net21474;
 wire net17393;
 wire net17376;
 wire net17368;
 wire net17367;
 wire net17364;
 wire net21477;
 wire net21481;
 wire net17365;
 wire net21483;
 wire net21482;
 wire net21544;
 wire clknet_leaf_32_clk;
 wire net17487;
 wire net17513;
 wire net17407;
 wire net17432;
 wire net17321;
 wire net17200;
 wire net21539;
 wire net17249;
 wire net17275;
 wire net17225;
 wire net17273;
 wire net17319;
 wire net17318;
 wire net17245;
 wire net17247;
 wire net17271;
 wire net17265;
 wire net17323;
 wire net17322;
 wire net17269;
 wire net17268;
 wire net17324;
 wire net17331;
 wire net17326;
 wire net17210;
 wire net17316;
 wire net17251;
 wire net17218;
 wire net17223;
 wire net17208;
 wire net17204;
 wire net17224;
 wire net17279;
 wire net17221;
 wire net17274;
 wire net17272;
 wire net17199;
 wire net17267;
 wire net17260;
 wire net17258;
 wire net17257;
 wire net17214;
 wire net17256;
 wire net17211;
 wire net17202;
 wire net17286;
 wire net17240;
 wire net17226;
 wire net17263;
 wire net17212;
 wire net17254;
 wire net17231;
 wire net17207;
 wire net17217;
 wire net17213;
 wire net17209;
 wire net17222;
 wire net20714;
 wire net20710;
 wire net20715;
 wire net20707;
 wire net20704;
 wire net20703;
 wire net18306;
 wire net18827;
 wire net18826;
 wire net18790;
 wire net18789;
 wire net18307;
 wire net18456;
 wire net18471;
 wire net18477;
 wire net18480;
 wire net18513;
 wire net18515;
 wire net18516;
 wire net18519;
 wire net18521;
 wire net18520;
 wire net18525;
 wire net18533;
 wire net18532;
 wire net18599;
 wire net18598;
 wire net18557;
 wire net18556;
 wire net18555;
 wire net18554;
 wire net18553;
 wire net18552;
 wire net18551;
 wire net18550;
 wire net18549;
 wire net18821;
 wire net18811;
 wire net18812;
 wire net18859;
 wire net18858;
 wire net18857;
 wire net18856;
 wire net18855;
 wire net18835;
 wire net18832;
 wire net18922;
 wire net18921;
 wire net18249;
 wire net19157;
 wire net19158;
 wire net19159;
 wire net20461;
 wire net20462;
 wire net20463;
 wire net20464;
 wire net20465;
 wire net20466;
 wire net20467;
 wire net20468;
 wire net20469;
 wire net20589;
 wire net20590;
 wire net20591;
 wire net20592;
 wire net21083;
 wire net21084;
 wire net21085;
 wire net21086;
 wire net21087;
 wire net21088;
 wire net21089;
 wire net21090;
 wire net21091;
 wire net21092;
 wire net21093;
 wire net21094;
 wire net21095;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_349_clk;
 wire clknet_leaf_352_clk;
 wire clknet_leaf_354_clk;
 wire clknet_leaf_355_clk;
 wire clknet_leaf_358_clk;
 wire clknet_leaf_362_clk;
 wire clknet_leaf_363_clk;
 wire clknet_leaf_369_clk;
 wire clknet_leaf_370_clk;
 wire clknet_leaf_372_clk;
 wire clknet_leaf_376_clk;
 wire clknet_leaf_377_clk;
 wire clknet_leaf_378_clk;
 wire clknet_leaf_382_clk;
 wire clknet_leaf_385_clk;
 wire clknet_leaf_389_clk;
 wire clknet_leaf_390_clk;
 wire clknet_leaf_394_clk;
 wire clknet_leaf_399_clk;
 wire clknet_leaf_410_clk;
 wire clknet_leaf_411_clk;
 wire clknet_leaf_412_clk;
 wire clknet_leaf_413_clk;
 wire clknet_leaf_415_clk;
 wire clknet_leaf_417_clk;
 wire clknet_leaf_423_clk;
 wire clknet_leaf_424_clk;
 wire clknet_leaf_425_clk;
 wire clknet_leaf_431_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net526;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net427;
 wire net428;
 wire net430;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net462;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net471;
 wire net473;
 wire net474;
 wire net475;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net528;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net419;
 wire net423;
 wire net435;
 wire net436;
 wire net438;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net461;
 wire net463;
 wire net464;
 wire net470;
 wire net472;
 wire net476;
 wire net477;
 wire net478;
 wire net493;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net523;
 wire net524;
 wire net525;
 wire net529;
 wire net530;
 wire net603;
 wire net604;
 wire net605;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net630;
 wire net631;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net668;
 wire net669;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire [0:0] _15537_;
 wire [0:0] _15538_;
 wire [0:0] _15539_;
 wire [0:0] _15540_;
 wire [0:0] _15541_;
 wire [0:0] _15542_;
 wire [0:0] _15543_;
 wire [0:0] _15544_;
 wire [0:0] _15545_;
 wire [0:0] _15546_;
 wire [0:0] _15547_;
 wire [0:0] _15548_;
 wire [0:0] _15549_;
 wire [0:0] _15550_;
 wire [0:0] _15551_;
 wire [0:0] _15552_;
 wire [0:0] _15553_;
 wire [0:0] _15554_;
 wire [0:0] _15555_;
 wire [0:0] _15556_;
 wire [0:0] _15558_;
 wire [0:0] _15559_;
 wire [0:0] _15560_;
 wire [0:0] _15561_;
 wire [0:0] _15563_;
 wire [0:0] _15564_;
 wire [0:0] _15565_;
 wire [0:0] _15566_;
 wire [0:0] _15567_;
 wire [0:0] _15568_;
 wire [0:0] _15569_;
 wire [0:0] _15570_;
 wire [0:0] _15571_;
 wire [0:0] _15572_;
 wire [0:0] _15573_;
 wire [0:0] _15574_;
 wire [0:0] _15575_;
 wire [0:0] _15576_;
 wire [0:0] _15577_;
 wire [0:0] _15578_;
 wire [0:0] _15579_;
 wire [0:0] _15580_;
 wire [0:0] _15581_;
 wire [0:0] _15582_;
 wire [0:0] _15583_;
 wire [0:0] _15584_;
 wire [0:0] _15585_;
 wire [0:0] _15586_;
 wire [0:0] _15587_;
 wire [0:0] _15588_;
 wire [0:0] _15589_;
 wire [0:0] _15590_;
 wire [0:0] _15592_;
 wire [0:0] _15593_;
 wire [0:0] _15594_;
 wire [0:0] _15595_;
 wire [0:0] _15597_;
 wire [0:0] _15598_;
 wire [0:0] _15599_;
 wire [0:0] _15600_;
 wire [0:0] _15601_;
 wire [0:0] _15602_;
 wire [0:0] _15603_;
 wire [0:0] _15604_;
 wire [0:0] _15605_;
 wire [0:0] _15606_;
 wire [0:0] _15607_;
 wire [0:0] _15608_;
 wire [0:0] _15609_;
 wire [0:0] _15610_;
 wire [0:0] _15611_;
 wire [0:0] _15612_;
 wire [0:0] _15613_;
 wire [0:0] _15614_;
 wire [0:0] _15615_;
 wire [0:0] _15616_;
 wire [0:0] _15617_;
 wire [0:0] _15618_;
 wire [0:0] _15619_;
 wire [0:0] _15620_;
 wire [0:0] _15621_;
 wire [0:0] _15622_;
 wire [0:0] _15623_;
 wire [0:0] _15624_;
 wire [0:0] _15626_;
 wire [0:0] _15627_;
 wire [0:0] _15628_;
 wire [0:0] _15629_;
 wire [0:0] _15631_;
 wire [0:0] _15632_;
 wire [0:0] _15633_;
 wire [0:0] _15634_;
 wire [0:0] _15635_;
 wire [0:0] _15636_;
 wire [0:0] _15637_;
 wire [0:0] _15638_;
 wire [0:0] _15639_;
 wire [0:0] _15640_;
 wire [0:0] _15641_;
 wire [0:0] _15642_;
 wire [0:0] _15643_;
 wire [0:0] _15644_;
 wire [0:0] _15645_;
 wire [0:0] _15646_;
 wire [0:0] _15647_;
 wire [0:0] _15648_;
 wire [0:0] _15649_;
 wire [0:0] _15650_;
 wire [0:0] _15651_;
 wire [0:0] _15652_;
 wire [0:0] _15653_;
 wire [0:0] _15654_;
 wire [0:0] _15655_;
 wire [0:0] _15656_;
 wire [0:0] _15657_;
 wire [0:0] _15658_;
 wire [0:0] _15660_;
 wire [0:0] _15661_;
 wire [0:0] _15662_;
 wire [0:0] _15663_;
 wire [0:0] _15665_;
 wire [0:0] _15666_;
 wire [0:0] _15667_;
 wire [0:0] _15668_;
 wire [0:0] _15669_;
 wire [0:0] _15670_;
 wire [0:0] _15671_;
 wire [0:0] _15672_;
 wire [0:0] _15673_;
 wire [0:0] _15674_;
 wire [0:0] _15675_;
 wire [0:0] _15676_;
 wire [0:0] _15677_;
 wire [0:0] _15678_;
 wire [0:0] _15679_;
 wire [0:0] _15680_;
 wire [0:0] _15681_;
 wire [0:0] _15682_;
 wire [0:0] _15683_;
 wire [0:0] _15684_;
 wire [0:0] _15685_;
 wire [0:0] _15686_;
 wire [0:0] _15687_;
 wire [0:0] _15688_;
 wire [0:0] _15689_;
 wire [0:0] _15690_;
 wire [0:0] _15692_;
 wire [0:0] _15693_;
 wire [0:0] _15694_;
 wire [0:0] _15695_;
 wire [0:0] _15696_;
 wire [0:0] _15697_;
 wire [0:0] _15699_;
 wire [0:0] _15700_;
 wire [0:0] _15701_;
 wire [0:0] _15702_;
 wire [0:0] _15703_;
 wire [0:0] _15704_;
 wire [0:0] _15705_;
 wire [0:0] _15706_;
 wire [0:0] _15707_;
 wire [0:0] _15708_;
 wire [0:0] _15709_;
 wire [0:0] _15710_;
 wire [0:0] _15712_;
 wire [0:0] _15713_;
 wire [0:0] _15714_;
 wire [0:0] _15715_;
 wire [0:0] _15716_;
 wire [0:0] _15717_;
 wire [0:0] _15718_;
 wire [0:0] _15719_;
 wire [0:0] _15720_;
 wire [0:0] _15721_;
 wire [0:0] _15722_;
 wire [0:0] _15724_;
 wire [0:0] _15725_;
 wire [0:0] _15726_;
 wire [0:0] _15727_;
 wire [0:0] _15728_;
 wire [0:0] _15729_;
 wire [0:0] _15731_;
 wire [0:0] _15732_;
 wire [0:0] _15733_;
 wire [0:0] _15734_;
 wire [0:0] _15735_;
 wire [0:0] _15736_;
 wire [0:0] _15737_;
 wire [0:0] _15738_;
 wire [0:0] _15739_;
 wire [0:0] _15740_;
 wire [0:0] _15741_;
 wire [0:0] _15742_;
 wire [0:0] _15744_;
 wire [0:0] _15745_;
 wire [0:0] _15746_;
 wire [0:0] _15747_;
 wire [0:0] _15748_;
 wire [0:0] _15749_;
 wire [0:0] _15750_;
 wire [0:0] _15751_;
 wire [0:0] _15752_;
 wire [0:0] _15753_;
 wire [0:0] _15754_;
 wire [0:0] _15756_;
 wire [0:0] _15757_;
 wire [0:0] _15758_;
 wire [0:0] _15759_;
 wire [0:0] _15760_;
 wire [0:0] _15761_;
 wire [0:0] _15763_;
 wire [0:0] _15764_;
 wire [0:0] _15765_;
 wire [0:0] _15766_;
 wire [0:0] _15767_;
 wire [0:0] _15768_;
 wire [0:0] _15769_;
 wire [0:0] _15770_;
 wire [0:0] _15771_;
 wire [0:0] _15772_;
 wire [0:0] _15773_;
 wire [0:0] _15774_;
 wire [0:0] _15775_;
 wire [0:0] _15776_;
 wire [0:0] _15777_;
 wire [0:0] _15778_;
 wire [0:0] _15779_;
 wire [0:0] _15780_;
 wire [0:0] _15781_;
 wire [0:0] _15782_;
 wire [0:0] _15783_;
 wire [0:0] _15784_;
 wire [0:0] _15785_;
 wire [0:0] _15786_;
 wire [0:0] _15788_;
 wire [0:0] _15789_;
 wire [0:0] _15790_;
 wire [0:0] _15791_;
 wire [0:0] _15792_;
 wire [0:0] _15793_;
 wire [0:0] _15795_;
 wire [0:0] _15796_;
 wire [0:0] _15797_;
 wire [0:0] _15798_;
 wire [0:0] _15799_;
 wire [0:0] _15800_;
 wire [0:0] _15801_;
 wire [0:0] _15802_;
 wire [0:0] _15803_;
 wire [0:0] _15804_;
 wire [0:0] _15805_;
 wire [0:0] _15806_;
 wire [0:0] _15807_;
 wire [0:0] _15808_;
 wire [0:0] _15809_;
 wire [0:0] _15810_;
 wire [0:0] _15811_;
 wire [0:0] _15812_;
 wire [0:0] _15813_;
 wire [0:0] _15814_;
 wire [0:0] _15815_;
 wire [0:0] _15816_;
 wire [0:0] _15817_;
 wire [0:0] _15818_;
 wire [0:0] _15820_;
 wire [0:0] _15821_;
 wire [0:0] _15822_;
 wire [0:0] _15823_;
 wire [0:0] _15824_;
 wire [0:0] _15825_;
 wire [0:0] _15827_;
 wire [0:0] _15828_;
 wire [0:0] _15829_;
 wire [0:0] _15830_;
 wire [0:0] _15831_;
 wire [0:0] _15832_;
 wire [0:0] _15833_;
 wire [0:0] _15834_;
 wire [0:0] _15835_;
 wire [0:0] _15836_;
 wire [0:0] _15837_;
 wire [0:0] _15838_;
 wire [0:0] _15839_;
 wire [0:0] _15840_;
 wire [0:0] _15841_;
 wire [0:0] _15842_;
 wire [0:0] _15843_;
 wire [0:0] _15844_;
 wire [0:0] _15845_;
 wire [0:0] _15846_;
 wire [0:0] _15847_;
 wire [0:0] _15848_;
 wire [0:0] _15849_;
 wire [0:0] _15850_;
 wire [0:0] _15852_;
 wire [0:0] _15853_;
 wire [0:0] _15854_;
 wire [0:0] _15855_;
 wire [0:0] _15856_;
 wire [0:0] _15857_;
 wire [0:0] _15859_;
 wire [0:0] _15860_;
 wire [0:0] _15861_;
 wire [0:0] _15862_;
 wire [0:0] _15863_;
 wire [0:0] _15864_;
 wire [0:0] _15865_;
 wire [0:0] _15866_;
 wire [0:0] _15867_;
 wire [0:0] _15868_;
 wire [0:0] _15869_;
 wire [0:0] _15870_;
 wire [0:0] _15871_;
 wire [0:0] _15872_;
 wire [0:0] _15873_;
 wire [0:0] _15874_;
 wire [0:0] _15875_;
 wire [0:0] _15876_;
 wire [0:0] _15877_;
 wire [0:0] _15878_;
 wire [0:0] _15879_;
 wire [0:0] _15880_;
 wire [0:0] _15881_;
 wire [0:0] _15882_;
 wire [0:0] _15884_;
 wire [0:0] _15885_;
 wire [0:0] _15886_;
 wire [0:0] _15887_;
 wire [0:0] _15888_;
 wire [0:0] _15889_;
 wire [0:0] _15891_;
 wire [0:0] _15892_;
 wire [0:0] _15893_;
 wire [0:0] _15894_;
 wire [0:0] _15895_;
 wire [0:0] _15896_;
 wire [0:0] _15897_;
 wire [0:0] _15898_;
 wire [0:0] _15899_;
 wire [0:0] _15900_;
 wire [0:0] _15901_;
 wire [0:0] _15902_;
 wire [0:0] _15903_;
 wire [0:0] _15904_;
 wire [0:0] _15905_;
 wire [0:0] _15906_;
 wire [0:0] _15907_;
 wire [0:0] _15908_;
 wire [0:0] _15909_;
 wire [0:0] _15910_;
 wire [0:0] _15911_;
 wire [0:0] _15912_;
 wire [0:0] _15913_;
 wire [0:0] _15914_;
 wire [0:0] _15916_;
 wire [0:0] _15917_;
 wire [0:0] _15918_;
 wire [0:0] _15919_;
 wire [0:0] _15920_;
 wire [0:0] _15921_;
 wire [0:0] _15923_;
 wire [0:0] _15924_;
 wire [0:0] _15925_;
 wire [0:0] _15926_;
 wire [0:0] _15927_;
 wire [0:0] _15928_;
 wire [0:0] _15929_;
 wire [0:0] _15930_;
 wire [0:0] _15931_;
 wire [0:0] _15932_;
 wire [0:0] _15933_;
 wire [0:0] _15934_;
 wire [0:0] _15935_;
 wire [0:0] _15936_;
 wire [0:0] _15937_;
 wire [0:0] _15938_;
 wire [0:0] _15939_;
 wire [0:0] _15940_;
 wire [0:0] _15941_;
 wire [0:0] _15942_;
 wire [0:0] _15943_;
 wire [0:0] _15944_;
 wire [0:0] _15945_;
 wire [0:0] _15946_;
 wire [0:0] _15947_;
 wire [0:0] _15948_;
 wire [0:0] _15950_;
 wire [0:0] _15951_;
 wire [0:0] _15952_;
 wire [0:0] _15953_;
 wire [0:0] _15954_;
 wire [0:0] _15955_;
 wire [0:0] _15957_;
 wire [0:0] _15958_;
 wire [0:0] _15959_;
 wire [0:0] _15960_;
 wire [0:0] _15961_;
 wire [0:0] _15962_;
 wire [0:0] _15963_;
 wire [0:0] _15964_;
 wire [0:0] _15965_;
 wire [0:0] _15966_;
 wire [0:0] _15967_;
 wire [0:0] _15968_;
 wire [0:0] _15969_;
 wire [0:0] _15970_;
 wire [0:0] _15971_;
 wire [0:0] _15972_;
 wire [0:0] _15973_;
 wire [0:0] _15974_;
 wire [0:0] _15975_;
 wire [0:0] _15976_;
 wire [0:0] _15977_;
 wire [0:0] _15978_;
 wire [0:0] _15979_;
 wire [0:0] _15980_;
 wire [0:0] _15981_;
 wire [0:0] _15982_;
 wire [0:0] _15983_;
 wire [0:0] _15984_;
 wire [0:0] _15986_;
 wire [0:0] _15987_;
 wire [0:0] _15988_;
 wire [0:0] _15989_;
 wire [0:0] _15990_;
 wire [0:0] _15991_;
 wire [0:0] _15993_;
 wire [0:0] _15994_;
 wire [0:0] _15995_;
 wire [0:0] _15996_;
 wire [0:0] _15997_;
 wire [0:0] _15998_;
 wire [0:0] _15999_;
 wire [0:0] _16000_;
 wire [0:0] _16001_;
 wire [0:0] _16002_;
 wire [0:0] _16003_;
 wire [0:0] _16004_;
 wire [0:0] _16005_;
 wire [0:0] _16006_;
 wire [0:0] _16007_;
 wire [0:0] _16008_;
 wire [0:0] _16009_;
 wire [0:0] _16010_;
 wire [0:0] _16011_;
 wire [0:0] _16012_;
 wire [0:0] _16013_;
 wire [0:0] _16014_;
 wire [0:0] _16015_;
 wire [0:0] _16016_;
 wire [0:0] _16017_;
 wire [0:0] _16018_;
 wire [0:0] _16019_;
 wire [0:0] _16020_;
 wire [0:0] _16022_;
 wire [0:0] _16023_;
 wire [0:0] _16024_;
 wire [0:0] _16025_;
 wire [0:0] _16026_;
 wire [0:0] _16027_;
 wire [0:0] _16029_;
 wire [0:0] _16030_;
 wire [0:0] _16031_;
 wire [0:0] _16032_;
 wire [0:0] _16033_;
 wire [0:0] _16034_;
 wire [0:0] _16035_;
 wire [0:0] _16036_;
 wire [0:0] _16037_;
 wire [0:0] _16038_;
 wire [0:0] _16039_;
 wire [0:0] _16040_;
 wire [0:0] _16041_;
 wire [0:0] _16042_;
 wire [0:0] _16043_;
 wire [0:0] _16044_;
 wire [0:0] _16045_;
 wire [0:0] _16046_;
 wire [0:0] _16047_;
 wire [0:0] _16048_;
 wire [0:0] _16049_;
 wire [0:0] _16050_;
 wire [0:0] _16051_;
 wire [0:0] _16052_;
 wire [0:0] _16053_;
 wire [0:0] _16054_;
 wire [0:0] _16055_;
 wire [0:0] _16056_;
 wire [0:0] _16058_;
 wire [0:0] _16059_;
 wire [0:0] _16060_;
 wire [0:0] _16061_;
 wire [0:0] _16062_;
 wire [0:0] _16063_;
 wire [0:0] _16065_;
 wire [0:0] _16066_;
 wire [0:0] _16067_;
 wire [0:0] _16068_;
 wire [0:0] _16069_;
 wire [0:0] _16070_;
 wire [0:0] _16071_;
 wire [0:0] _16072_;
 wire [0:0] _16074_;
 wire [0:0] _16075_;
 wire [0:0] _16076_;
 wire [0:0] _16077_;
 wire [0:0] _16078_;
 wire [0:0] _16079_;
 wire [0:0] _16080_;
 wire [0:0] _16081_;
 wire [0:0] _16082_;
 wire [0:0] _16083_;
 wire [0:0] _16084_;
 wire [0:0] _16085_;
 wire [0:0] _16086_;
 wire [0:0] _16087_;
 wire [0:0] _16088_;
 wire [0:0] _16089_;
 wire [0:0] _16090_;
 wire [0:0] _16092_;
 wire [0:0] _16093_;
 wire [0:0] _16094_;
 wire [0:0] _16095_;
 wire [0:0] _16096_;
 wire [0:0] _16097_;
 wire [0:0] _16099_;
 wire [0:0] _16100_;
 wire [0:0] _16101_;
 wire [0:0] _16102_;
 wire [0:0] _16103_;
 wire [0:0] _16104_;
 wire [0:0] _16105_;
 wire [0:0] _16106_;
 wire [0:0] _16107_;
 wire [0:0] _16108_;
 wire [0:0] _16109_;
 wire [0:0] _16110_;
 wire [0:0] _16111_;
 wire [0:0] _16112_;
 wire [0:0] _16113_;
 wire [0:0] _16114_;
 wire [0:0] _16115_;
 wire [0:0] _16116_;
 wire [0:0] _16117_;
 wire [0:0] _16118_;
 wire [0:0] _16119_;
 wire [0:0] _16120_;
 wire [0:0] _16121_;
 wire [0:0] _16122_;
 wire [0:0] _16124_;
 wire [0:0] _16125_;
 wire [0:0] _16126_;
 wire [0:0] _16127_;
 wire [0:0] _16128_;
 wire [0:0] _16129_;
 wire [0:0] _16131_;
 wire [0:0] _16132_;
 wire [0:0] _16133_;
 wire [0:0] _16134_;
 wire [0:0] _16135_;
 wire [0:0] _16136_;
 wire [0:0] _16137_;
 wire [0:0] _16138_;
 wire [0:0] _16139_;
 wire [0:0] _16140_;
 wire [0:0] _16141_;
 wire [0:0] _16142_;
 wire [0:0] _16144_;
 wire [0:0] _16145_;
 wire [0:0] _16146_;
 wire [0:0] _16147_;
 wire [0:0] _16148_;
 wire [0:0] _16149_;
 wire [0:0] _16150_;
 wire [0:0] _16151_;
 wire [0:0] _16152_;
 wire [0:0] _16153_;
 wire [0:0] _16154_;
 wire [0:0] _16156_;
 wire [0:0] _16157_;
 wire [0:0] _16158_;
 wire [0:0] _16159_;
 wire [0:0] _16160_;
 wire [0:0] _16161_;
 wire [0:0] _16163_;
 wire [0:0] _16164_;
 wire [0:0] _16165_;
 wire [0:0] _16166_;
 wire [0:0] _16167_;
 wire [0:0] _16168_;
 wire [0:0] _16169_;
 wire [0:0] _16170_;
 wire [0:0] _16171_;
 wire [0:0] _16172_;
 wire [0:0] _16173_;
 wire [0:0] _16174_;
 wire [0:0] _16176_;
 wire [0:0] _16177_;
 wire [0:0] _16178_;
 wire [0:0] _16179_;
 wire [0:0] _16180_;
 wire [0:0] _16181_;
 wire [0:0] _16182_;
 wire [0:0] _16183_;
 wire [0:0] _16184_;
 wire [0:0] _16185_;
 wire [0:0] _16186_;
 wire [0:0] _16188_;
 wire [0:0] _16189_;
 wire [0:0] _16190_;
 wire [0:0] _16191_;
 wire [0:0] _16192_;
 wire [0:0] _16193_;
 wire [0:0] _16195_;
 wire [0:0] _16196_;
 wire [0:0] _16197_;
 wire [0:0] _16198_;
 wire [0:0] _16199_;
 wire [0:0] _16200_;
 wire [0:0] _16201_;
 wire [0:0] _16202_;
 wire [0:0] _16203_;
 wire [0:0] _16204_;
 wire [0:0] _16205_;
 wire [0:0] _16206_;
 wire [0:0] _16207_;
 wire [0:0] _16208_;
 wire [0:0] _16209_;
 wire [0:0] _16210_;

 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16211_ (.A1(\u0.w[0][19] ),
    .A2(\u0.w[2][19] ),
    .ZN(_07232_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16212_ (.A1(\u0.w[1][19] ),
    .A2(\u0.subword[19] ),
    .Z(_07243_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16213_ (.A1(\u0.tmp_w[19] ),
    .A2(_07243_),
    .Z(_07254_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16214_ (.A1(_07232_),
    .A2(_07254_),
    .Z(_07265_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16215_ (.I(net129),
    .ZN(_07276_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17768 (.I(_01805_),
    .Z(net17768));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16217_ (.A1(_07265_),
    .A2(net21518),
    .ZN(_07297_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16218_ (.A1(net21530),
    .A2(net39),
    .Z(_07308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16219_ (.A1(_07297_),
    .A2(_07308_),
    .ZN(_07319_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _16220_ (.I(_07319_),
    .ZN(_07330_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17800 (.I(_01076_),
    .Z(net17800));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17777 (.I(_01753_),
    .Z(net17777));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16223_ (.A1(\u0.w[0][16] ),
    .A2(\u0.w[2][16] ),
    .ZN(_07361_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16224_ (.A1(\u0.w[1][16] ),
    .A2(\u0.subword[16] ),
    .Z(_07372_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16225_ (.A1(_07372_),
    .A2(\u0.tmp_w[16] ),
    .Z(_07383_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16226_ (.A1(_07383_),
    .A2(_07361_),
    .Z(_07394_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17769 (.I(_01799_),
    .Z(net17769));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16228_ (.A1(_07394_),
    .A2(net21530),
    .ZN(_07415_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16229_ (.I(net36),
    .ZN(_07426_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17803 (.I(_01046_),
    .Z(net17803));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16231_ (.A1(_07426_),
    .A2(net21542),
    .Z(_07448_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16232_ (.I(net21133),
    .ZN(_07458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16233_ (.A1(_07415_),
    .A2(_07458_),
    .ZN(_15543_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16234_ (.A1(\u0.w[0][17] ),
    .A2(\u0.w[2][17] ),
    .ZN(_07463_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16235_ (.A1(\u0.w[1][17] ),
    .A2(\u0.subword[17] ),
    .Z(_07464_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16236_ (.A1(\u0.tmp_w[17] ),
    .A2(_07464_),
    .Z(_07465_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16237_ (.A1(_07463_),
    .A2(_07465_),
    .Z(_07466_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17775 (.I(_01775_),
    .Z(net17775));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17785 (.I(net17784),
    .Z(net17785));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16240_ (.A1(_07466_),
    .A2(net21530),
    .ZN(_07469_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16241_ (.I(net37),
    .ZN(_07470_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16242_ (.A1(_07470_),
    .A2(net21542),
    .Z(_07471_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16243_ (.I(_07471_),
    .ZN(_07472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16244_ (.A1(_07469_),
    .A2(_07472_),
    .ZN(_15548_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16245_ (.A1(\u0.w[0][21] ),
    .A2(\u0.w[2][21] ),
    .ZN(_07473_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16246_ (.A1(\u0.w[1][21] ),
    .A2(\u0.subword[21] ),
    .Z(_07475_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16247_ (.A1(\u0.tmp_w[21] ),
    .A2(_07475_),
    .Z(_07477_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16248_ (.A1(_07473_),
    .A2(_07477_),
    .Z(_07479_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16249_ (.A1(_07479_),
    .A2(net21530),
    .Z(_07481_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16250_ (.A1(net21530),
    .A2(net42),
    .ZN(_07482_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16251_ (.A1(_07481_),
    .A2(_07482_),
    .ZN(_07484_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17790 (.I(_01253_),
    .Z(net17790));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17793 (.I(_01232_),
    .Z(net17793));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16254_ (.A1(\u0.w[0][20] ),
    .A2(\u0.w[2][20] ),
    .ZN(_07489_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16255_ (.A1(\u0.w[1][20] ),
    .A2(\u0.subword[20] ),
    .Z(_07491_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16256_ (.A1(\u0.tmp_w[20] ),
    .A2(_07491_),
    .Z(_07493_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16257_ (.A1(_07489_),
    .A2(_07493_),
    .Z(_07495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16258_ (.A1(_07495_),
    .A2(net21530),
    .Z(_07497_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16259_ (.I(net41),
    .ZN(_07498_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16260_ (.A1(_07498_),
    .A2(net21544),
    .Z(_07504_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16261_ (.A1(_07497_),
    .A2(_07504_),
    .ZN(_07513_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17792 (.I(_01243_),
    .Z(net17792));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16263_ (.A1(\u0.w[0][18] ),
    .A2(\u0.w[2][18] ),
    .Z(_07526_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16264_ (.A1(\u0.subword[18] ),
    .A2(\u0.w[1][18] ),
    .Z(_07531_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16265_ (.A1(\u0.tmp_w[18] ),
    .A2(_07531_),
    .Z(_07532_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16266_ (.A1(_07526_),
    .A2(_07532_),
    .Z(_07533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16267_ (.A1(_07533_),
    .A2(net21530),
    .ZN(_07534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16268_ (.A1(net21544),
    .A2(net38),
    .ZN(_07535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16269_ (.A1(_07534_),
    .A2(_07535_),
    .ZN(_07536_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17748 (.I(_02535_),
    .Z(net17748));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17755 (.I(_02472_),
    .Z(net17755));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16272_ (.A1(\u0.w[0][0] ),
    .A2(\u0.w[2][0] ),
    .ZN(_07538_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16273_ (.A1(\u0.w[1][0] ),
    .A2(\u0.subword[0] ),
    .Z(_07539_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16274_ (.A1(\u0.tmp_w[0] ),
    .A2(_07539_),
    .Z(_07540_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16275_ (.A1(_07538_),
    .A2(_07540_),
    .Z(_07541_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17751 (.I(_02525_),
    .Z(net17751));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16277_ (.A1(net20923),
    .A2(net21527),
    .ZN(_07543_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16278_ (.I(net1),
    .ZN(_07544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16279_ (.A1(_07544_),
    .A2(net21531),
    .Z(_07545_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16280_ (.I(_07545_),
    .ZN(_07546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16281_ (.A1(_07546_),
    .A2(_07543_),
    .ZN(_15611_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16282_ (.A1(\u0.w[0][1] ),
    .A2(\u0.w[2][1] ),
    .ZN(_07547_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16283_ (.A1(\u0.w[1][1] ),
    .A2(\u0.subword[1] ),
    .Z(_07548_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16284_ (.A1(\u0.tmp_w[1] ),
    .A2(_07548_),
    .Z(_07549_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16285_ (.A1(_07549_),
    .A2(_07547_),
    .Z(_07550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16286_ (.A1(_07550_),
    .A2(net21527),
    .ZN(_07551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16287_ (.I(net40),
    .ZN(_07552_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16288_ (.A1(_07552_),
    .A2(net21531),
    .Z(_07553_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16289_ (.I(_07553_),
    .ZN(_07554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16290_ (.A1(_07554_),
    .A2(_07551_),
    .ZN(_15616_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16291_ (.A1(\u0.w[0][2] ),
    .A2(\u0.w[2][2] ),
    .ZN(_07555_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16292_ (.I(\u0.tmp_w[2] ),
    .ZN(_07556_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16293_ (.A1(\u0.subword[2] ),
    .A2(\u0.w[1][2] ),
    .Z(_07557_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16294_ (.A1(_07556_),
    .A2(_07557_),
    .Z(_07558_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16295_ (.A1(_07555_),
    .A2(_07558_),
    .Z(_07559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16296_ (.A1(_07559_),
    .A2(net21526),
    .ZN(_07560_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16297_ (.A1(net21533),
    .A2(net51),
    .Z(_07561_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16298_ (.I(_07561_),
    .ZN(_07562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16299_ (.A1(_07560_),
    .A2(_07562_),
    .ZN(_07563_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17745 (.I(_02585_),
    .Z(net17745));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16301_ (.A1(\u0.w[0][3] ),
    .A2(\u0.w[2][3] ),
    .ZN(_07564_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16302_ (.A1(\u0.w[1][3] ),
    .A2(\u0.subword[3] ),
    .Z(_07565_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16303_ (.A1(\u0.tmp_w[3] ),
    .A2(_07565_),
    .Z(_07566_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16304_ (.A1(_07564_),
    .A2(_07566_),
    .Z(_07567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16305_ (.A1(_07567_),
    .A2(net21518),
    .ZN(_07568_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16306_ (.A1(net21518),
    .A2(net62),
    .Z(_07569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16307_ (.A1(_07568_),
    .A2(_07569_),
    .ZN(_07570_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _16308_ (.I(_07570_),
    .ZN(_07571_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17744 (.I(_02597_),
    .Z(net17744));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17794 (.I(_01232_),
    .Z(net17794));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16311_ (.A1(\u0.w[0][4] ),
    .A2(\u0.w[2][4] ),
    .ZN(_07573_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16312_ (.A1(\u0.w[1][4] ),
    .A2(\u0.subword[4] ),
    .Z(_07574_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16313_ (.A1(\u0.tmp_w[4] ),
    .A2(_07574_),
    .Z(_07575_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16314_ (.A1(_07573_),
    .A2(_07575_),
    .Z(_07576_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16315_ (.A1(net21523),
    .A2(net73),
    .ZN(_07577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16316_ (.A1(_07576_),
    .A2(net21523),
    .B(_07577_),
    .ZN(_07578_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17747 (.I(_02573_),
    .Z(net17747));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17758 (.I(_02425_),
    .Z(net17758));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16319_ (.A1(\u0.w[0][5] ),
    .A2(\u0.w[2][5] ),
    .ZN(_07580_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16320_ (.A1(\u0.w[1][5] ),
    .A2(\u0.subword[5] ),
    .Z(_07581_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16321_ (.A1(\u0.tmp_w[5] ),
    .A2(_07581_),
    .Z(_07582_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16322_ (.A1(_07580_),
    .A2(_07582_),
    .Z(_07583_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16323_ (.A1(_07583_),
    .A2(net21520),
    .Z(_07584_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16324_ (.A1(net21520),
    .A2(net84),
    .ZN(_07585_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16325_ (.A1(_07584_),
    .A2(_07585_),
    .ZN(_07586_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17739 (.I(_02699_),
    .Z(net17739));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16327_ (.A1(\u0.w[1][6] ),
    .A2(\u0.subword[6] ),
    .Z(_07587_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16328_ (.A1(\u0.w[0][6] ),
    .A2(\u0.w[2][6] ),
    .ZN(_07588_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16329_ (.A1(\u0.tmp_w[6] ),
    .A2(_07587_),
    .A3(_07588_),
    .Z(_07589_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16330_ (.A1(_07589_),
    .A2(net21525),
    .Z(_07590_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16331_ (.A1(net21525),
    .A2(net95),
    .ZN(_07591_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16332_ (.A1(_07590_),
    .A2(_07591_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16333_ (.A1(\u0.w[1][7] ),
    .A2(\u0.subword[7] ),
    .Z(_07592_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16334_ (.A1(\u0.w[0][7] ),
    .A2(\u0.w[2][7] ),
    .ZN(_07593_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16335_ (.A1(\u0.tmp_w[7] ),
    .A2(_07592_),
    .A3(_07593_),
    .Z(_07594_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16336_ (.A1(_07594_),
    .A2(net21525),
    .Z(_07595_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17757 (.I(_02425_),
    .Z(net17757));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16338_ (.A1(net21525),
    .A2(net106),
    .ZN(_07597_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16339_ (.A1(_07595_),
    .A2(_07597_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16340_ (.A1(\u0.w[0][8] ),
    .A2(\u0.w[2][8] ),
    .ZN(_07598_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16341_ (.A1(\u0.w[1][8] ),
    .A2(\u0.subword[8] ),
    .Z(_07599_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16342_ (.A1(\u0.tmp_w[8] ),
    .A2(_07599_),
    .Z(_07600_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16343_ (.A1(_07598_),
    .A2(_07600_),
    .Z(_07601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16344_ (.A1(_07601_),
    .A2(net21518),
    .ZN(_07602_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16345_ (.I(net117),
    .ZN(_07603_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16346_ (.A1(_07603_),
    .A2(net21531),
    .Z(_07604_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16347_ (.I(net21120),
    .ZN(_07605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16348_ (.A1(_07602_),
    .A2(_07605_),
    .ZN(_15577_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16349_ (.A1(\u0.w[0][9] ),
    .A2(\u0.w[2][9] ),
    .ZN(_07606_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16350_ (.A1(\u0.w[1][9] ),
    .A2(\u0.subword[9] ),
    .Z(_07607_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16351_ (.A1(\u0.tmp_w[9] ),
    .A2(_07607_),
    .Z(_07608_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16352_ (.A1(_07608_),
    .A2(_07606_),
    .Z(_07609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16353_ (.A1(_07609_),
    .A2(net21518),
    .ZN(_07610_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16354_ (.I(net128),
    .ZN(_07611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16355_ (.A1(_07611_),
    .A2(net21542),
    .Z(_07612_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16356_ (.I(_07612_),
    .ZN(_07613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16357_ (.A1(_07613_),
    .A2(_07610_),
    .ZN(_15582_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16358_ (.A1(\u0.w[0][10] ),
    .A2(\u0.w[2][10] ),
    .ZN(_07614_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16359_ (.I(\u0.tmp_w[10] ),
    .ZN(_07615_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16360_ (.A1(\u0.subword[10] ),
    .A2(\u0.w[1][10] ),
    .Z(_07616_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16361_ (.A1(_07615_),
    .A2(_07616_),
    .Z(_07617_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16362_ (.A1(_07614_),
    .A2(_07617_),
    .Z(_07618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16363_ (.A1(_07618_),
    .A2(net21524),
    .ZN(_07619_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16364_ (.A1(net21543),
    .A2(net12),
    .Z(_07620_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16365_ (.I(_07620_),
    .ZN(_07621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16366_ (.A1(_07619_),
    .A2(_07621_),
    .ZN(_07622_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17736 (.I(_02939_),
    .Z(net17736));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16368_ (.A1(\u0.w[0][11] ),
    .A2(\u0.w[2][11] ),
    .ZN(_07623_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16369_ (.A1(\u0.w[1][11] ),
    .A2(\u0.subword[11] ),
    .Z(_07624_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16370_ (.A1(\u0.tmp_w[11] ),
    .A2(_07624_),
    .Z(_07625_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16371_ (.A1(_07623_),
    .A2(_07625_),
    .Z(_07626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16372_ (.A1(_07626_),
    .A2(net21518),
    .ZN(_07627_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16373_ (.A1(net21518),
    .A2(net23),
    .Z(_07628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16374_ (.A1(_07627_),
    .A2(_07628_),
    .ZN(_07629_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _16375_ (.I(_07629_),
    .ZN(_07630_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17754 (.I(net17753),
    .Z(net17754));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17762 (.I(net444),
    .Z(net17762));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16378_ (.A1(\u0.w[0][12] ),
    .A2(\u0.w[2][12] ),
    .ZN(_07632_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16379_ (.A1(\u0.w[1][12] ),
    .A2(\u0.subword[12] ),
    .Z(_07633_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16380_ (.A1(\u0.tmp_w[12] ),
    .A2(_07633_),
    .Z(_07634_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16381_ (.A1(_07632_),
    .A2(_07634_),
    .Z(_07635_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16382_ (.I(net32),
    .ZN(_07636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16383_ (.I0(_07635_),
    .I1(_07636_),
    .S(net21532),
    .Z(_07637_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17734 (.I(_03201_),
    .Z(net17734));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _16385_ (.I(_07637_),
    .ZN(_07639_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17733 (.I(_03223_),
    .Z(net17733));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17731 (.I(_03229_),
    .Z(net17731));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16388_ (.A1(\u0.w[0][13] ),
    .A2(\u0.w[2][13] ),
    .ZN(_07641_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16389_ (.A1(\u0.w[1][13] ),
    .A2(\u0.subword[13] ),
    .Z(_07642_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16390_ (.A1(\u0.tmp_w[13] ),
    .A2(_07642_),
    .Z(_07643_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16391_ (.A1(_07641_),
    .A2(_07643_),
    .Z(_07644_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16392_ (.A1(_07644_),
    .A2(net21523),
    .Z(_07645_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16393_ (.A1(net21523),
    .A2(net33),
    .ZN(_07646_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16394_ (.A1(_07645_),
    .A2(_07646_),
    .ZN(_07647_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17735 (.I(_03147_),
    .Z(net17735));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16396_ (.A1(\u0.w[0][14] ),
    .A2(\u0.w[2][14] ),
    .ZN(_07648_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16397_ (.A1(\u0.w[1][14] ),
    .A2(\u0.subword[14] ),
    .Z(_07649_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16398_ (.A1(\u0.tmp_w[14] ),
    .A2(_07649_),
    .Z(_07650_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16399_ (.A1(_07648_),
    .A2(_07650_),
    .Z(_07651_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16400_ (.A1(_07651_),
    .A2(net21521),
    .Z(_07652_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16401_ (.A1(net21521),
    .A2(net34),
    .ZN(_07653_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16402_ (.A1(_07652_),
    .A2(_07653_),
    .ZN(_07654_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17737 (.I(_02788_),
    .Z(net17737));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16404_ (.A1(\u0.w[1][15] ),
    .A2(\u0.subword[15] ),
    .Z(_07655_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16405_ (.A1(\u0.w[0][15] ),
    .A2(\u0.w[2][15] ),
    .ZN(_07656_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16406_ (.A1(\u0.tmp_w[15] ),
    .A2(_07655_),
    .A3(_07656_),
    .Z(_07657_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16407_ (.A1(_07657_),
    .A2(net21521),
    .Z(_07658_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16408_ (.A1(net21521),
    .A2(net35),
    .ZN(_07659_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16409_ (.A1(_07658_),
    .A2(_07659_),
    .ZN(_07660_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17732 (.I(_03229_),
    .Z(net17732));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16411_ (.A1(\u0.w[1][22] ),
    .A2(\u0.subword[22] ),
    .Z(_07661_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16412_ (.A1(\u0.w[0][22] ),
    .A2(\u0.w[2][22] ),
    .ZN(_07662_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16413_ (.A1(\u0.tmp_w[22] ),
    .A2(_07661_),
    .A3(_07662_),
    .Z(_07663_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16414_ (.A1(_07663_),
    .A2(net21530),
    .Z(_07664_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16415_ (.A1(net21530),
    .A2(net43),
    .ZN(_07665_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16416_ (.A1(_07664_),
    .A2(_07665_),
    .ZN(_07666_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17727 (.I(_03282_),
    .Z(net17727));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16418_ (.A1(\u0.w[1][23] ),
    .A2(\u0.subword[23] ),
    .Z(_07667_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16419_ (.A1(\u0.w[0][23] ),
    .A2(\u0.w[2][23] ),
    .ZN(_07668_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16420_ (.A1(\u0.tmp_w[23] ),
    .A2(_07667_),
    .A3(_07668_),
    .Z(_07669_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16421_ (.A1(_07669_),
    .A2(net21521),
    .Z(_07670_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16422_ (.A1(net21530),
    .A2(net44),
    .ZN(_07671_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16423_ (.A1(_07670_),
    .A2(_07671_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16424_ (.I(\u0.w[0][24] ),
    .ZN(_07672_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16425_ (.A1(\u0.w[2][24] ),
    .A2(\u0.r0.out[24] ),
    .Z(_07673_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16426_ (.A1(_07673_),
    .A2(_07672_),
    .Z(_07674_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16427_ (.A1(\u0.subword[24] ),
    .A2(\u0.w[1][24] ),
    .Z(_07675_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16428_ (.A1(\u0.tmp_w[24] ),
    .A2(_07675_),
    .Z(_07676_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16429_ (.A1(_07676_),
    .A2(_07674_),
    .Z(_07677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16430_ (.A1(_07674_),
    .A2(_07676_),
    .ZN(_07678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16431_ (.A1(_07678_),
    .A2(_07677_),
    .ZN(_07679_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16432_ (.A1(net21531),
    .A2(net45),
    .Z(_07680_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16433_ (.A1(net21526),
    .A2(net20844),
    .B(_07680_),
    .ZN(_15645_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16434_ (.A1(\u0.w[0][25] ),
    .A2(\u0.w[2][25] ),
    .Z(_07681_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16435_ (.A1(_07681_),
    .A2(\u0.r0.out[25] ),
    .Z(_07682_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16436_ (.A1(\u0.tmp_w[25] ),
    .A2(\u0.w[1][25] ),
    .Z(_07683_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16437_ (.A1(\u0.subword[25] ),
    .A2(_07683_),
    .Z(_07684_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16438_ (.A1(_07682_),
    .A2(_07684_),
    .Z(_07685_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16439_ (.A1(_07682_),
    .A2(_07684_),
    .ZN(_07686_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16440_ (.A1(_07685_),
    .A2(_07686_),
    .B(_07276_),
    .ZN(_07687_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16441_ (.A1(_07276_),
    .A2(net46),
    .Z(_07688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16442_ (.A1(_07687_),
    .A2(_07688_),
    .ZN(_15650_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16443_ (.I(\u0.w[0][26] ),
    .ZN(_07689_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16444_ (.A1(\u0.w[2][26] ),
    .A2(\u0.r0.out[26] ),
    .Z(_07690_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16445_ (.A1(_07689_),
    .A2(_07690_),
    .Z(_07691_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16446_ (.A1(\u0.w[1][26] ),
    .A2(\u0.subword[26] ),
    .Z(_07692_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16447_ (.A1(\u0.tmp_w[26] ),
    .A2(_07692_),
    .Z(_07693_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16448_ (.A1(_07691_),
    .A2(_07693_),
    .Z(_07694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16449_ (.A1(_07694_),
    .A2(net21529),
    .ZN(_07695_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16450_ (.A1(net21529),
    .A2(net47),
    .Z(_07696_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16451_ (.A1(_07695_),
    .A2(_07696_),
    .ZN(_07697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17808 (.I(_01020_),
    .Z(net17808));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16453_ (.A1(\u0.w[0][27] ),
    .A2(\u0.w[2][27] ),
    .Z(_07698_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16454_ (.A1(\u0.r0.out[27] ),
    .A2(_07698_),
    .Z(_07699_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16455_ (.A1(\u0.tmp_w[27] ),
    .A2(\u0.w[1][27] ),
    .Z(_07700_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16456_ (.A1(\u0.subword[27] ),
    .A2(_07700_),
    .Z(_07701_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16457_ (.A1(_07699_),
    .A2(_07701_),
    .Z(_07702_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16458_ (.A1(_07699_),
    .A2(_07701_),
    .ZN(_07703_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16459_ (.A1(_07702_),
    .A2(net21540),
    .A3(_07703_),
    .Z(_07704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16460_ (.A1(net21540),
    .A2(net48),
    .ZN(_07705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16461_ (.A1(_07704_),
    .A2(_07705_),
    .ZN(_07706_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17721 (.I(_03303_),
    .Z(net17721));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17726 (.I(_03282_),
    .Z(net17726));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16464_ (.A1(\u0.w[0][28] ),
    .A2(\u0.w[2][28] ),
    .Z(_07708_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16465_ (.A1(\u0.r0.out[28] ),
    .A2(_07708_),
    .Z(_07709_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16466_ (.A1(\u0.tmp_w[28] ),
    .A2(\u0.w[1][28] ),
    .Z(_07710_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16467_ (.A1(\u0.subword[28] ),
    .A2(_07710_),
    .Z(_07711_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16468_ (.A1(_07709_),
    .A2(_07711_),
    .Z(_07712_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16469_ (.A1(_07709_),
    .A2(_07711_),
    .ZN(_07713_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16470_ (.A1(_07712_),
    .A2(_07713_),
    .B(net21520),
    .ZN(_07714_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16471_ (.A1(net21519),
    .A2(net49),
    .Z(_07715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16472_ (.A1(_07714_),
    .A2(_07715_),
    .ZN(_07716_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _16473_ (.I(net20669),
    .ZN(_07717_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17761 (.I(_02410_),
    .Z(net17761));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16475_ (.A1(\u0.w[0][29] ),
    .A2(\u0.w[2][29] ),
    .Z(_07718_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16476_ (.A1(\u0.r0.out[29] ),
    .A2(_07718_),
    .Z(_07719_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16477_ (.A1(\u0.tmp_w[29] ),
    .A2(\u0.w[1][29] ),
    .Z(_07720_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16478_ (.A1(\u0.subword[29] ),
    .A2(_07720_),
    .Z(_07721_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16479_ (.A1(_07719_),
    .A2(_07721_),
    .Z(_07722_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16480_ (.A1(_07719_),
    .A2(_07721_),
    .ZN(_07723_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16481_ (.A1(_07722_),
    .A2(_07723_),
    .B(net21528),
    .ZN(_07724_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16482_ (.A1(net21528),
    .A2(net50),
    .Z(_07725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16483_ (.A1(_07724_),
    .A2(_07725_),
    .ZN(_07726_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _16484_ (.I(_07726_),
    .ZN(_07727_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17723 (.I(_03287_),
    .Z(net17723));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16486_ (.A1(\u0.w[0][30] ),
    .A2(\u0.w[2][30] ),
    .A3(\u0.r0.out[30] ),
    .Z(_07728_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16487_ (.I(\u0.w[1][30] ),
    .ZN(_07729_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16488_ (.A1(\u0.tmp_w[30] ),
    .A2(\u0.subword[30] ),
    .A3(_07729_),
    .Z(_07730_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16489_ (.A1(_07728_),
    .A2(_07730_),
    .Z(_07731_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16490_ (.I(net52),
    .ZN(_07732_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17717 (.I(_03319_),
    .Z(net17717));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16492_ (.A1(_07732_),
    .A2(net21538),
    .Z(_07734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16493_ (.A1(_07731_),
    .A2(net21525),
    .B(_07734_),
    .ZN(_07735_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17729 (.I(_03266_),
    .Z(net17729));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16495_ (.A1(\u0.w[0][31] ),
    .A2(\u0.w[2][31] ),
    .Z(_07736_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16496_ (.A1(\u0.r0.out[31] ),
    .A2(_07736_),
    .Z(_07737_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16497_ (.A1(\u0.w[1][31] ),
    .A2(\u0.subword[31] ),
    .A3(_07737_),
    .Z(_07738_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16498_ (.I(\u0.tmp_w[31] ),
    .ZN(_07739_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16499_ (.A1(_07738_),
    .A2(_07739_),
    .Z(_07740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16500_ (.A1(_07738_),
    .A2(_07739_),
    .ZN(_07741_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16501_ (.A1(_07740_),
    .A2(net21528),
    .A3(_07741_),
    .Z(_07742_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16502_ (.A1(net21528),
    .A2(net53),
    .ZN(_07743_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16503_ (.A1(_07742_),
    .A2(_07743_),
    .Z(_07744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16504_ (.I(_07744_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16505_ (.A1(net21127),
    .A2(net21128),
    .ZN(_07745_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17730 (.I(_03251_),
    .Z(net17730));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17759 (.I(_02425_),
    .Z(net17759));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16508_ (.I0(_07745_),
    .I1(net54),
    .S(net21535),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16509_ (.A1(net21126),
    .A2(_07547_),
    .ZN(_07748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16510_ (.I0(_07748_),
    .I1(net55),
    .S(net21535),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16511_ (.A1(_07557_),
    .A2(net21125),
    .ZN(_07749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16512_ (.I0(_07749_),
    .I1(net56),
    .S(net21535),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16513_ (.A1(net21122),
    .A2(_07564_),
    .ZN(_07750_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place17760 (.I(_02425_),
    .Z(net17760));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16515_ (.I0(_07750_),
    .I1(net57),
    .S(net21535),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16516_ (.A1(_07574_),
    .A2(_07573_),
    .ZN(_07752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16517_ (.I0(_07752_),
    .I1(net58),
    .S(net21535),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16518_ (.A1(_07581_),
    .A2(_07580_),
    .ZN(_07753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16519_ (.I0(_07753_),
    .I1(net59),
    .S(net21539),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16520_ (.A1(_07587_),
    .A2(_07588_),
    .ZN(_07754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16521_ (.I0(_07754_),
    .I1(net60),
    .S(net21539),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16522_ (.A1(_07592_),
    .A2(_07593_),
    .ZN(_07755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16523_ (.I0(_07755_),
    .I1(net61),
    .S(net21539),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16524_ (.A1(net21121),
    .A2(_07598_),
    .ZN(_07756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16525_ (.I0(_07756_),
    .I1(net63),
    .S(net21538),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16526_ (.A1(net21119),
    .A2(_07606_),
    .ZN(_07757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16527_ (.I0(_07757_),
    .I1(net64),
    .S(net21534),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16528_ (.A1(net21117),
    .A2(_07614_),
    .ZN(_07758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16529_ (.I0(_07758_),
    .I1(net65),
    .S(net21538),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16530_ (.A1(net21115),
    .A2(_07623_),
    .ZN(_07759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16531_ (.I0(_07759_),
    .I1(net66),
    .S(net21534),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16532_ (.A1(_07633_),
    .A2(_07632_),
    .ZN(_07760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16533_ (.I0(_07760_),
    .I1(net67),
    .S(net21534),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16534_ (.A1(_07642_),
    .A2(_07641_),
    .ZN(_07761_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17749 (.I(_02527_),
    .Z(net17749));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16536_ (.I0(_07761_),
    .I1(net68),
    .S(net21534),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16537_ (.A1(_07649_),
    .A2(_07648_),
    .ZN(_07763_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16538_ (.I0(_07763_),
    .I1(net69),
    .S(net21535),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16539_ (.A1(_07655_),
    .A2(_07656_),
    .ZN(_07764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16540_ (.I0(_07764_),
    .I1(net70),
    .S(net21535),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16541_ (.A1(net21134),
    .A2(_07361_),
    .ZN(_07765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16542_ (.I0(_07765_),
    .I1(net71),
    .S(net21535),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16543_ (.A1(net21131),
    .A2(net21132),
    .ZN(_07766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16544_ (.I0(_07766_),
    .I1(net72),
    .S(net21535),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16545_ (.A1(_07526_),
    .A2(net21129),
    .Z(_07767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16546_ (.I0(_07767_),
    .I1(net74),
    .S(net21535),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16547_ (.A1(net21135),
    .A2(_07232_),
    .ZN(_07768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16548_ (.I0(_07768_),
    .I1(net75),
    .S(net21535),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16549_ (.A1(net21130),
    .A2(_07489_),
    .ZN(_07769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16550_ (.I0(_07769_),
    .I1(net76),
    .S(net21538),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16551_ (.A1(_07475_),
    .A2(_07473_),
    .ZN(_07770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16552_ (.I0(_07770_),
    .I1(net77),
    .S(net21539),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16553_ (.A1(_07661_),
    .A2(_07662_),
    .ZN(_07771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16554_ (.I0(_07771_),
    .I1(net78),
    .S(net21538),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16555_ (.A1(_07667_),
    .A2(_07668_),
    .ZN(_07772_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17716 (.I(_03352_),
    .Z(net17716));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17718 (.I(_03309_),
    .Z(net17718));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16558_ (.I0(_07772_),
    .I1(net79),
    .S(net21535),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16559_ (.A1(net21113),
    .A2(_07674_),
    .ZN(_07775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16560_ (.I0(_07775_),
    .I1(net80),
    .S(net21535),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16561_ (.A1(net21194),
    .A2(net21253),
    .A3(net20962),
    .Z(_07776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16562_ (.I0(_07776_),
    .I1(net81),
    .S(net21535),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16563_ (.A1(net21111),
    .A2(net20961),
    .ZN(_07777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16564_ (.I0(_07777_),
    .I1(net82),
    .S(net21535),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16565_ (.A1(net21192),
    .A2(net21251),
    .A3(net20960),
    .Z(_07778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16566_ (.I0(_07778_),
    .I1(net83),
    .S(net21535),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16567_ (.A1(net21191),
    .A2(\u0.subword[28] ),
    .A3(_07709_),
    .Z(_07779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16568_ (.I0(_07779_),
    .I1(net85),
    .S(net21535),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16569_ (.A1(net21190),
    .A2(\u0.subword[29] ),
    .A3(_07719_),
    .Z(_07780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16570_ (.I0(_07780_),
    .I1(net86),
    .S(net21539),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16571_ (.A1(\u0.w[1][30] ),
    .A2(\u0.subword[30] ),
    .A3(_07728_),
    .Z(_07781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16572_ (.I0(_07781_),
    .I1(net87),
    .S(net21535),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16573_ (.I0(_07738_),
    .I1(net88),
    .S(net21535),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16574_ (.I(net21208),
    .ZN(_07782_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17741 (.I(_02680_),
    .Z(net17741));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16576_ (.I0(net21208),
    .I1(net89),
    .S(net21535),
    .Z(_07784_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16577_ (.A1(net21236),
    .A2(net21240),
    .Z(_07785_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17714 (.I(net17713),
    .Z(net17714));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16579_ (.A1(net21236),
    .A2(net21240),
    .ZN(_07787_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16580_ (.A1(_07785_),
    .A2(net21535),
    .A3(_07787_),
    .Z(_07788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16581_ (.I0(net21109),
    .I1(_07784_),
    .S(_07788_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17740 (.I(_02688_),
    .Z(net17740));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16583_ (.I0(net21199),
    .I1(net90),
    .S(net21535),
    .Z(_07790_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16584_ (.I(net21199),
    .ZN(_07791_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16585_ (.A1(net21226),
    .A2(net21239),
    .Z(_07792_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17724 (.I(_03287_),
    .Z(net17724));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16587_ (.A1(net21226),
    .A2(net21239),
    .ZN(_07794_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16588_ (.A1(_07792_),
    .A2(net21522),
    .A3(_07794_),
    .Z(_07795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16589_ (.I0(_07790_),
    .I1(_07791_),
    .S(_07795_),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16590_ (.I(net21189),
    .ZN(_07796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16591_ (.I0(net21189),
    .I1(net91),
    .S(net21535),
    .Z(_07797_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16592_ (.A1(net21238),
    .A2(net21217),
    .Z(_07798_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16593_ (.A1(net21238),
    .A2(net21217),
    .ZN(_07799_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16594_ (.A1(_07798_),
    .A2(net21535),
    .A3(_07799_),
    .Z(_07800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16595_ (.I0(_07796_),
    .I1(_07797_),
    .S(_07800_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16596_ (.I(net21188),
    .ZN(_07801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16597_ (.I0(net21188),
    .I1(net92),
    .S(net21535),
    .Z(_07802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16598_ (.A1(net21214),
    .A2(net21237),
    .Z(_07803_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16599_ (.A1(net21214),
    .A2(net21237),
    .ZN(_07804_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16600_ (.A1(_07803_),
    .A2(net21535),
    .A3(_07804_),
    .Z(_07805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16601_ (.I0(_07801_),
    .I1(_07802_),
    .S(_07805_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17725 (.I(_03282_),
    .Z(net17725));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16603_ (.I0(net21187),
    .I1(net93),
    .S(net21535),
    .Z(_07807_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16604_ (.I(net21187),
    .ZN(_07808_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16605_ (.A1(net21213),
    .A2(\u0.subword[4] ),
    .Z(_07809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16606_ (.A1(net21213),
    .A2(\u0.subword[4] ),
    .ZN(_07810_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16607_ (.A1(_07809_),
    .A2(net21522),
    .A3(_07810_),
    .Z(_07811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16608_ (.I0(_07807_),
    .I1(_07808_),
    .S(_07811_),
    .Z(_00347_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16609_ (.A1(net21212),
    .A2(\u0.subword[5] ),
    .Z(_07812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16610_ (.A1(net21212),
    .A2(\u0.subword[5] ),
    .ZN(_07813_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16611_ (.A1(_07812_),
    .A2(net21525),
    .A3(_07813_),
    .Z(_07814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16612_ (.I0(net21186),
    .I1(net94),
    .S(net21535),
    .Z(_07815_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16613_ (.A1(_07814_),
    .A2(_07815_),
    .ZN(_07816_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16614_ (.A1(net21186),
    .A2(_07814_),
    .B(_07816_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16615_ (.A1(\u0.w[0][6] ),
    .A2(\u0.subword[6] ),
    .Z(_07817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16616_ (.A1(\u0.w[0][6] ),
    .A2(\u0.subword[6] ),
    .ZN(_07818_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16617_ (.A1(_07817_),
    .A2(net21525),
    .A3(_07818_),
    .Z(_07819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16618_ (.I0(net21185),
    .I1(net96),
    .S(net21539),
    .Z(_07820_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16619_ (.A1(_07819_),
    .A2(_07820_),
    .ZN(_07821_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16620_ (.A1(net21185),
    .A2(_07819_),
    .B(_07821_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16621_ (.A1(\u0.w[0][7] ),
    .A2(\u0.subword[7] ),
    .Z(_07822_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16622_ (.A1(\u0.w[0][7] ),
    .A2(\u0.subword[7] ),
    .ZN(_07823_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16623_ (.A1(_07822_),
    .A2(net21539),
    .A3(_07823_),
    .Z(_07824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16624_ (.I0(net21184),
    .I1(net97),
    .S(net21539),
    .Z(_07825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16625_ (.A1(_07824_),
    .A2(_07825_),
    .ZN(_07826_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16626_ (.A1(net21184),
    .A2(_07824_),
    .B(_07826_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16627_ (.I0(net21183),
    .I1(net98),
    .S(net21534),
    .Z(_07827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16628_ (.I(net21183),
    .ZN(_07828_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16629_ (.A1(net21211),
    .A2(net21245),
    .Z(_07829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16630_ (.A1(net21211),
    .A2(net21245),
    .ZN(_07830_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16631_ (.A1(_07829_),
    .A2(net21523),
    .A3(_07830_),
    .Z(_07831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16632_ (.I0(_07827_),
    .I1(net21108),
    .S(_07831_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16633_ (.I0(net21182),
    .I1(net99),
    .S(net21534),
    .Z(_07832_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16634_ (.I(net21182),
    .ZN(_07833_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16635_ (.A1(net21209),
    .A2(net21244),
    .Z(_07834_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17706 (.I(_03887_),
    .Z(net17706));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16637_ (.A1(net21209),
    .A2(net21244),
    .ZN(_07836_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16638_ (.A1(_07834_),
    .A2(net21521),
    .A3(_07836_),
    .Z(_07837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16639_ (.I0(_07832_),
    .I1(_07833_),
    .S(_07837_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16640_ (.I0(net21207),
    .I1(net100),
    .S(net21535),
    .Z(_07838_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16641_ (.I(net21207),
    .ZN(_07839_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16642_ (.A1(net21243),
    .A2(net21235),
    .Z(_07840_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16643_ (.A1(net21243),
    .A2(net21235),
    .ZN(_07841_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16644_ (.A1(_07840_),
    .A2(net21521),
    .A3(_07841_),
    .Z(_07842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16645_ (.I0(_07838_),
    .I1(_07839_),
    .S(_07842_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16646_ (.I(net21206),
    .ZN(_07843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16647_ (.I0(net21206),
    .I1(net101),
    .S(net21534),
    .Z(_07844_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16648_ (.A1(net21234),
    .A2(net21242),
    .Z(_07845_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16649_ (.A1(net21234),
    .A2(net21242),
    .ZN(_07846_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16650_ (.A1(_07845_),
    .A2(net21534),
    .A3(_07846_),
    .Z(_07847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16651_ (.I0(_07843_),
    .I1(_07844_),
    .S(_07847_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16652_ (.I0(net21205),
    .I1(net102),
    .S(net21534),
    .Z(_07848_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16653_ (.I(net21205),
    .ZN(_07849_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16654_ (.A1(net21233),
    .A2(net21241),
    .Z(_07850_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16655_ (.A1(net21233),
    .A2(net21241),
    .ZN(_07851_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16656_ (.A1(_07850_),
    .A2(net21523),
    .A3(_07851_),
    .Z(_07852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16657_ (.I0(_07848_),
    .I1(_07849_),
    .S(_07852_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16658_ (.A1(net21232),
    .A2(\u0.subword[13] ),
    .Z(_07853_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16659_ (.A1(net21232),
    .A2(\u0.subword[13] ),
    .ZN(_07854_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16660_ (.A1(_07853_),
    .A2(net21534),
    .A3(_07854_),
    .Z(_07855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16661_ (.I0(net21204),
    .I1(net103),
    .S(net21534),
    .Z(_07856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16662_ (.A1(_07855_),
    .A2(_07856_),
    .ZN(_07857_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16663_ (.A1(net21204),
    .A2(_07855_),
    .B(_07857_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16664_ (.A1(net21231),
    .A2(\u0.subword[14] ),
    .Z(_07858_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16665_ (.A1(net21231),
    .A2(\u0.subword[14] ),
    .ZN(_07859_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16666_ (.A1(_07858_),
    .A2(net21535),
    .A3(_07859_),
    .Z(_07860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16667_ (.I0(\u0.w[1][14] ),
    .I1(net104),
    .S(net21535),
    .Z(_07861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16668_ (.A1(_07860_),
    .A2(_07861_),
    .ZN(_07862_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16669_ (.A1(\u0.w[1][14] ),
    .A2(_07860_),
    .B(_07862_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16670_ (.A1(\u0.w[0][15] ),
    .A2(\u0.subword[15] ),
    .Z(_07863_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16671_ (.A1(\u0.w[0][15] ),
    .A2(\u0.subword[15] ),
    .ZN(_07864_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16672_ (.A1(_07863_),
    .A2(net21535),
    .A3(_07864_),
    .Z(_07865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16673_ (.I0(\u0.w[1][15] ),
    .I1(net105),
    .S(net21535),
    .Z(_07866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16674_ (.A1(_07865_),
    .A2(_07866_),
    .ZN(_07867_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16675_ (.A1(\u0.w[1][15] ),
    .A2(_07865_),
    .B(_07867_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16676_ (.I0(net21203),
    .I1(net107),
    .S(net21535),
    .Z(_07868_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16677_ (.I(net21203),
    .ZN(_07869_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16678_ (.A1(net21230),
    .A2(net21250),
    .Z(_07870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16679_ (.A1(net21230),
    .A2(net21250),
    .ZN(_07871_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16680_ (.A1(_07870_),
    .A2(net21521),
    .A3(_07871_),
    .Z(_07872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16681_ (.I0(_07868_),
    .I1(net21107),
    .S(_07872_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16682_ (.I0(net21202),
    .I1(net108),
    .S(net21534),
    .Z(_07873_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16683_ (.I(net21202),
    .ZN(_07874_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16684_ (.A1(net21229),
    .A2(net21249),
    .Z(_07875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16685_ (.A1(net21229),
    .A2(net21249),
    .ZN(_07876_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16686_ (.A1(_07875_),
    .A2(net21521),
    .A3(_07876_),
    .Z(_07877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16687_ (.I0(_07873_),
    .I1(net21106),
    .S(_07877_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16688_ (.I0(net21201),
    .I1(net109),
    .S(net21535),
    .Z(_07878_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16689_ (.I(net21201),
    .ZN(_07879_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16690_ (.A1(\u0.subword[18] ),
    .A2(net21228),
    .Z(_07880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16691_ (.A1(\u0.subword[18] ),
    .A2(net21228),
    .ZN(_07881_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16692_ (.A1(_07880_),
    .A2(net21521),
    .A3(_07881_),
    .Z(_07882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16693_ (.I0(_07878_),
    .I1(_07879_),
    .S(_07882_),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16694_ (.I0(net21200),
    .I1(net110),
    .S(net21535),
    .Z(_07883_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16695_ (.I(net21200),
    .ZN(_07884_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16696_ (.A1(net21227),
    .A2(net21248),
    .Z(_07885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16697_ (.A1(net21227),
    .A2(net21248),
    .ZN(_07886_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16698_ (.A1(_07885_),
    .A2(net21521),
    .A3(_07886_),
    .Z(_07887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16699_ (.I0(_07883_),
    .I1(_07884_),
    .S(_07887_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16700_ (.I(net21198),
    .ZN(_07888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16701_ (.I0(net21198),
    .I1(net111),
    .S(net21535),
    .Z(_07889_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16702_ (.A1(net21225),
    .A2(net21247),
    .Z(_07890_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16703_ (.A1(net21225),
    .A2(net21247),
    .ZN(_07891_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16704_ (.A1(_07890_),
    .A2(net21538),
    .A3(_07891_),
    .Z(_07892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16705_ (.I0(_07888_),
    .I1(_07889_),
    .S(_07892_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16706_ (.I(net21197),
    .ZN(_07893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16707_ (.I0(net21197),
    .I1(net112),
    .S(net21535),
    .Z(_07894_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16708_ (.A1(net21224),
    .A2(net21246),
    .Z(_07895_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16709_ (.A1(net21224),
    .A2(net21246),
    .ZN(_07896_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16710_ (.A1(_07895_),
    .A2(net21538),
    .A3(_07896_),
    .Z(_07897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16711_ (.I0(_07893_),
    .I1(_07894_),
    .S(_07897_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16712_ (.I0(net21196),
    .I1(net113),
    .S(net21538),
    .Z(_07898_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16713_ (.I(net21196),
    .ZN(_07899_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16714_ (.A1(\u0.w[0][22] ),
    .A2(\u0.subword[22] ),
    .Z(_07900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16715_ (.A1(\u0.w[0][22] ),
    .A2(\u0.subword[22] ),
    .ZN(_07901_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16716_ (.A1(_07900_),
    .A2(net21521),
    .A3(_07901_),
    .Z(_07902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16717_ (.I0(_07898_),
    .I1(_07899_),
    .S(_07902_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16718_ (.I0(\u0.w[1][23] ),
    .I1(net114),
    .S(net21535),
    .Z(_07903_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16719_ (.I(\u0.w[1][23] ),
    .ZN(_07904_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16720_ (.A1(\u0.w[0][23] ),
    .A2(\u0.subword[23] ),
    .Z(_07905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16721_ (.A1(\u0.w[0][23] ),
    .A2(\u0.subword[23] ),
    .ZN(_07906_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16722_ (.A1(_07905_),
    .A2(net21521),
    .A3(_07906_),
    .Z(_07907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16723_ (.I0(_07903_),
    .I1(_07904_),
    .S(_07907_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16724_ (.I(net21195),
    .ZN(_07908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16725_ (.I0(net21195),
    .I1(net115),
    .S(net21535),
    .Z(_07909_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16726_ (.A1(net21223),
    .A2(net21254),
    .A3(net21257),
    .Z(_07910_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17713 (.I(_03367_),
    .Z(net17713));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16728_ (.A1(_07910_),
    .A2(net21522),
    .ZN(_07912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16729_ (.I0(net21105),
    .I1(_07909_),
    .S(_07912_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16730_ (.I(net21194),
    .ZN(_07913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16731_ (.I0(net21194),
    .I1(net116),
    .S(net21535),
    .Z(_07914_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16732_ (.A1(net21222),
    .A2(net21253),
    .A3(net21256),
    .Z(_07915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16733_ (.A1(_07915_),
    .A2(net21522),
    .ZN(_07916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16734_ (.I0(net21104),
    .I1(_07914_),
    .S(_07916_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16735_ (.I(net21193),
    .ZN(_07917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16736_ (.I0(net21193),
    .I1(net118),
    .S(net21535),
    .Z(_07918_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16737_ (.A1(net21221),
    .A2(net21252),
    .A3(net21255),
    .Z(_07919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16738_ (.A1(_07919_),
    .A2(net21522),
    .ZN(_07920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16739_ (.I0(_07917_),
    .I1(_07918_),
    .S(_07920_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16740_ (.I(net21192),
    .ZN(_07921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16741_ (.I0(net21192),
    .I1(net119),
    .S(net21535),
    .Z(_07922_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16742_ (.A1(net21220),
    .A2(net21251),
    .A3(\u0.r0.out[27] ),
    .Z(_07923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16743_ (.A1(_07923_),
    .A2(net21522),
    .ZN(_07924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16744_ (.I0(_07921_),
    .I1(_07922_),
    .S(_07924_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16745_ (.I(net21191),
    .ZN(_07925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16746_ (.I0(net21191),
    .I1(net120),
    .S(net21535),
    .Z(_07926_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16747_ (.A1(net21219),
    .A2(\u0.subword[28] ),
    .A3(\u0.r0.out[28] ),
    .Z(_07927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16748_ (.A1(_07927_),
    .A2(net21521),
    .ZN(_07928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16749_ (.I0(_07925_),
    .I1(_07926_),
    .S(_07928_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16750_ (.I(net21190),
    .ZN(_07929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16751_ (.I0(net21190),
    .I1(net121),
    .S(net21539),
    .Z(_07930_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16752_ (.A1(net21218),
    .A2(\u0.subword[29] ),
    .A3(\u0.r0.out[29] ),
    .Z(_07931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16753_ (.A1(_07931_),
    .A2(net21525),
    .ZN(_07932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16754_ (.I0(_07929_),
    .I1(_07930_),
    .S(_07932_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16755_ (.I0(\u0.w[1][30] ),
    .I1(net122),
    .S(net21535),
    .Z(_07933_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16756_ (.A1(net21216),
    .A2(\u0.subword[30] ),
    .A3(\u0.r0.out[30] ),
    .Z(_07934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16757_ (.A1(_07934_),
    .A2(net21522),
    .ZN(_07935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16758_ (.I0(_07729_),
    .I1(_07933_),
    .S(_07935_),
    .Z(_00344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16759_ (.I(\u0.w[1][31] ),
    .ZN(_07936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16760_ (.I0(\u0.w[1][31] ),
    .I1(net123),
    .S(net21535),
    .Z(_07937_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _16761_ (.A1(net21215),
    .A2(\u0.subword[31] ),
    .A3(\u0.r0.out[31] ),
    .Z(_07938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16762_ (.A1(_07938_),
    .A2(net21522),
    .ZN(_07939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16763_ (.I0(_07936_),
    .I1(_07937_),
    .S(_07939_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17719 (.I(net17718),
    .Z(net17719));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16765_ (.A1(net21535),
    .A2(net124),
    .ZN(_07941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16766_ (.A1(_07788_),
    .A2(_07941_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17703 (.I(_03933_),
    .Z(net17703));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16768_ (.A1(net21535),
    .A2(net125),
    .Z(_07943_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16769_ (.A1(_07795_),
    .A2(_07943_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16770_ (.A1(net21535),
    .A2(net126),
    .ZN(_07944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16771_ (.A1(_07800_),
    .A2(_07944_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16772_ (.A1(net21535),
    .A2(net127),
    .ZN(_07945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16773_ (.A1(_07805_),
    .A2(_07945_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16774_ (.A1(net21535),
    .A2(net2),
    .Z(_07946_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16775_ (.A1(_07811_),
    .A2(_07946_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16776_ (.A1(net21535),
    .A2(net3),
    .Z(_07947_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16777_ (.A1(_07814_),
    .A2(_07947_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17702 (.I(net17701),
    .Z(net17702));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16779_ (.A1(net21539),
    .A2(net4),
    .Z(_07949_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16780_ (.A1(_07819_),
    .A2(_07949_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16781_ (.A1(net21539),
    .A2(net5),
    .ZN(_07950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16782_ (.A1(_07824_),
    .A2(_07950_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16783_ (.A1(net21534),
    .A2(net6),
    .Z(_07951_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16784_ (.A1(_07831_),
    .A2(_07951_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16785_ (.A1(net21534),
    .A2(net7),
    .Z(_07952_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16786_ (.A1(_07837_),
    .A2(_07952_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16787_ (.A1(net21535),
    .A2(net8),
    .Z(_07953_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16788_ (.A1(_07842_),
    .A2(_07953_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17704 (.I(_03903_),
    .Z(net17704));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16790_ (.A1(net21534),
    .A2(net9),
    .ZN(_07955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16791_ (.A1(_07847_),
    .A2(_07955_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16792_ (.A1(net21534),
    .A2(net10),
    .Z(_07956_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16793_ (.A1(_07852_),
    .A2(_07956_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16794_ (.A1(net21534),
    .A2(net11),
    .ZN(_07957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16795_ (.A1(_07855_),
    .A2(_07957_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16796_ (.A1(net21535),
    .A2(net13),
    .ZN(_07958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16797_ (.A1(_07860_),
    .A2(_07958_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16798_ (.A1(net21535),
    .A2(net14),
    .ZN(_07959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16799_ (.A1(_07865_),
    .A2(_07959_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16800_ (.A1(net21535),
    .A2(net15),
    .Z(_07960_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16801_ (.A1(_07872_),
    .A2(_07960_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16802_ (.A1(net21534),
    .A2(net16),
    .Z(_07961_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16803_ (.A1(_07877_),
    .A2(_07961_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16804_ (.A1(net21535),
    .A2(net17),
    .Z(_07962_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16805_ (.A1(_07882_),
    .A2(_07962_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16806_ (.A1(net21535),
    .A2(net18),
    .Z(_07963_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16807_ (.A1(_07887_),
    .A2(_07963_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16808_ (.A1(net21538),
    .A2(net19),
    .ZN(_07964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16809_ (.A1(_07892_),
    .A2(_07964_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16810_ (.A1(net21538),
    .A2(net20),
    .ZN(_07965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16811_ (.A1(_07897_),
    .A2(_07965_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16812_ (.A1(net21538),
    .A2(net21),
    .Z(_07966_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16813_ (.A1(_07902_),
    .A2(_07966_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16814_ (.A1(net21535),
    .A2(net22),
    .Z(_07967_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16815_ (.A1(_07907_),
    .A2(_07967_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16816_ (.A1(net21535),
    .A2(net24),
    .ZN(_07968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16817_ (.A1(_07912_),
    .A2(_07968_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16818_ (.A1(net21535),
    .A2(net25),
    .ZN(_07969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16819_ (.A1(_07916_),
    .A2(_07969_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16820_ (.A1(net21535),
    .A2(net26),
    .ZN(_07970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16821_ (.A1(_07920_),
    .A2(_07970_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16822_ (.A1(net21535),
    .A2(net27),
    .ZN(_07971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16823_ (.A1(_07924_),
    .A2(_07971_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16824_ (.A1(net21535),
    .A2(net28),
    .ZN(_07972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16825_ (.A1(_07928_),
    .A2(_07972_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16826_ (.A1(net21539),
    .A2(net29),
    .ZN(_07973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16827_ (.A1(_07932_),
    .A2(_07973_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16828_ (.A1(net21535),
    .A2(net30),
    .ZN(_07974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16829_ (.A1(_07935_),
    .A2(_07974_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16830_ (.A1(net21535),
    .A2(net31),
    .ZN(_07975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16831_ (.A1(_07939_),
    .A2(_07975_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16832_ (.A1(net21530),
    .A2(_07466_),
    .B(_07471_),
    .ZN(_15537_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16833_ (.I(_07536_),
    .ZN(_07976_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17695 (.I(_04022_),
    .Z(net17695));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16835_ (.A1(net21530),
    .A2(_07394_),
    .B(_07448_),
    .ZN(_15538_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16836_ (.I(_15553_[0]),
    .ZN(_07977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16837_ (.A1(net20556),
    .A2(_07977_),
    .ZN(_07978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16838_ (.I(_07978_),
    .ZN(_07979_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16839_ (.I(_15549_[0]),
    .ZN(_07980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16840_ (.A1(net20778),
    .A2(_07980_),
    .ZN(_07981_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16841_ (.I(_07981_),
    .ZN(_07982_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16842_ (.A1(_07979_),
    .A2(_07982_),
    .B(net20610),
    .ZN(_07983_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16843_ (.I(_07513_),
    .ZN(_07984_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17709 (.I(_03881_),
    .Z(net17709));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17710 (.I(_03837_),
    .Z(net17710));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16846_ (.I(_15540_[0]),
    .ZN(_07987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16847_ (.A1(_07536_),
    .A2(_07987_),
    .ZN(_07988_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17707 (.I(_03881_),
    .Z(net17707));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16849_ (.A1(net20794),
    .A2(_07988_),
    .Z(_07990_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17693 (.I(_04091_),
    .Z(net17693));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17697 (.I(_03988_),
    .Z(net17697));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16852_ (.A1(net20863),
    .A2(_15539_[0]),
    .A3(net21517),
    .ZN(_07993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16853_ (.A1(_07990_),
    .A2(net20541),
    .ZN(_07994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16854_ (.A1(_07994_),
    .A2(net20551),
    .A3(_07983_),
    .ZN(_07995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16855_ (.A1(net20779),
    .A2(net20833),
    .ZN(_07996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16856_ (.A1(_07996_),
    .A2(net20794),
    .Z(_07997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16857_ (.A1(net20793),
    .A2(net20792),
    .ZN(_07998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16858_ (.A1(_07997_),
    .A2(_07998_),
    .ZN(_07999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16859_ (.A1(_07998_),
    .A2(_07996_),
    .ZN(_08000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17746 (.I(_02585_),
    .Z(net17746));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16861_ (.A1(_08000_),
    .A2(net20608),
    .ZN(_08002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16862_ (.A1(_07999_),
    .A2(_08002_),
    .A3(net20782),
    .ZN(_08003_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16863_ (.A1(_07995_),
    .A2(_08003_),
    .A3(net20789),
    .ZN(_08004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16864_ (.A1(net20554),
    .A2(net20836),
    .ZN(_08005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16865_ (.A1(net20777),
    .A2(net20624),
    .ZN(_08006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16866_ (.A1(_08005_),
    .A2(_08006_),
    .ZN(_08007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17700 (.I(_03971_),
    .Z(net17700));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17701 (.I(_03963_),
    .Z(net17701));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16869_ (.A1(_08007_),
    .A2(net20794),
    .ZN(_08010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16870_ (.A1(net20863),
    .A2(net21515),
    .A3(_07987_),
    .ZN(_08011_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16871_ (.I(_08011_),
    .ZN(_08012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16872_ (.A1(net20614),
    .A2(_08012_),
    .ZN(_08013_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16873_ (.A1(_08010_),
    .A2(net20782),
    .A3(_08013_),
    .ZN(_08014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16874_ (.A1(net20777),
    .A2(_07977_),
    .ZN(_08015_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16875_ (.I(_08015_),
    .ZN(_08016_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17690 (.I(_04608_),
    .Z(net17690));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17689 (.I(_04661_),
    .Z(net17689));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16878_ (.A1(_08016_),
    .A2(net20794),
    .B(net20782),
    .ZN(_08019_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16879_ (.A1(net20864),
    .A2(net20386),
    .A3(net21517),
    .ZN(_08020_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17818 (.I(_00940_),
    .Z(net17818));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16881_ (.A1(net20366),
    .A2(_08020_),
    .A3(_07330_),
    .ZN(_08022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16882_ (.A1(net20555),
    .A2(_07980_),
    .ZN(_08023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16883_ (.I(_08023_),
    .ZN(_08024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16884_ (.A1(_08024_),
    .A2(net20802),
    .ZN(_08025_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16885_ (.A1(_08019_),
    .A2(_08022_),
    .A3(_08025_),
    .ZN(_08026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16886_ (.I(_07484_),
    .ZN(_08027_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17686 (.I(_04768_),
    .Z(net17686));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16888_ (.A1(_08014_),
    .A2(_08026_),
    .A3(net20536),
    .ZN(_08029_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _16889_ (.I(_07666_),
    .ZN(_08030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17711 (.I(_03373_),
    .Z(net17711));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16891_ (.A1(_08030_),
    .A2(_08029_),
    .A3(_08004_),
    .ZN(_08032_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16892_ (.A1(net20777),
    .A2(net20836),
    .ZN(_08033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16893_ (.A1(_08033_),
    .A2(net20794),
    .ZN(_08034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17684 (.I(_04777_),
    .Z(net17684));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16895_ (.A1(_08034_),
    .A2(net20542),
    .Z(_08036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16896_ (.A1(_07976_),
    .A2(net20793),
    .ZN(_08037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16897_ (.A1(net20778),
    .A2(_15539_[0]),
    .ZN(_08038_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16898_ (.A1(_08037_),
    .A2(net20607),
    .A3(_08038_),
    .ZN(_08039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16899_ (.A1(net20777),
    .A2(_15555_[0]),
    .Z(_08040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16900_ (.A1(_08040_),
    .A2(net20794),
    .ZN(_08041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16901_ (.A1(_08036_),
    .A2(_08039_),
    .A3(_08041_),
    .ZN(_08042_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16902_ (.I(_15541_[0]),
    .ZN(_08043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16903_ (.A1(net20780),
    .A2(_08043_),
    .ZN(_08044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16904_ (.A1(_08044_),
    .A2(net20607),
    .Z(_08045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16905_ (.A1(_08045_),
    .A2(net20364),
    .ZN(_08046_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17683 (.I(_04782_),
    .Z(net17683));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16907_ (.A1(net20792),
    .A2(net20777),
    .ZN(_08048_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17682 (.I(_04971_),
    .Z(net17682));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16909_ (.A1(net20863),
    .A2(net20388),
    .A3(net21516),
    .ZN(_08050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16910_ (.A1(net20528),
    .A2(net20794),
    .A3(net20359),
    .ZN(_08051_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16911_ (.A1(_08046_),
    .A2(net20783),
    .A3(_08051_),
    .ZN(_08052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16912_ (.A1(_08042_),
    .A2(_08052_),
    .A3(net20536),
    .ZN(_08053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16913_ (.A1(_08050_),
    .A2(net20794),
    .ZN(_08054_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16914_ (.I(_08054_),
    .ZN(_08055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16915_ (.A1(net20793),
    .A2(net20777),
    .ZN(_08056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16916_ (.A1(_08055_),
    .A2(net20525),
    .ZN(_08057_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16917_ (.A1(net20863),
    .A2(_08043_),
    .A3(net21515),
    .ZN(_08058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16918_ (.A1(_08058_),
    .A2(net20603),
    .ZN(_08059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _16919_ (.I(_08059_),
    .ZN(_08060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16920_ (.A1(_08060_),
    .A2(net20366),
    .ZN(_08061_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16921_ (.A1(_08057_),
    .A2(_08061_),
    .A3(net20783),
    .ZN(_08062_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17681 (.I(_04993_),
    .Z(net17681));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16923_ (.A1(_08050_),
    .A2(net20611),
    .ZN(_08064_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _16924_ (.I(_08064_),
    .ZN(_08065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16925_ (.I(_15546_[0]),
    .ZN(_08066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16926_ (.A1(net20777),
    .A2(_08066_),
    .ZN(_08067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16927_ (.A1(_08065_),
    .A2(net20145),
    .ZN(_08068_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17685 (.I(_04775_),
    .Z(net17685));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16929_ (.A1(_08037_),
    .A2(net20794),
    .ZN(_08070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16930_ (.A1(_08068_),
    .A2(net20544),
    .A3(net20143),
    .ZN(_08071_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17679 (.I(_05012_),
    .Z(net17679));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16932_ (.A1(_08062_),
    .A2(_08071_),
    .A3(net20789),
    .ZN(_08073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16933_ (.A1(_08053_),
    .A2(_08073_),
    .A3(net20846),
    .ZN(_08074_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _16934_ (.I(_00394_),
    .ZN(_08075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17691 (.I(_04328_),
    .Z(net17691));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16936_ (.A1(_08032_),
    .A2(_08074_),
    .A3(_08075_),
    .ZN(_08077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16937_ (.A1(_07979_),
    .A2(net20363),
    .B(net20799),
    .ZN(_08078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16938_ (.A1(_08067_),
    .A2(_07330_),
    .Z(_08079_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17743 (.I(_02632_),
    .Z(net17743));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16940_ (.A1(_08079_),
    .A2(net20542),
    .ZN(_08081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17687 (.I(_04768_),
    .Z(net17687));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16942_ (.A1(_08078_),
    .A2(_08081_),
    .B(net20536),
    .ZN(_08083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16943_ (.A1(net20778),
    .A2(net20835),
    .ZN(_08084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16944_ (.A1(_08084_),
    .A2(net20794),
    .Z(_08085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16945_ (.A1(net20863),
    .A2(net20624),
    .A3(net21515),
    .ZN(_08086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16946_ (.A1(_08085_),
    .A2(net20522),
    .ZN(_08087_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16947_ (.A1(net20863),
    .A2(_15549_[0]),
    .A3(net21515),
    .ZN(_08088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16948_ (.A1(net20526),
    .A2(net20613),
    .A3(net20354),
    .ZN(_08089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16949_ (.A1(_08087_),
    .A2(net20542),
    .A3(_08089_),
    .ZN(_08090_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17675 (.I(_05371_),
    .Z(net17675));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16951_ (.A1(_08083_),
    .A2(_08090_),
    .B(_08030_),
    .ZN(_08092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16952_ (.A1(_07988_),
    .A2(_07330_),
    .ZN(_08093_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16953_ (.I(_08093_),
    .ZN(_08094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16954_ (.I(_15551_[0]),
    .ZN(_08095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16955_ (.A1(net20863),
    .A2(net21515),
    .B(_08095_),
    .ZN(_08096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16956_ (.A1(_08096_),
    .A2(net20794),
    .Z(_08097_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16957_ (.A1(_08094_),
    .A2(_08097_),
    .A3(net20553),
    .ZN(_08098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16958_ (.A1(_08039_),
    .A2(net20542),
    .Z(_08099_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16959_ (.A1(net20863),
    .A2(_15546_[0]),
    .A3(net21517),
    .ZN(_08100_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16960_ (.A1(_08100_),
    .A2(_07330_),
    .Z(_08101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16961_ (.A1(_08099_),
    .A2(_08098_),
    .B(net20139),
    .ZN(_08102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16962_ (.A1(_08102_),
    .A2(net20535),
    .ZN(_08103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16963_ (.A1(_08103_),
    .A2(_08092_),
    .ZN(_08104_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16964_ (.I(_15544_[0]),
    .ZN(_08105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16965_ (.A1(net20778),
    .A2(_08105_),
    .Z(_08106_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17674 (.I(_05371_),
    .Z(net17674));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16967_ (.A1(_08106_),
    .A2(net20798),
    .B(net20542),
    .ZN(_08108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16968_ (.A1(_08040_),
    .A2(_07330_),
    .ZN(_08109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16969_ (.A1(_08108_),
    .A2(_08025_),
    .A3(net20138),
    .ZN(_08110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16970_ (.A1(net20863),
    .A2(net21515),
    .A3(_08095_),
    .ZN(_08111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16971_ (.A1(_08111_),
    .A2(_07330_),
    .ZN(_08112_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16972_ (.I(_08112_),
    .ZN(_08113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16973_ (.A1(net20778),
    .A2(_15544_[0]),
    .ZN(_08114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16974_ (.A1(_08113_),
    .A2(_08114_),
    .ZN(_08115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17669 (.I(_05398_),
    .Z(net17669));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16976_ (.A1(_08115_),
    .A2(net20550),
    .A3(_08041_),
    .ZN(_08117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16977_ (.A1(_08110_),
    .A2(_08117_),
    .A3(net20789),
    .ZN(_08118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16978_ (.A1(net20777),
    .A2(net20386),
    .ZN(_08119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16979_ (.A1(_08037_),
    .A2(net20614),
    .A3(_08119_),
    .ZN(_08120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16980_ (.A1(_07976_),
    .A2(net20833),
    .ZN(_08121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16981_ (.A1(net20347),
    .A2(net20798),
    .A3(_08114_),
    .ZN(_08122_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16982_ (.A1(net20136),
    .A2(_08122_),
    .A3(net20553),
    .ZN(_08123_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17666 (.I(_05432_),
    .Z(net17666));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17673 (.I(net17672),
    .Z(net17673));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16985_ (.A1(net20614),
    .A2(_15565_[0]),
    .ZN(_08126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17665 (.I(_05443_),
    .Z(net17665));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16987_ (.A1(net20614),
    .A2(net20522),
    .B(_08126_),
    .C(net20782),
    .ZN(_08128_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16988_ (.A1(_08123_),
    .A2(net20535),
    .A3(_08128_),
    .ZN(_08129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16989_ (.A1(_08118_),
    .A2(_08129_),
    .A3(_08030_),
    .ZN(_08130_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16990_ (.A1(_08104_),
    .A2(_08130_),
    .A3(net20845),
    .ZN(_08131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16991_ (.A1(_08131_),
    .A2(_08077_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16992_ (.A1(_08056_),
    .A2(net20794),
    .Z(_08132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16993_ (.A1(_08132_),
    .A2(_08020_),
    .ZN(_08133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16994_ (.A1(_08065_),
    .A2(net20529),
    .ZN(_08134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16995_ (.A1(_08133_),
    .A2(net20789),
    .A3(_08134_),
    .ZN(_08135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16996_ (.A1(_08135_),
    .A2(net20787),
    .ZN(_08136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16997_ (.A1(_07997_),
    .A2(_08005_),
    .ZN(_08137_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16998_ (.I(_08033_),
    .ZN(_08138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16999_ (.A1(_08079_),
    .A2(_08138_),
    .ZN(_08139_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17000_ (.A1(_08137_),
    .A2(_08139_),
    .A3(net20532),
    .Z(_08140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17001_ (.A1(_08088_),
    .A2(net20794),
    .ZN(_08141_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17002_ (.I(_08141_),
    .ZN(_08142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17003_ (.A1(_08142_),
    .A2(_08038_),
    .ZN(_08143_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17004_ (.I(_08143_),
    .ZN(_08144_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17005_ (.I(_15567_[0]),
    .ZN(_08145_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17006_ (.A1(_08027_),
    .A2(_08145_),
    .A3(net20605),
    .Z(_08146_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17007_ (.A1(_08144_),
    .A2(_08146_),
    .B(net20548),
    .ZN(_08147_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17008_ (.A1(_08136_),
    .A2(_08140_),
    .B(_08030_),
    .C(_08147_),
    .ZN(_08148_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17009_ (.I(_08121_),
    .ZN(_08149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17010_ (.A1(_08149_),
    .A2(net20794),
    .ZN(_08150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17011_ (.A1(_08150_),
    .A2(_08041_),
    .Z(_08151_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17012_ (.I(_08086_),
    .ZN(_08152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17013_ (.A1(_08152_),
    .A2(net20605),
    .ZN(_08153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17014_ (.A1(_08153_),
    .A2(net20782),
    .Z(_08154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17015_ (.A1(_08016_),
    .A2(net20613),
    .ZN(_08155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17016_ (.A1(_08151_),
    .A2(_08154_),
    .A3(net19445),
    .ZN(_08156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17017_ (.A1(_07997_),
    .A2(_08020_),
    .ZN(_08157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17018_ (.A1(_08157_),
    .A2(_08139_),
    .A3(net20550),
    .ZN(_08158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17019_ (.A1(_08156_),
    .A2(net20789),
    .A3(_08158_),
    .ZN(_08159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17020_ (.A1(net20349),
    .A2(net20542),
    .ZN(_08160_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17021_ (.A1(_08094_),
    .A2(_08160_),
    .ZN(_08161_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17022_ (.I(_15539_[0]),
    .ZN(_08162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17023_ (.A1(net20778),
    .A2(_08162_),
    .ZN(_08163_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17024_ (.A1(_08163_),
    .A2(net20608),
    .Z(_08164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17025_ (.A1(_08161_),
    .A2(_08164_),
    .B(net20790),
    .ZN(_08165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17026_ (.A1(_08044_),
    .A2(net20794),
    .ZN(_08166_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17027_ (.I(_08166_),
    .ZN(_08167_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17028_ (.A1(net20778),
    .A2(_15555_[0]),
    .Z(_08168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17029_ (.A1(_08167_),
    .A2(net20344),
    .ZN(_08169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17030_ (.A1(_07993_),
    .A2(net20606),
    .ZN(_08170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17031_ (.I(_08170_),
    .ZN(_08171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17032_ (.A1(_08171_),
    .A2(net20538),
    .ZN(_08172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17033_ (.A1(_08169_),
    .A2(_08172_),
    .A3(net20784),
    .ZN(_08173_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17034_ (.A1(_08165_),
    .A2(_08173_),
    .B(_08030_),
    .ZN(_08174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17035_ (.A1(_08159_),
    .A2(_08174_),
    .ZN(_08175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17036_ (.A1(_08148_),
    .A2(_08175_),
    .A3(_08075_),
    .ZN(_08176_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17037_ (.A1(net20777),
    .A2(net20387),
    .Z(_08177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17038_ (.A1(_08177_),
    .A2(net20794),
    .B(net20782),
    .ZN(_08178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17039_ (.A1(_08178_),
    .A2(_08172_),
    .B(net20537),
    .ZN(_08179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17040_ (.A1(_08060_),
    .A2(net20528),
    .ZN(_08180_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17041_ (.A1(_08180_),
    .A2(net20785),
    .A3(_08164_),
    .ZN(_08181_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17042_ (.A1(_08179_),
    .A2(_08181_),
    .B(_08030_),
    .ZN(_08182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17043_ (.A1(_07997_),
    .A2(net20365),
    .ZN(_08183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17044_ (.A1(net20833),
    .A2(net20835),
    .ZN(_08184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17045_ (.A1(_08056_),
    .A2(_08184_),
    .A3(net20613),
    .ZN(_08185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17046_ (.A1(_08183_),
    .A2(net20542),
    .A3(_08185_),
    .ZN(_08186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17047_ (.A1(_08094_),
    .A2(net20352),
    .ZN(_08187_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17048_ (.A1(net20347),
    .A2(net20797),
    .A3(net20148),
    .ZN(_08188_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17049_ (.A1(_08187_),
    .A2(_08188_),
    .A3(net20782),
    .ZN(_08189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17050_ (.A1(_08186_),
    .A2(_08189_),
    .ZN(_08190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17051_ (.A1(_08190_),
    .A2(net20537),
    .ZN(_08191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17052_ (.A1(_08182_),
    .A2(_08191_),
    .B(_08075_),
    .ZN(_08192_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17053_ (.I(_08037_),
    .ZN(_08193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17054_ (.A1(_08067_),
    .A2(net20794),
    .ZN(_08194_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17055_ (.A1(net20131),
    .A2(net20141),
    .B1(_08194_),
    .B2(_08149_),
    .ZN(_08195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17056_ (.A1(_08085_),
    .A2(_07998_),
    .ZN(_08196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17057_ (.A1(net20608),
    .A2(net20555),
    .Z(_08197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17058_ (.A1(_08197_),
    .A2(_08105_),
    .ZN(_08198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17059_ (.A1(_08196_),
    .A2(net20552),
    .A3(_08198_),
    .ZN(_08199_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17060_ (.A1(_08195_),
    .A2(net20552),
    .B(_08199_),
    .C(net20789),
    .ZN(_08200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17061_ (.A1(net20794),
    .A2(net20792),
    .ZN(_08201_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17062_ (.A1(_08201_),
    .A2(_07976_),
    .Z(_08202_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17063_ (.A1(net20794),
    .A2(_15558_[0]),
    .Z(_08203_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17064_ (.A1(_08202_),
    .A2(_08203_),
    .Z(_08204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17065_ (.A1(_08101_),
    .A2(net20782),
    .Z(_08205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17066_ (.A1(_08204_),
    .A2(_08205_),
    .B(net20789),
    .ZN(_08206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17067_ (.A1(_08106_),
    .A2(net20796),
    .ZN(_08207_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17068_ (.A1(_08207_),
    .A2(net20542),
    .A3(_08101_),
    .Z(_08208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17069_ (.A1(_08045_),
    .A2(net20365),
    .ZN(_08209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17070_ (.A1(_08208_),
    .A2(_08209_),
    .ZN(_08210_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17071_ (.A1(_08206_),
    .A2(_08210_),
    .B(net20846),
    .ZN(_08211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17072_ (.A1(_08200_),
    .A2(_08211_),
    .ZN(_08212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17073_ (.A1(_08192_),
    .A2(_08212_),
    .ZN(_08213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17074_ (.A1(_08176_),
    .A2(_08213_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17075_ (.A1(_08056_),
    .A2(net20794),
    .A3(net20137),
    .Z(_08214_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17076_ (.A1(net20366),
    .A2(net20604),
    .A3(net20522),
    .Z(_08215_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17077_ (.A1(net19911),
    .A2(_08215_),
    .B(net20548),
    .ZN(_08216_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17078_ (.I(_08096_),
    .ZN(_08217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17079_ (.A1(net20346),
    .A2(net19910),
    .A3(net20604),
    .ZN(_08218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17080_ (.A1(net20863),
    .A2(net20623),
    .A3(net21515),
    .ZN(_08219_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17081_ (.A1(_07996_),
    .A2(net20795),
    .A3(_08219_),
    .ZN(_08220_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17082_ (.A1(_08218_),
    .A2(net20782),
    .A3(net20343),
    .ZN(_08221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17083_ (.A1(_08216_),
    .A2(_08221_),
    .ZN(_08222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17084_ (.A1(_08222_),
    .A2(net20789),
    .ZN(_08223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17085_ (.A1(net19909),
    .A2(net20353),
    .ZN(_08224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17086_ (.A1(_08224_),
    .A2(net20795),
    .ZN(_08225_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17087_ (.A1(net20554),
    .A2(net20355),
    .ZN(_08226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17088_ (.A1(_08226_),
    .A2(net20602),
    .A3(net20528),
    .ZN(_08227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17089_ (.A1(_08225_),
    .A2(_08227_),
    .A3(net20548),
    .ZN(_08228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17090_ (.A1(net20140),
    .A2(net20795),
    .B(net20548),
    .ZN(_08229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17091_ (.A1(_08226_),
    .A2(net20604),
    .A3(_08056_),
    .ZN(_08230_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17092_ (.A1(_08219_),
    .A2(net20604),
    .Z(_08231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17093_ (.A1(_08229_),
    .A2(_08230_),
    .A3(_08231_),
    .ZN(_08232_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17094_ (.A1(_08228_),
    .A2(_08232_),
    .A3(net20532),
    .ZN(_08233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17095_ (.A1(_08223_),
    .A2(net20846),
    .A3(_08233_),
    .ZN(_08234_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17096_ (.I(_08087_),
    .ZN(_08235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17097_ (.A1(_08100_),
    .A2(net20606),
    .ZN(_08236_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17098_ (.A1(_08236_),
    .A2(_08106_),
    .B(net20542),
    .ZN(_08237_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17099_ (.A1(_08235_),
    .A2(net19908),
    .ZN(_08238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17100_ (.A1(_08065_),
    .A2(net20523),
    .ZN(_08239_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17101_ (.A1(net20144),
    .A2(net20357),
    .A3(net20794),
    .ZN(_08240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17102_ (.A1(_08239_),
    .A2(_08240_),
    .B(net20549),
    .ZN(_08241_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17103_ (.A1(_08238_),
    .A2(_08241_),
    .B(net20532),
    .ZN(_08242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17104_ (.A1(net20554),
    .A2(_15555_[0]),
    .ZN(_08243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17105_ (.I(_08243_),
    .ZN(_08244_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17106_ (.I(_07996_),
    .ZN(_08245_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17107_ (.A1(net20130),
    .A2(net20342),
    .B(net20605),
    .ZN(_08246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17108_ (.A1(_08005_),
    .A2(net20794),
    .A3(net20366),
    .ZN(_08247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17109_ (.A1(_08246_),
    .A2(net20782),
    .A3(_08247_),
    .ZN(_08248_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17110_ (.A1(net20147),
    .A2(net20543),
    .Z(_08249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17111_ (.A1(net20132),
    .A2(net20361),
    .ZN(_08250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17112_ (.A1(_08249_),
    .A2(_08250_),
    .B(net20536),
    .ZN(_08251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17113_ (.A1(_08248_),
    .A2(_08251_),
    .ZN(_08252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17114_ (.A1(_08242_),
    .A2(_08030_),
    .A3(_08252_),
    .ZN(_08253_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17115_ (.A1(_08234_),
    .A2(_08253_),
    .A3(_08075_),
    .ZN(_08254_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17116_ (.A1(_08245_),
    .A2(_15560_[0]),
    .B(net20605),
    .ZN(_08255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17117_ (.A1(net20142),
    .A2(_08255_),
    .B(net20549),
    .ZN(_08256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17118_ (.A1(_08114_),
    .A2(net20606),
    .ZN(_08257_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17119_ (.A1(_08257_),
    .A2(_08012_),
    .Z(_08258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17120_ (.A1(net20797),
    .A2(_15565_[0]),
    .ZN(_08259_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17664 (.I(_05480_),
    .Z(net17664));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17122_ (.A1(_08258_),
    .A2(_08259_),
    .B(net20782),
    .ZN(_08261_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17123_ (.A1(_08256_),
    .A2(_08261_),
    .B(net20846),
    .ZN(_08262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17124_ (.A1(_08094_),
    .A2(_08226_),
    .ZN(_08263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17125_ (.A1(_08263_),
    .A2(_08019_),
    .B(net20846),
    .ZN(_08264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17126_ (.A1(net20132),
    .A2(net20540),
    .ZN(_08265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17127_ (.A1(_08143_),
    .A2(_08265_),
    .A3(net20787),
    .ZN(_08266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17128_ (.A1(_08264_),
    .A2(_08266_),
    .B(net20533),
    .ZN(_08267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17129_ (.A1(_08262_),
    .A2(_08267_),
    .ZN(_08268_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17130_ (.A1(net20795),
    .A2(_15563_[0]),
    .Z(_08269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17131_ (.A1(_08269_),
    .A2(_08249_),
    .B(net20846),
    .ZN(_08270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17132_ (.A1(net20794),
    .A2(net20160),
    .ZN(_08271_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17133_ (.A1(_08239_),
    .A2(net20787),
    .A3(_08271_),
    .ZN(_08272_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17134_ (.A1(_08270_),
    .A2(_08272_),
    .B(net20789),
    .ZN(_08273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17135_ (.A1(net20151),
    .A2(_08084_),
    .ZN(_08274_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17136_ (.A1(_08274_),
    .A2(net20794),
    .ZN(_08275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17137_ (.A1(_07982_),
    .A2(net20610),
    .ZN(_08276_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17138_ (.A1(_08154_),
    .A2(_08275_),
    .A3(_08276_),
    .ZN(_08277_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17139_ (.A1(_07998_),
    .A2(net20524),
    .A3(net20613),
    .ZN(_08278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17140_ (.A1(net20794),
    .A2(net20134),
    .ZN(_08279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17141_ (.A1(_08278_),
    .A2(net20549),
    .A3(_08279_),
    .ZN(_08280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17142_ (.A1(_08277_),
    .A2(net20846),
    .A3(_08280_),
    .ZN(_08281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17143_ (.A1(_08273_),
    .A2(_08281_),
    .ZN(_08282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17144_ (.A1(_08268_),
    .A2(net20845),
    .A3(_08282_),
    .ZN(_08283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17145_ (.A1(_08254_),
    .A2(_08283_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17146_ (.I(_08214_),
    .ZN(_08284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17147_ (.A1(net20140),
    .A2(_07330_),
    .ZN(_08285_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17148_ (.A1(_08284_),
    .A2(net20788),
    .A3(_08285_),
    .ZN(_08286_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17149_ (.I(_08070_),
    .ZN(_08287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17150_ (.A1(_08287_),
    .A2(net20366),
    .ZN(_08288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17151_ (.A1(_08060_),
    .A2(net20540),
    .ZN(_08289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17152_ (.A1(_08288_),
    .A2(net20537),
    .A3(_08289_),
    .ZN(_08290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17153_ (.A1(_08286_),
    .A2(_08290_),
    .ZN(_08291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17154_ (.A1(_08291_),
    .A2(net20542),
    .ZN(_08292_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17155_ (.A1(_08142_),
    .A2(net20523),
    .Z(_08293_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17156_ (.I(_08013_),
    .ZN(_08294_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17157_ (.A1(_08293_),
    .A2(_08294_),
    .B(net20536),
    .ZN(_08295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17158_ (.A1(_08109_),
    .A2(net20782),
    .Z(_08296_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17159_ (.A1(_08027_),
    .A2(net20366),
    .A3(_07330_),
    .Z(_08297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17160_ (.A1(_08296_),
    .A2(_08297_),
    .Z(_08298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17161_ (.A1(_08298_),
    .A2(_08295_),
    .B(net20846),
    .ZN(_08299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17162_ (.A1(_08292_),
    .A2(_08299_),
    .ZN(_08300_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17163_ (.A1(_08193_),
    .A2(_08096_),
    .B(net20614),
    .ZN(_08301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17164_ (.A1(_07990_),
    .A2(net20356),
    .ZN(_08302_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17165_ (.A1(_08301_),
    .A2(_08302_),
    .A3(net20782),
    .ZN(_08303_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17166_ (.A1(_08196_),
    .A2(_08120_),
    .A3(net20542),
    .ZN(_08304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17167_ (.A1(_08303_),
    .A2(_08304_),
    .ZN(_08305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17168_ (.A1(_08305_),
    .A2(net20790),
    .ZN(_08306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17169_ (.A1(_08113_),
    .A2(_07996_),
    .ZN(_08307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17170_ (.A1(_08143_),
    .A2(_08307_),
    .ZN(_08308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17171_ (.A1(_08308_),
    .A2(net20542),
    .ZN(_08309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17172_ (.A1(_08220_),
    .A2(net20782),
    .B(net20788),
    .ZN(_08310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17173_ (.A1(_08309_),
    .A2(_08310_),
    .B(_08030_),
    .ZN(_08311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17174_ (.A1(_08306_),
    .A2(_08311_),
    .ZN(_08312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17175_ (.A1(_08300_),
    .A2(_08312_),
    .ZN(_08313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17176_ (.A1(_08313_),
    .A2(_08075_),
    .ZN(_08314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17177_ (.A1(_08038_),
    .A2(net20794),
    .Z(_08315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17178_ (.A1(_08315_),
    .A2(net20365),
    .ZN(_08316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17179_ (.A1(net20555),
    .A2(_08105_),
    .ZN(_08317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17180_ (.A1(_08317_),
    .A2(_07981_),
    .ZN(_08318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17181_ (.A1(_08318_),
    .A2(net20608),
    .ZN(_08319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17182_ (.A1(_08316_),
    .A2(_08319_),
    .ZN(_08320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17183_ (.A1(_08320_),
    .A2(net20547),
    .ZN(_08321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17184_ (.A1(_07990_),
    .A2(_08023_),
    .ZN(_08322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17185_ (.A1(_08322_),
    .A2(_08002_),
    .A3(net20782),
    .ZN(_08323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17186_ (.A1(_08321_),
    .A2(_08323_),
    .ZN(_08324_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17187_ (.A1(_08324_),
    .A2(net20790),
    .ZN(_08325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17188_ (.A1(net20348),
    .A2(_07998_),
    .ZN(_08326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17189_ (.A1(_08326_),
    .A2(net20802),
    .ZN(_08327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17190_ (.A1(_08064_),
    .A2(net20542),
    .Z(_08328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17191_ (.A1(_08327_),
    .A2(_08328_),
    .B(net20790),
    .ZN(_08329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17192_ (.A1(_08111_),
    .A2(net20794),
    .ZN(_08330_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17193_ (.I(_08330_),
    .ZN(_08331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17194_ (.A1(_08331_),
    .A2(net20538),
    .ZN(_08332_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17195_ (.A1(_08180_),
    .A2(_08332_),
    .A3(net20785),
    .ZN(_08333_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17196_ (.A1(_08329_),
    .A2(_08333_),
    .B(_08030_),
    .ZN(_08334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17197_ (.A1(_08325_),
    .A2(_08334_),
    .B(_08075_),
    .ZN(_08335_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17198_ (.A1(_08155_),
    .A2(net20782),
    .Z(_08336_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17199_ (.A1(net20133),
    .A2(_07982_),
    .B(net20799),
    .ZN(_08337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17200_ (.A1(_08336_),
    .A2(_08337_),
    .A3(_08013_),
    .ZN(_08338_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17201_ (.I(_08006_),
    .ZN(_08339_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17202_ (.A1(_08339_),
    .A2(net20608),
    .A3(_08033_),
    .Z(_08340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17203_ (.A1(_08045_),
    .A2(_08226_),
    .ZN(_08341_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17204_ (.A1(_08340_),
    .A2(net20544),
    .A3(_08341_),
    .ZN(_08342_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17205_ (.A1(_08338_),
    .A2(_08342_),
    .A3(net20789),
    .ZN(_08343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17206_ (.A1(_08094_),
    .A2(_08138_),
    .ZN(_08344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17207_ (.A1(_08327_),
    .A2(_08344_),
    .B(net20782),
    .ZN(_08345_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17208_ (.A1(_08245_),
    .A2(_15560_[0]),
    .ZN(_08346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17209_ (.A1(net20782),
    .A2(_08013_),
    .ZN(_08347_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17210_ (.A1(net20794),
    .A2(_08346_),
    .B(_08347_),
    .ZN(_08348_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17211_ (.A1(_08348_),
    .A2(_08345_),
    .B(net20536),
    .ZN(_08349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17212_ (.A1(_08343_),
    .A2(_08030_),
    .A3(_08349_),
    .ZN(_08350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17213_ (.A1(_08335_),
    .A2(_08350_),
    .ZN(_08351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17214_ (.A1(_08351_),
    .A2(_08314_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17215_ (.A1(_08078_),
    .A2(net20551),
    .A3(_08002_),
    .ZN(_08352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17216_ (.A1(_08048_),
    .A2(_08184_),
    .ZN(_08353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17217_ (.A1(net20341),
    .A2(net20794),
    .ZN(_08354_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17218_ (.A1(_08354_),
    .A2(_08307_),
    .A3(net20782),
    .ZN(_08355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17219_ (.A1(_08352_),
    .A2(net20536),
    .A3(_08355_),
    .ZN(_08356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17220_ (.A1(_08113_),
    .A2(net20527),
    .ZN(_08357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17221_ (.A1(_08108_),
    .A2(_08357_),
    .ZN(_08358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17222_ (.A1(net20799),
    .A2(net20521),
    .ZN(_08359_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17223_ (.A1(net20345),
    .A2(net20799),
    .B(net20551),
    .C(_08359_),
    .ZN(_08360_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17224_ (.A1(_08358_),
    .A2(_08360_),
    .A3(net20789),
    .ZN(_08361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17225_ (.A1(_08356_),
    .A2(_08030_),
    .A3(_08361_),
    .ZN(_08362_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17226_ (.A1(_08194_),
    .A2(net20345),
    .Z(_08363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17227_ (.A1(_08099_),
    .A2(_08363_),
    .ZN(_08364_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17228_ (.A1(_08170_),
    .A2(net20782),
    .Z(_08365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17229_ (.A1(_08168_),
    .A2(net20794),
    .ZN(_08366_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17230_ (.A1(_08365_),
    .A2(_08366_),
    .B(net20532),
    .ZN(_08367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17231_ (.A1(_08364_),
    .A2(_08367_),
    .ZN(_08368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17232_ (.A1(_07997_),
    .A2(net20358),
    .ZN(_08369_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17233_ (.A1(_08197_),
    .A2(net20782),
    .ZN(_08370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17234_ (.A1(_08369_),
    .A2(_08370_),
    .B(net20789),
    .ZN(_08371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17235_ (.A1(_08016_),
    .A2(net20797),
    .B(net20542),
    .ZN(_08372_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17236_ (.A1(_08139_),
    .A2(_08372_),
    .A3(_08034_),
    .ZN(_08373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17237_ (.A1(_08371_),
    .A2(_08373_),
    .ZN(_08374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17238_ (.A1(_08368_),
    .A2(_08374_),
    .A3(net20846),
    .ZN(_08375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17239_ (.A1(_08362_),
    .A2(_08075_),
    .A3(_08375_),
    .ZN(_08376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17240_ (.A1(_08005_),
    .A2(net20148),
    .ZN(_08377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17241_ (.A1(_08377_),
    .A2(net20606),
    .ZN(_08378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17242_ (.A1(_08208_),
    .A2(_08378_),
    .ZN(_08379_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17243_ (.A1(net20531),
    .A2(net20129),
    .B(_08240_),
    .C(net20782),
    .ZN(_08380_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17244_ (.A1(_08379_),
    .A2(_08380_),
    .A3(net20535),
    .ZN(_08381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17245_ (.A1(_08153_),
    .A2(_08217_),
    .Z(_08382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17246_ (.A1(_08205_),
    .A2(_08382_),
    .B(net20533),
    .ZN(_08383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17247_ (.A1(_08167_),
    .A2(net20365),
    .ZN(_08384_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17248_ (.A1(_08384_),
    .A2(_08115_),
    .A3(net20550),
    .ZN(_08385_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17249_ (.A1(_08383_),
    .A2(_08385_),
    .B(net20846),
    .ZN(_08386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17250_ (.A1(_08381_),
    .A2(_08386_),
    .ZN(_08387_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17251_ (.A1(_08245_),
    .A2(net20159),
    .B(net20605),
    .ZN(_08388_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17252_ (.A1(_08133_),
    .A2(_08388_),
    .A3(net20549),
    .ZN(_08389_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17253_ (.A1(net20362),
    .A2(net20548),
    .ZN(_08390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17254_ (.A1(_08390_),
    .A2(net19912),
    .B(net20532),
    .ZN(_08391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17255_ (.A1(_08389_),
    .A2(_08391_),
    .B(_08030_),
    .ZN(_08392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17256_ (.A1(_08353_),
    .A2(net20605),
    .Z(_08393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17257_ (.A1(_08274_),
    .A2(net20605),
    .ZN(_08394_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17258_ (.A1(_08393_),
    .A2(_08394_),
    .A3(net20782),
    .ZN(_08395_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17259_ (.A1(_08137_),
    .A2(net20549),
    .A3(_08278_),
    .ZN(_08396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17260_ (.A1(_08395_),
    .A2(_08396_),
    .A3(net20534),
    .ZN(_08397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17261_ (.A1(_08392_),
    .A2(_08397_),
    .ZN(_08398_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17262_ (.A1(_08387_),
    .A2(net20845),
    .A3(_08398_),
    .ZN(_08399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17263_ (.A1(_08376_),
    .A2(_08399_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17264_ (.A1(net20610),
    .A2(net20833),
    .ZN(_08400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17265_ (.A1(_07999_),
    .A2(net20545),
    .A3(_08400_),
    .ZN(_08401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17266_ (.A1(_08331_),
    .A2(net20528),
    .ZN(_08402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17267_ (.A1(_08065_),
    .A2(net20366),
    .ZN(_08403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17268_ (.A1(_08402_),
    .A2(_08403_),
    .A3(net20786),
    .ZN(_08404_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17269_ (.A1(_08401_),
    .A2(_08404_),
    .A3(net20790),
    .ZN(_08405_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17270_ (.A1(_08024_),
    .A2(net20609),
    .B(net20547),
    .ZN(_08406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17271_ (.A1(_08315_),
    .A2(net20356),
    .ZN(_08407_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17272_ (.A1(_08406_),
    .A2(_08407_),
    .B(net20790),
    .ZN(_08408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17273_ (.A1(_08132_),
    .A2(_08226_),
    .ZN(_08409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17274_ (.A1(_08099_),
    .A2(_08409_),
    .ZN(_08410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17275_ (.A1(_08408_),
    .A2(_08410_),
    .ZN(_08411_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17276_ (.A1(_08405_),
    .A2(_08411_),
    .A3(_08075_),
    .ZN(_08412_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17277_ (.I(_07990_),
    .ZN(_08413_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17278_ (.A1(_08301_),
    .A2(net20546),
    .A3(_08413_),
    .ZN(_08414_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17279_ (.A1(_08194_),
    .A2(net20782),
    .A3(_08317_),
    .Z(_08415_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17280_ (.A1(_08415_),
    .A2(net20790),
    .ZN(_08416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17281_ (.A1(_08414_),
    .A2(_08416_),
    .B(_08075_),
    .ZN(_08417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17282_ (.A1(_08079_),
    .A2(net20357),
    .ZN(_08418_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17283_ (.A1(_08036_),
    .A2(_08418_),
    .A3(_08041_),
    .ZN(_08419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17284_ (.A1(net20540),
    .A2(net20602),
    .Z(_08420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17285_ (.A1(_08420_),
    .A2(_08226_),
    .ZN(_08421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17286_ (.A1(_08331_),
    .A2(net20351),
    .ZN(_08422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17287_ (.A1(_08421_),
    .A2(net20786),
    .A3(_08422_),
    .ZN(_08423_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17288_ (.A1(_08419_),
    .A2(_08423_),
    .A3(net20790),
    .ZN(_08424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17289_ (.A1(_08417_),
    .A2(_08424_),
    .ZN(_08425_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17290_ (.A1(_08412_),
    .A2(_08425_),
    .A3(net20846),
    .ZN(_08426_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17291_ (.I(_08366_),
    .ZN(_08427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17292_ (.A1(_08427_),
    .A2(net20523),
    .ZN(_08428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17293_ (.A1(_08428_),
    .A2(_08154_),
    .B(net20789),
    .ZN(_08429_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17294_ (.A1(net20151),
    .A2(net20366),
    .Z(_08430_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17295_ (.A1(_08430_),
    .A2(net20794),
    .B(net20549),
    .C(_08231_),
    .ZN(_08431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17296_ (.A1(_08429_),
    .A2(_08431_),
    .ZN(_08432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17297_ (.A1(net20801),
    .A2(net20833),
    .ZN(_08433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17298_ (.A1(_08433_),
    .A2(net20835),
    .ZN(_08434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17299_ (.A1(_08036_),
    .A2(_08434_),
    .B(net20536),
    .ZN(_08435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17300_ (.A1(_08023_),
    .A2(_08163_),
    .ZN(_08436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17301_ (.A1(_08436_),
    .A2(net20609),
    .ZN(_08437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17302_ (.A1(net20364),
    .A2(net20667),
    .ZN(_08438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17303_ (.A1(_08438_),
    .A2(net20801),
    .ZN(_08439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17304_ (.A1(_08437_),
    .A2(_08439_),
    .A3(net20782),
    .ZN(_08440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17305_ (.A1(_08435_),
    .A2(_08440_),
    .ZN(_08441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17306_ (.A1(_08432_),
    .A2(_08441_),
    .A3(net20845),
    .ZN(_08442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17307_ (.A1(_08094_),
    .A2(net20354),
    .ZN(_08443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17308_ (.A1(net20538),
    .A2(net20356),
    .A3(net20800),
    .ZN(_08444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17309_ (.A1(_08443_),
    .A2(net20782),
    .A3(_08444_),
    .ZN(_08445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17310_ (.A1(net20602),
    .A2(_07980_),
    .Z(_08446_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17311_ (.A1(_08315_),
    .A2(net20782),
    .A3(_08446_),
    .Z(_08447_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17312_ (.A1(_08445_),
    .A2(_08447_),
    .A3(net20537),
    .ZN(_08448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17313_ (.A1(_08055_),
    .A2(net20530),
    .ZN(_08449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17314_ (.I(_08420_),
    .ZN(_08450_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17315_ (.A1(_08449_),
    .A2(_08450_),
    .A3(net20543),
    .ZN(_08451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17316_ (.A1(_08205_),
    .A2(net20146),
    .ZN(_08452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17317_ (.A1(_08451_),
    .A2(_08452_),
    .A3(net20790),
    .ZN(_08453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17318_ (.A1(_08448_),
    .A2(_08075_),
    .A3(_08453_),
    .ZN(_08454_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17319_ (.A1(_08442_),
    .A2(_08454_),
    .A3(_08030_),
    .ZN(_08455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17320_ (.A1(_08426_),
    .A2(_08455_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17321_ (.A1(_08060_),
    .A2(net20538),
    .ZN(_08456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17322_ (.A1(_08456_),
    .A2(_08150_),
    .A3(net20782),
    .ZN(_08457_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17323_ (.A1(net20794),
    .A2(_15559_[0]),
    .Z(_08458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17324_ (.A1(_08402_),
    .A2(net20543),
    .A3(_08458_),
    .ZN(_08459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17325_ (.A1(_08457_),
    .A2(_08459_),
    .ZN(_08460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17326_ (.A1(_08460_),
    .A2(net20790),
    .ZN(_08461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17327_ (.A1(_08357_),
    .A2(net20135),
    .ZN(_08462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17328_ (.A1(_08462_),
    .A2(net20784),
    .ZN(_08463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17329_ (.A1(_08237_),
    .A2(net20537),
    .Z(_08464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17330_ (.A1(_08463_),
    .A2(_08464_),
    .ZN(_08465_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17331_ (.A1(_08461_),
    .A2(_08030_),
    .A3(_08465_),
    .ZN(_08466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17332_ (.A1(_08339_),
    .A2(net20800),
    .ZN(_08467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17333_ (.A1(_08301_),
    .A2(_08467_),
    .ZN(_08468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17334_ (.A1(_08468_),
    .A2(net20546),
    .ZN(_08469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17335_ (.A1(_08057_),
    .A2(_08203_),
    .ZN(_08470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17336_ (.A1(_08470_),
    .A2(net20785),
    .ZN(_08471_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17337_ (.A1(_08469_),
    .A2(net20537),
    .A3(_08471_),
    .ZN(_08472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17338_ (.A1(_07998_),
    .A2(net20608),
    .ZN(_08473_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17339_ (.A1(_08473_),
    .A2(_08149_),
    .Z(_08474_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17340_ (.A1(_08048_),
    .A2(net20794),
    .Z(_08475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17341_ (.A1(_08475_),
    .A2(net20128),
    .ZN(_08476_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17342_ (.A1(_08474_),
    .A2(_08476_),
    .A3(net20547),
    .ZN(_08477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17343_ (.A1(_08473_),
    .A2(_08166_),
    .ZN(_08478_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17344_ (.A1(net20349),
    .A2(net20782),
    .Z(_08479_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17345_ (.A1(_08478_),
    .A2(_08479_),
    .B(net20537),
    .ZN(_08480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17346_ (.A1(_08477_),
    .A2(_08480_),
    .B(_08030_),
    .ZN(_08481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17347_ (.A1(_08472_),
    .A2(_08481_),
    .ZN(_08482_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17348_ (.A1(_08466_),
    .A2(_08482_),
    .ZN(_08483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17349_ (.A1(_08483_),
    .A2(_08075_),
    .ZN(_08484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17350_ (.A1(_08243_),
    .A2(_08217_),
    .ZN(_08485_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17351_ (.A1(_08485_),
    .A2(net20605),
    .ZN(_08486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17352_ (.A1(_08486_),
    .A2(_08372_),
    .B(net20534),
    .ZN(_08487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17353_ (.A1(_08353_),
    .A2(net20605),
    .ZN(_08488_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17354_ (.A1(_08488_),
    .A2(net20549),
    .A3(net20520),
    .ZN(_08489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17355_ (.A1(_08487_),
    .A2(_08489_),
    .B(_08030_),
    .ZN(_08490_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17356_ (.A1(_07997_),
    .A2(net20522),
    .ZN(_08491_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17357_ (.A1(_08301_),
    .A2(_08491_),
    .A3(net20785),
    .ZN(_08492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17358_ (.A1(net20363),
    .A2(net20610),
    .B(net20782),
    .ZN(_08493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17359_ (.A1(_08331_),
    .A2(net20360),
    .ZN(_08494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17360_ (.A1(_08197_),
    .A2(net20521),
    .ZN(_08495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17361_ (.A1(_08493_),
    .A2(_08494_),
    .A3(_08495_),
    .ZN(_08496_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17362_ (.A1(_08492_),
    .A2(net20537),
    .A3(_08496_),
    .ZN(_08497_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17363_ (.A1(_08490_),
    .A2(_08497_),
    .B(_08075_),
    .ZN(_08498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17364_ (.A1(_08005_),
    .A2(net20351),
    .ZN(_08499_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17365_ (.A1(net20800),
    .A2(_08499_),
    .B(_08025_),
    .C(net20786),
    .ZN(_08500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17366_ (.A1(net20350),
    .A2(net20612),
    .A3(net20351),
    .ZN(_08501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17367_ (.A1(_08491_),
    .A2(net20546),
    .A3(_08501_),
    .ZN(_08502_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17368_ (.A1(_08500_),
    .A2(net20537),
    .A3(_08502_),
    .ZN(_08503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17369_ (.A1(_08427_),
    .A2(net20538),
    .ZN(_08504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17370_ (.A1(_08065_),
    .A2(net20528),
    .ZN(_08505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17371_ (.A1(_08504_),
    .A2(net20543),
    .A3(_08505_),
    .ZN(_08506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17372_ (.A1(net20150),
    .A2(net20359),
    .ZN(_08507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17373_ (.A1(_08507_),
    .A2(net20783),
    .A3(_08269_),
    .ZN(_08508_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17374_ (.A1(_08506_),
    .A2(_08508_),
    .A3(net20790),
    .ZN(_08509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17375_ (.A1(_08503_),
    .A2(_08509_),
    .A3(_08030_),
    .ZN(_08510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17376_ (.A1(_08498_),
    .A2(_08510_),
    .ZN(_08511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17377_ (.A1(_08484_),
    .A2(_08511_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17378_ (.A1(_08287_),
    .A2(net20351),
    .ZN(_08512_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17379_ (.A1(_08336_),
    .A2(_08512_),
    .A3(_08495_),
    .ZN(_08513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17380_ (.A1(_08166_),
    .A2(net20542),
    .Z(_08514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17381_ (.A1(_08514_),
    .A2(_08357_),
    .B(net20536),
    .ZN(_08515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17382_ (.A1(_08513_),
    .A2(_08515_),
    .B(_08030_),
    .ZN(_08516_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17383_ (.A1(_08288_),
    .A2(net20783),
    .A3(_08209_),
    .ZN(_08517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17384_ (.A1(_08255_),
    .A2(_08494_),
    .A3(net20550),
    .ZN(_08518_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17385_ (.A1(_08517_),
    .A2(_08518_),
    .A3(net20536),
    .ZN(_08519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17386_ (.A1(_08516_),
    .A2(_08519_),
    .ZN(_08520_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17387_ (.A1(_08006_),
    .A2(_07993_),
    .A3(net20797),
    .ZN(_08521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17388_ (.A1(_08521_),
    .A2(_08257_),
    .ZN(_08522_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17389_ (.A1(_08522_),
    .A2(net20782),
    .ZN(_08523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17390_ (.A1(_08163_),
    .A2(net20608),
    .ZN(_08524_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17391_ (.A1(_08413_),
    .A2(_08524_),
    .A3(net20546),
    .ZN(_08525_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17392_ (.A1(_08523_),
    .A2(_08525_),
    .ZN(_08526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17393_ (.A1(_08526_),
    .A2(net20537),
    .ZN(_08527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17394_ (.A1(_08420_),
    .A2(_08138_),
    .ZN(_08528_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17395_ (.A1(_08433_),
    .A2(net20782),
    .Z(_08529_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17396_ (.A1(_08528_),
    .A2(_08529_),
    .B(net20536),
    .ZN(_08530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17397_ (.A1(_08475_),
    .A2(net20541),
    .ZN(_08531_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17398_ (.A1(_08531_),
    .A2(net20544),
    .A3(_08278_),
    .ZN(_08532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17399_ (.A1(_08530_),
    .A2(_08532_),
    .ZN(_08533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17400_ (.A1(_08527_),
    .A2(_08533_),
    .A3(_08030_),
    .ZN(_08534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17401_ (.A1(_08520_),
    .A2(_08534_),
    .A3(_08075_),
    .ZN(_08535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17402_ (.A1(_08085_),
    .A2(net20541),
    .ZN(_08536_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17403_ (.A1(_08536_),
    .A2(net20782),
    .A3(_08307_),
    .ZN(_08537_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17404_ (.A1(net20539),
    .A2(net20354),
    .A3(net20614),
    .ZN(_08538_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17405_ (.A1(_08119_),
    .A2(net20541),
    .A3(net20798),
    .ZN(_08539_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17406_ (.A1(_08538_),
    .A2(_08539_),
    .A3(net20542),
    .ZN(_08540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17407_ (.A1(_08537_),
    .A2(_08540_),
    .A3(net20789),
    .ZN(_08541_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17408_ (.A1(net20796),
    .A2(net20387),
    .ZN(_08542_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17409_ (.A1(_08488_),
    .A2(net20782),
    .A3(_08542_),
    .ZN(_08543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17410_ (.A1(net20531),
    .A2(net20606),
    .B(net20782),
    .ZN(_08544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17411_ (.A1(_08244_),
    .A2(net20794),
    .ZN(_08545_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17412_ (.A1(_08544_),
    .A2(_08545_),
    .A3(net20148),
    .ZN(_08546_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17413_ (.A1(_08543_),
    .A2(_08546_),
    .A3(net20535),
    .ZN(_08547_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17414_ (.A1(_08541_),
    .A2(_08547_),
    .A3(net20846),
    .ZN(_08548_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17415_ (.A1(net20539),
    .A2(net20365),
    .A3(net20614),
    .ZN(_08549_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _17416_ (.A1(net20782),
    .A2(_08150_),
    .A3(_08549_),
    .A4(_08259_),
    .ZN(_08550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17417_ (.A1(_07330_),
    .A2(_15569_[0]),
    .ZN(_08551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17418_ (.A1(_08551_),
    .A2(net20542),
    .ZN(_08552_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17419_ (.A1(_08552_),
    .A2(_08097_),
    .ZN(_08553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17420_ (.A1(net20149),
    .A2(net20798),
    .ZN(_08554_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17421_ (.A1(_08553_),
    .A2(_08554_),
    .B(net20789),
    .ZN(_08555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17422_ (.A1(_08550_),
    .A2(_08555_),
    .ZN(_08556_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17423_ (.A1(net20625),
    .A2(net20794),
    .B(net20542),
    .ZN(_08557_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17424_ (.I(_08557_),
    .ZN(_08558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17425_ (.A1(_08558_),
    .A2(_08545_),
    .B(net20534),
    .ZN(_08559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17426_ (.A1(_08139_),
    .A2(_08108_),
    .A3(_08034_),
    .ZN(_08560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17427_ (.A1(_08559_),
    .A2(_08560_),
    .ZN(_08561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17428_ (.A1(_08556_),
    .A2(_08561_),
    .A3(_08030_),
    .ZN(_08562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17429_ (.A1(_08548_),
    .A2(_08562_),
    .A3(net20845),
    .ZN(_08563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17430_ (.A1(_08535_),
    .A2(_08563_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17431_ (.A1(net21518),
    .A2(_07609_),
    .B(_07612_),
    .ZN(_15571_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17432_ (.A1(_07618_),
    .A2(net21524),
    .B(_07620_),
    .ZN(_08564_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17662 (.I(_05497_),
    .Z(net17662));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17434_ (.A1(net21518),
    .A2(_07601_),
    .B(_07604_),
    .ZN(_15572_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17435_ (.A1(net20743),
    .A2(net20823),
    .ZN(_08565_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17436_ (.I(_08565_),
    .ZN(_08566_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17667 (.I(_05424_),
    .Z(net17667));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17438_ (.A1(_08566_),
    .A2(net20721),
    .ZN(_08568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17439_ (.A1(net20740),
    .A2(_15589_[0]),
    .Z(_08569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17440_ (.A1(_08569_),
    .A2(net20721),
    .ZN(_08570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17441_ (.A1(_08568_),
    .A2(_08570_),
    .ZN(_08571_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17442_ (.I(_08571_),
    .ZN(_08572_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17672 (.I(_05374_),
    .Z(net17672));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17680 (.I(_05003_),
    .Z(net17680));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17445_ (.A1(net20827),
    .A2(net20821),
    .ZN(_08575_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _17446_ (.I(_08575_),
    .ZN(_08576_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17447_ (.I(_15573_[0]),
    .ZN(_08577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17448_ (.A1(net20740),
    .A2(_08577_),
    .ZN(_08578_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17449_ (.I(_08578_),
    .ZN(_08579_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17661 (.I(_05539_),
    .Z(net17661));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17451_ (.A1(_08576_),
    .A2(_08579_),
    .B(net20580),
    .ZN(_08581_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17452_ (.A1(_08572_),
    .A2(net20854),
    .A3(_08581_),
    .ZN(_08582_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17670 (.I(_05398_),
    .Z(net17670));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17454_ (.A1(net20827),
    .A2(_15578_[0]),
    .ZN(_08584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17455_ (.A1(_08584_),
    .A2(net20721),
    .ZN(_08585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17456_ (.I(_08585_),
    .ZN(_08586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17457_ (.A1(net20743),
    .A2(net20740),
    .ZN(_08587_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17668 (.I(_05398_),
    .Z(net17668));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17459_ (.A1(_08586_),
    .A2(net20515),
    .ZN(_08589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17460_ (.A1(net20745),
    .A2(net20823),
    .ZN(_08590_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17461_ (.I(_15575_[0]),
    .ZN(_08591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17462_ (.A1(_08591_),
    .A2(net20738),
    .ZN(_08592_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17463_ (.A1(net20513),
    .A2(net20334),
    .A3(net20589),
    .ZN(_08593_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17464_ (.A1(_08589_),
    .A2(_08593_),
    .A3(_07639_),
    .ZN(_08594_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _17465_ (.I(net20712),
    .ZN(_08595_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17660 (.I(_05551_),
    .Z(net17660));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17676 (.I(_05339_),
    .Z(net17676));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17468_ (.A1(_08582_),
    .A2(_08594_),
    .A3(_08595_),
    .ZN(_08598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17469_ (.A1(net20827),
    .A2(_08591_),
    .ZN(_08599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17470_ (.A1(_08599_),
    .A2(_07630_),
    .ZN(_08600_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17471_ (.I(_08600_),
    .ZN(_08601_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17472_ (.I(_15574_[0]),
    .ZN(_08602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17473_ (.A1(_08602_),
    .A2(net20740),
    .ZN(_08603_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17656 (.I(_05708_),
    .Z(net17656));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17475_ (.A1(_08601_),
    .A2(net20331),
    .ZN(_08605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17476_ (.A1(net20747),
    .A2(net20739),
    .ZN(_08606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17477_ (.A1(_08586_),
    .A2(_08606_),
    .ZN(_08607_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17478_ (.A1(_08605_),
    .A2(_08607_),
    .A3(_07639_),
    .ZN(_08608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17479_ (.A1(_08584_),
    .A2(net20587),
    .ZN(_08609_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17480_ (.I(_08609_),
    .ZN(_08610_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17481_ (.I(_15580_[0]),
    .ZN(_08611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17482_ (.A1(net20738),
    .A2(_08611_),
    .ZN(_08612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17483_ (.A1(_08610_),
    .A2(net20121),
    .ZN(_08613_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17663 (.I(_05482_),
    .Z(net17663));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17677 (.I(_05105_),
    .Z(net17677));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17486_ (.A1(_08590_),
    .A2(net20724),
    .Z(_08616_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17487_ (.I(_08616_),
    .ZN(_08617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17488_ (.A1(_08613_),
    .A2(net20855),
    .A3(_08617_),
    .ZN(_08618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17489_ (.A1(_08608_),
    .A2(_08618_),
    .A3(net20712),
    .ZN(_08619_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17490_ (.A1(_08598_),
    .A2(_08619_),
    .A3(net20710),
    .ZN(_08620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17491_ (.A1(net20738),
    .A2(net20821),
    .ZN(_08621_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17492_ (.A1(_08621_),
    .A2(net20721),
    .Z(_08622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17493_ (.A1(net20745),
    .A2(net20744),
    .ZN(_08623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17494_ (.A1(_08622_),
    .A2(_08623_),
    .ZN(_08624_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17495_ (.I(_08621_),
    .ZN(_08625_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17496_ (.A1(net20821),
    .A2(net20830),
    .ZN(_08626_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17708 (.I(_03881_),
    .Z(net17708));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17498_ (.A1(_08625_),
    .A2(_08626_),
    .B(net20585),
    .ZN(_08628_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17499_ (.A1(_08624_),
    .A2(_08628_),
    .A3(net20717),
    .ZN(_08629_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17500_ (.I(_15583_[0]),
    .ZN(_08630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17501_ (.A1(net20740),
    .A2(_08630_),
    .ZN(_08631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17502_ (.I(_08631_),
    .ZN(_08632_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17503_ (.I(_15587_[0]),
    .ZN(_08633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17504_ (.A1(net20823),
    .A2(_08633_),
    .ZN(_08634_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17505_ (.I(_08634_),
    .ZN(_08635_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17506_ (.A1(_08632_),
    .A2(_08635_),
    .B(net20586),
    .ZN(_08636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17507_ (.A1(net20823),
    .A2(net20622),
    .ZN(_08637_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17650 (.I(_06085_),
    .Z(net17650));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17509_ (.A1(net20330),
    .A2(_08637_),
    .A3(net20733),
    .ZN(_08639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17510_ (.A1(_08639_),
    .A2(net20851),
    .A3(_08636_),
    .ZN(_08640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17511_ (.A1(_08629_),
    .A2(_08640_),
    .A3(net20712),
    .ZN(_08641_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _17512_ (.I(net20708),
    .ZN(_08642_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17648 (.I(net17647),
    .Z(net17648));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17514_ (.A1(net20823),
    .A2(_08630_),
    .ZN(_08644_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17515_ (.I(_08644_),
    .ZN(_08645_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _17516_ (.A1(net20823),
    .A2(net20381),
    .ZN(_08646_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17517_ (.A1(_08645_),
    .A2(_08646_),
    .B(net20732),
    .ZN(_08647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17518_ (.A1(net20823),
    .A2(net20382),
    .ZN(_08648_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place17820 (.I(_00940_),
    .Z(net17820));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17520_ (.A1(net20330),
    .A2(_08648_),
    .A3(net20584),
    .ZN(_08650_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17822 (.I(net17820),
    .Z(net17822));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17522_ (.A1(_08647_),
    .A2(_08650_),
    .A3(net20851),
    .ZN(_08652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17523_ (.A1(net20826),
    .A2(net20830),
    .ZN(_08653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17524_ (.A1(net20740),
    .A2(net20621),
    .ZN(_08654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17525_ (.A1(_08653_),
    .A2(_08654_),
    .ZN(_08655_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17649 (.I(_06085_),
    .Z(net17649));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17821 (.I(net17820),
    .Z(net17821));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17528_ (.A1(_08655_),
    .A2(net20733),
    .ZN(_08658_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17643 (.I(_06177_),
    .Z(net17643));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17530_ (.A1(_08602_),
    .A2(net20823),
    .ZN(_08660_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17531_ (.I(_08660_),
    .ZN(_08661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17532_ (.A1(_08661_),
    .A2(net20586),
    .ZN(_08662_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17533_ (.A1(_08658_),
    .A2(net20717),
    .A3(net19906),
    .ZN(_08663_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17642 (.I(_06198_),
    .Z(net17642));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17535_ (.A1(_08652_),
    .A2(_08663_),
    .A3(_08595_),
    .ZN(_08665_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17536_ (.A1(_08665_),
    .A2(_08642_),
    .A3(_08641_),
    .ZN(_08666_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _17537_ (.I(net20847),
    .ZN(_08667_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17671 (.I(_05374_),
    .Z(net17671));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17539_ (.A1(_08620_),
    .A2(_08666_),
    .A3(_08667_),
    .ZN(_08669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17540_ (.A1(_08569_),
    .A2(_07630_),
    .ZN(_08670_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place17819 (.I(_00940_),
    .Z(net17819));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17542_ (.A1(_08645_),
    .A2(net20728),
    .ZN(_08672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17543_ (.A1(_08670_),
    .A2(_08672_),
    .Z(_08673_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17544_ (.I(_15578_[0]),
    .ZN(_08674_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17545_ (.A1(net20739),
    .A2(_08674_),
    .Z(_08675_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17546_ (.A1(_08675_),
    .A2(net20734),
    .B(net20848),
    .ZN(_08676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17547_ (.A1(_08673_),
    .A2(_08676_),
    .B(net20708),
    .ZN(_08677_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17548_ (.I(_15585_[0]),
    .ZN(_08678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17549_ (.A1(net20827),
    .A2(_08678_),
    .ZN(_08679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17550_ (.A1(_08679_),
    .A2(_07630_),
    .ZN(_08680_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17551_ (.I(_08680_),
    .ZN(_08681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17552_ (.A1(net20738),
    .A2(_15578_[0]),
    .ZN(_08682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17553_ (.A1(net19444),
    .A2(net20323),
    .ZN(_08683_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17554_ (.A1(_08683_),
    .A2(net20848),
    .A3(net20126),
    .ZN(_08684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17555_ (.A1(_08677_),
    .A2(_08684_),
    .B(_08595_),
    .ZN(_08685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17556_ (.A1(net20740),
    .A2(net20829),
    .ZN(_08686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17557_ (.A1(_08686_),
    .A2(net20721),
    .Z(_08687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17558_ (.A1(net20620),
    .A2(net20823),
    .ZN(_08688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17559_ (.A1(_08687_),
    .A2(net20504),
    .ZN(_08689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17560_ (.A1(net20825),
    .A2(net20384),
    .ZN(_08690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17561_ (.A1(net20512),
    .A2(_08690_),
    .A3(_07630_),
    .ZN(_08691_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17562_ (.A1(_08689_),
    .A2(_08691_),
    .B(_07639_),
    .ZN(_08692_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17653 (.I(_06080_),
    .Z(net17653));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17564_ (.A1(net20338),
    .A2(_08635_),
    .B(net20737),
    .ZN(_08694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17565_ (.A1(_08612_),
    .A2(net20580),
    .ZN(_08695_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17644 (.I(_06176_),
    .Z(net17644));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17567_ (.A1(_08694_),
    .A2(_08695_),
    .B(net20848),
    .ZN(_08697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17637 (.I(net17636),
    .Z(net17637));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17569_ (.A1(_08692_),
    .A2(_08697_),
    .B(net20708),
    .ZN(_08699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17570_ (.A1(_08685_),
    .A2(_08699_),
    .ZN(_08700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17571_ (.A1(net20827),
    .A2(_15580_[0]),
    .ZN(_08701_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17572_ (.I(_08701_),
    .ZN(_08702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17573_ (.A1(_08702_),
    .A2(net20723),
    .ZN(_08703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17574_ (.A1(_08581_),
    .A2(net20854),
    .A3(_08703_),
    .ZN(_08704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17575_ (.A1(net20738),
    .A2(net20383),
    .ZN(_08705_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17576_ (.I(_08705_),
    .ZN(_08706_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17577_ (.A1(net20113),
    .A2(_08702_),
    .B(net20721),
    .ZN(_08707_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17635 (.I(_06380_),
    .Z(net17635));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17579_ (.A1(net20589),
    .A2(_08603_),
    .ZN(_08709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17580_ (.A1(_08707_),
    .A2(_07639_),
    .A3(net20111),
    .ZN(_08710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17581_ (.A1(_08704_),
    .A2(_08710_),
    .A3(net20710),
    .ZN(_08711_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17582_ (.A1(_08576_),
    .A2(_08646_),
    .B(net20583),
    .ZN(_08712_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17583_ (.A1(net20666),
    .A2(net20323),
    .A3(net20728),
    .ZN(_08713_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17584_ (.A1(_08712_),
    .A2(_08713_),
    .A3(net20850),
    .ZN(_08714_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17585_ (.A1(net20578),
    .A2(_15599_[0]),
    .ZN(_08715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17586_ (.A1(_08715_),
    .A2(_07639_),
    .ZN(_08716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17587_ (.I(_08716_),
    .ZN(_08717_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17588_ (.I(net20504),
    .ZN(_08718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17589_ (.A1(_08718_),
    .A2(net20721),
    .ZN(_08719_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17590_ (.A1(_08717_),
    .A2(_08719_),
    .B(net20708),
    .ZN(_08720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17591_ (.A1(_08714_),
    .A2(_08720_),
    .ZN(_08721_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17592_ (.A1(_08711_),
    .A2(_08595_),
    .A3(_08721_),
    .ZN(_08722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17593_ (.A1(_08700_),
    .A2(_08722_),
    .A3(net20847),
    .ZN(_08723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17594_ (.A1(_08669_),
    .A2(_08723_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17595_ (.A1(net20722),
    .A2(_15592_[0]),
    .B(_07639_),
    .ZN(_08724_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17596_ (.I(_08724_),
    .ZN(_08725_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17597_ (.A1(_08611_),
    .A2(net20856),
    .A3(net21116),
    .ZN(_08726_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17598_ (.A1(net20321),
    .A2(net20110),
    .ZN(_08727_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17658 (.I(_05620_),
    .Z(net17658));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17600_ (.A1(_08725_),
    .A2(_08727_),
    .B(net20712),
    .ZN(_08729_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17601_ (.A1(net20334),
    .A2(net20325),
    .A3(net20582),
    .ZN(_08730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17602_ (.A1(net20323),
    .A2(net20110),
    .A3(net20725),
    .ZN(_08731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17603_ (.A1(_08730_),
    .A2(_08731_),
    .A3(net20850),
    .ZN(_08732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17604_ (.A1(_08729_),
    .A2(_08732_),
    .B(net20710),
    .ZN(_08733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17605_ (.A1(_08612_),
    .A2(net20721),
    .Z(_08734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17606_ (.A1(net19904),
    .A2(net20666),
    .ZN(_08735_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17607_ (.I(_08709_),
    .ZN(_08736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17608_ (.A1(_08736_),
    .A2(net20513),
    .ZN(_08737_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17609_ (.A1(_08735_),
    .A2(_08737_),
    .A3(net20714),
    .ZN(_08738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17610_ (.A1(_08687_),
    .A2(_08623_),
    .ZN(_08739_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17611_ (.A1(net20579),
    .A2(net20823),
    .Z(_08740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17612_ (.A1(_08740_),
    .A2(net20324),
    .ZN(_08741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17613_ (.A1(net20109),
    .A2(net20848),
    .A3(_08741_),
    .ZN(_08742_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17614_ (.A1(_08738_),
    .A2(_08742_),
    .A3(net20712),
    .ZN(_08743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17615_ (.A1(_08743_),
    .A2(_08733_),
    .ZN(_08744_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17616_ (.A1(net20747),
    .A2(net20830),
    .B(net20513),
    .C(net20578),
    .ZN(_08745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17617_ (.A1(_08606_),
    .A2(net20721),
    .Z(_08746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17618_ (.A1(_08746_),
    .A2(net20505),
    .ZN(_08747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17619_ (.A1(_08745_),
    .A2(net20853),
    .A3(_08747_),
    .ZN(_08748_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17620_ (.A1(_08576_),
    .A2(net20726),
    .B(net20848),
    .ZN(_08749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17621_ (.A1(_08726_),
    .A2(net20587),
    .ZN(_08750_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17622_ (.I(_08750_),
    .ZN(_08751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17623_ (.A1(net19443),
    .A2(net20507),
    .ZN(_08752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17624_ (.A1(_08646_),
    .A2(net20729),
    .ZN(_08753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17625_ (.A1(_08749_),
    .A2(_08752_),
    .A3(net20108),
    .ZN(_08754_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17626_ (.A1(_08748_),
    .A2(_08754_),
    .A3(_08595_),
    .ZN(_08755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17627_ (.A1(net20738),
    .A2(net20385),
    .Z(_08756_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17627 (.I(_06838_),
    .Z(net17627));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17629_ (.A1(_08756_),
    .A2(net20721),
    .B(net20714),
    .ZN(_08758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17630_ (.A1(_08637_),
    .A2(net20579),
    .ZN(_08759_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17631_ (.I(_08759_),
    .ZN(_08760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17632_ (.A1(_08760_),
    .A2(net20507),
    .ZN(_08761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17633_ (.A1(_08758_),
    .A2(_08761_),
    .B(_08595_),
    .ZN(_08762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17634_ (.A1(_08601_),
    .A2(_08587_),
    .ZN(_08763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17635_ (.A1(net20721),
    .A2(_08579_),
    .ZN(_08764_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17636_ (.A1(net19442),
    .A2(net20714),
    .A3(net19903),
    .ZN(_08765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17637_ (.A1(_08762_),
    .A2(_08765_),
    .B(_08642_),
    .ZN(_08766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17638_ (.A1(_08755_),
    .A2(_08766_),
    .ZN(_08767_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17639_ (.A1(_08744_),
    .A2(_08767_),
    .A3(net20847),
    .ZN(_08768_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17640_ (.A1(_08695_),
    .A2(net20339),
    .Z(_08769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17641_ (.A1(_08622_),
    .A2(net20664),
    .ZN(_08770_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17642_ (.A1(_08769_),
    .A2(_08770_),
    .A3(_08595_),
    .ZN(_08771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17643_ (.A1(_08746_),
    .A2(_08648_),
    .ZN(_08772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17644_ (.A1(net20125),
    .A2(net20581),
    .B(_08595_),
    .ZN(_08773_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17645_ (.A1(_08772_),
    .A2(_08773_),
    .A3(_08741_),
    .ZN(_08774_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17646_ (.A1(_08771_),
    .A2(_08774_),
    .A3(net20716),
    .ZN(_08775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17647_ (.A1(_08578_),
    .A2(_08644_),
    .B(net20584),
    .ZN(_08776_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17648_ (.I(_08776_),
    .ZN(_08777_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17649_ (.A1(net20712),
    .A2(_15601_[0]),
    .A3(net20726),
    .Z(_08778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17650_ (.A1(_08777_),
    .A2(_08778_),
    .ZN(_08779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17651_ (.A1(_08779_),
    .A2(net20848),
    .B(net20711),
    .ZN(_08780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17652_ (.A1(_08775_),
    .A2(_08780_),
    .B(net20847),
    .ZN(_08781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17653_ (.A1(_08646_),
    .A2(net20592),
    .ZN(_08782_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17654_ (.A1(net20721),
    .A2(_08688_),
    .ZN(_08783_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17655_ (.I(_08783_),
    .ZN(_08784_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _17656_ (.A1(net20126),
    .A2(_08749_),
    .A3(_08782_),
    .A4(_08784_),
    .ZN(_08785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17657_ (.A1(net20329),
    .A2(_08648_),
    .ZN(_08786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17658_ (.A1(_08769_),
    .A2(_08786_),
    .A3(net20848),
    .ZN(_08787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17659_ (.A1(_08785_),
    .A2(net20712),
    .A3(_08787_),
    .ZN(_08788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17660_ (.A1(_08764_),
    .A2(net20853),
    .ZN(_08789_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17661_ (.I(_08789_),
    .ZN(_08790_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17662_ (.A1(_08709_),
    .A2(net20666),
    .Z(_08791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17663_ (.A1(_08791_),
    .A2(_08790_),
    .B(net20712),
    .ZN(_08792_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17664_ (.I(_15589_[0]),
    .ZN(_08793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17665_ (.A1(net20825),
    .A2(_08793_),
    .ZN(_08794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17666_ (.A1(_08794_),
    .A2(net20721),
    .ZN(_08795_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _17667_ (.I(_08795_),
    .ZN(_08796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17668_ (.A1(_08796_),
    .A2(net20335),
    .ZN(_08797_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17669_ (.A1(_08761_),
    .A2(_08797_),
    .A3(net20714),
    .ZN(_08798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17670_ (.A1(_08792_),
    .A2(_08798_),
    .B(_08642_),
    .ZN(_08799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17671_ (.A1(_08799_),
    .A2(_08788_),
    .ZN(_08800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17672_ (.A1(_08781_),
    .A2(_08800_),
    .ZN(_08801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17673_ (.A1(_08768_),
    .A2(_08801_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17674_ (.A1(net20827),
    .A2(net20619),
    .ZN(_08802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17675_ (.A1(_08622_),
    .A2(_08802_),
    .ZN(_08803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17676_ (.A1(net20519),
    .A2(net20320),
    .A3(net20584),
    .ZN(_08804_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17677_ (.A1(_08803_),
    .A2(_08804_),
    .A3(net20718),
    .ZN(_08805_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17678_ (.A1(_08606_),
    .A2(net20114),
    .A3(net20727),
    .ZN(_08806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17679_ (.A1(_08603_),
    .A2(net20504),
    .A3(net20588),
    .ZN(_08807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17680_ (.A1(_08806_),
    .A2(_08807_),
    .ZN(_08808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17681_ (.A1(_08808_),
    .A2(net20848),
    .ZN(_08809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17682_ (.A1(_08805_),
    .A2(_08809_),
    .ZN(_08810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17683_ (.A1(_08810_),
    .A2(net20712),
    .ZN(_08811_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17684_ (.A1(_08751_),
    .A2(net20515),
    .ZN(_08812_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17685_ (.A1(_08707_),
    .A2(_08812_),
    .A3(net20854),
    .ZN(_08813_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17686_ (.I(_08802_),
    .ZN(_08814_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17687_ (.A1(_08814_),
    .A2(net20727),
    .B(net20848),
    .ZN(_08815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17688_ (.A1(_08751_),
    .A2(_08606_),
    .ZN(_08816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17689_ (.A1(_08706_),
    .A2(net20726),
    .ZN(_08817_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17690_ (.A1(_08815_),
    .A2(_08816_),
    .A3(_08817_),
    .ZN(_08818_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17691_ (.A1(_08813_),
    .A2(_08818_),
    .A3(_08595_),
    .ZN(_08819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17692_ (.A1(_08811_),
    .A2(_08819_),
    .A3(net20709),
    .ZN(_08820_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17693_ (.I(_08689_),
    .ZN(_08821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17694_ (.A1(_08701_),
    .A2(net20579),
    .ZN(_08822_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17695_ (.A1(_08822_),
    .A2(_08675_),
    .B(net20848),
    .ZN(_08823_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17696_ (.A1(_08821_),
    .A2(_08823_),
    .ZN(_08824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17697_ (.A1(net20506),
    .A2(net20336),
    .A3(net20582),
    .ZN(_08825_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17698_ (.A1(net20122),
    .A2(net20332),
    .A3(net20725),
    .ZN(_08826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17699_ (.A1(_08825_),
    .A2(_08826_),
    .B(net20850),
    .ZN(_08827_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17700_ (.A1(_08824_),
    .A2(_08827_),
    .B(_08595_),
    .ZN(_08828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17701_ (.A1(net20124),
    .A2(net20848),
    .Z(_08829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17702_ (.A1(_08760_),
    .A2(net20334),
    .ZN(_08830_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17703_ (.A1(_08829_),
    .A2(_08830_),
    .B(_08595_),
    .ZN(_08831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17704_ (.A1(net20825),
    .A2(net20380),
    .ZN(_08832_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17705_ (.I(_08832_),
    .ZN(_08833_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17706_ (.A1(net20327),
    .A2(_08833_),
    .B(net20586),
    .ZN(_08834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17707_ (.A1(net20664),
    .A2(_08603_),
    .A3(net20732),
    .ZN(_08835_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17708_ (.A1(_08834_),
    .A2(net20717),
    .A3(_08835_),
    .ZN(_08836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17709_ (.A1(_08831_),
    .A2(_08836_),
    .ZN(_08837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17710_ (.A1(_08828_),
    .A2(_08642_),
    .A3(_08837_),
    .ZN(_08838_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17711_ (.A1(_08820_),
    .A2(_08838_),
    .A3(_08667_),
    .ZN(_08839_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17712_ (.A1(_08623_),
    .A2(net20506),
    .A3(net20590),
    .ZN(_08840_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17713_ (.A1(net20379),
    .A2(net20590),
    .B(_08840_),
    .C(net20848),
    .ZN(_08841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17714_ (.A1(_08784_),
    .A2(_07639_),
    .Z(_08842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17715_ (.A1(_08632_),
    .A2(net20586),
    .ZN(_08843_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17716_ (.A1(net20516),
    .A2(_08648_),
    .A3(net20737),
    .ZN(_08844_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17717_ (.A1(_08842_),
    .A2(_08843_),
    .A3(_08844_),
    .ZN(_08845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17718_ (.A1(_08841_),
    .A2(_08595_),
    .A3(_08845_),
    .ZN(_08846_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17719_ (.A1(net20327),
    .A2(net20618),
    .B(net20586),
    .ZN(_08847_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17720_ (.A1(_08689_),
    .A2(_08847_),
    .A3(net20717),
    .ZN(_08848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17721_ (.A1(_08682_),
    .A2(net20583),
    .ZN(_08849_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17722_ (.A1(net20721),
    .A2(_15599_[0]),
    .Z(_08850_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17723_ (.I(_08850_),
    .ZN(_08851_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17724_ (.A1(net20107),
    .A2(net20115),
    .B(_08851_),
    .C(net20849),
    .ZN(_08852_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17725_ (.A1(_08848_),
    .A2(net20712),
    .A3(_08852_),
    .ZN(_08853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17726_ (.A1(_08846_),
    .A2(_08853_),
    .A3(net20708),
    .ZN(_08854_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17727_ (.A1(net20721),
    .A2(_15597_[0]),
    .Z(_08855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17728_ (.A1(_08829_),
    .A2(_08855_),
    .B(net20713),
    .ZN(_08856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17729_ (.A1(net20730),
    .A2(net20618),
    .ZN(_08857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17730_ (.A1(_08825_),
    .A2(net20716),
    .A3(_08857_),
    .ZN(_08858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17731_ (.A1(_08856_),
    .A2(_08858_),
    .B(net20709),
    .ZN(_08859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17732_ (.A1(_08760_),
    .A2(net20510),
    .ZN(_08860_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17733_ (.A1(_08777_),
    .A2(_08860_),
    .A3(net20715),
    .ZN(_08861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17734_ (.A1(_08736_),
    .A2(net20110),
    .ZN(_08862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17735_ (.A1(_08862_),
    .A2(net20850),
    .A3(_08753_),
    .ZN(_08863_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17736_ (.A1(_08861_),
    .A2(_08863_),
    .A3(net20713),
    .ZN(_08864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17737_ (.A1(_08859_),
    .A2(_08864_),
    .B(_08667_),
    .ZN(_08865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17738_ (.A1(_08854_),
    .A2(_08865_),
    .ZN(_08866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17739_ (.A1(_08839_),
    .A2(_08866_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17740_ (.A1(_08576_),
    .A2(net20665),
    .B(net20727),
    .ZN(_08867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17741_ (.A1(_08655_),
    .A2(net20584),
    .ZN(_08868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17742_ (.A1(_08867_),
    .A2(_08868_),
    .A3(net20851),
    .ZN(_08869_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17743_ (.I(_15594_[0]),
    .ZN(_08870_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17744_ (.A1(net20511),
    .A2(_08870_),
    .A3(net20733),
    .ZN(_08871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17745_ (.A1(_08871_),
    .A2(_08662_),
    .ZN(_08872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17746_ (.A1(_08872_),
    .A2(net20717),
    .ZN(_08873_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17747_ (.A1(_08869_),
    .A2(_08873_),
    .A3(_08595_),
    .ZN(_08874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17748_ (.A1(net20666),
    .A2(net20119),
    .ZN(_08875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17749_ (.A1(_08875_),
    .A2(net20731),
    .ZN(_08876_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17628 (.I(_06833_),
    .Z(net17628));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17751_ (.A1(_08646_),
    .A2(net20585),
    .B(net20848),
    .ZN(_08878_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17752_ (.A1(_08876_),
    .A2(_08878_),
    .A3(net19906),
    .ZN(_08879_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17753_ (.A1(net20519),
    .A2(_08654_),
    .A3(net20732),
    .ZN(_08880_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17754_ (.A1(_08592_),
    .A2(net20110),
    .A3(_07630_),
    .ZN(_08881_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17755_ (.A1(_08880_),
    .A2(_08881_),
    .A3(net20848),
    .ZN(_08882_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17756_ (.A1(_08879_),
    .A2(_08882_),
    .A3(net20712),
    .ZN(_08883_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17757_ (.A1(_08874_),
    .A2(_08883_),
    .A3(_08642_),
    .ZN(_08884_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17758_ (.A1(_08609_),
    .A2(net20848),
    .Z(_08885_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17759_ (.A1(_08867_),
    .A2(_08885_),
    .B(net20712),
    .ZN(_08886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17760_ (.A1(_08679_),
    .A2(net20721),
    .ZN(_08887_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17761_ (.I(_08887_),
    .ZN(_08888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17762_ (.A1(_08888_),
    .A2(net20507),
    .ZN(_08889_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17763_ (.A1(_08763_),
    .A2(_08889_),
    .A3(net20715),
    .ZN(_08890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17764_ (.A1(_08886_),
    .A2(_08890_),
    .B(_08642_),
    .ZN(_08891_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17765_ (.A1(net20330),
    .A2(net20117),
    .A3(net20733),
    .ZN(_08892_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17766_ (.A1(_08628_),
    .A2(net20717),
    .A3(_08892_),
    .ZN(_08893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17767_ (.A1(net20827),
    .A2(_08674_),
    .ZN(_08894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17768_ (.A1(net20119),
    .A2(_08894_),
    .B(net20731),
    .ZN(_08895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17769_ (.A1(_08578_),
    .A2(net20504),
    .B(net20584),
    .ZN(_08896_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17770_ (.A1(_08895_),
    .A2(_08896_),
    .B(net20848),
    .ZN(_08897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17771_ (.A1(_08893_),
    .A2(_08897_),
    .ZN(_08898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17772_ (.A1(_08898_),
    .A2(net20712),
    .ZN(_08899_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17773_ (.A1(_08891_),
    .A2(_08899_),
    .ZN(_08900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17774_ (.A1(_08884_),
    .A2(_08900_),
    .B(_08667_),
    .ZN(_08901_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17775_ (.A1(_08670_),
    .A2(_07639_),
    .Z(_08902_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17776_ (.A1(net20823),
    .A2(net20621),
    .ZN(_08903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17777_ (.A1(_08903_),
    .A2(net20721),
    .Z(_08904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17778_ (.A1(_08904_),
    .A2(net20712),
    .ZN(_08905_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17779_ (.A1(_08902_),
    .A2(_08905_),
    .Z(_08906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17780_ (.A1(_08587_),
    .A2(net20116),
    .B(net20586),
    .ZN(_08907_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17781_ (.I(_08662_),
    .ZN(_08908_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17782_ (.A1(_08907_),
    .A2(_08908_),
    .B(_08595_),
    .ZN(_08909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17783_ (.A1(_08906_),
    .A2(_08909_),
    .ZN(_08910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17784_ (.A1(_08910_),
    .A2(_08642_),
    .ZN(_08911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17785_ (.A1(_08601_),
    .A2(net20510),
    .ZN(_08912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17786_ (.A1(_08590_),
    .A2(_08603_),
    .A3(net20727),
    .ZN(_08913_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17787_ (.A1(_08912_),
    .A2(_08913_),
    .A3(_08595_),
    .ZN(_08914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17788_ (.A1(_08706_),
    .A2(net20583),
    .ZN(_08915_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17789_ (.A1(_08806_),
    .A2(net20712),
    .A3(_08915_),
    .ZN(_08916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17790_ (.A1(_08914_),
    .A2(_08916_),
    .B(net20718),
    .ZN(_08917_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17791_ (.A1(_08911_),
    .A2(_08917_),
    .B(_08667_),
    .ZN(_08918_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17792_ (.A1(_08680_),
    .A2(_08625_),
    .ZN(_08919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17793_ (.A1(_08919_),
    .A2(_08776_),
    .B(net20848),
    .ZN(_08920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17794_ (.A1(_08803_),
    .A2(net20718),
    .ZN(_08921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17795_ (.A1(_08920_),
    .A2(_08921_),
    .ZN(_08922_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17796_ (.A1(_08922_),
    .A2(_08595_),
    .ZN(_08923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17797_ (.A1(_08739_),
    .A2(_08712_),
    .A3(net20848),
    .ZN(_08924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17798_ (.A1(_08590_),
    .A2(_08705_),
    .ZN(_08925_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17799_ (.A1(_08925_),
    .A2(net20588),
    .ZN(_08926_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17800_ (.A1(_08603_),
    .A2(net20332),
    .A3(net20727),
    .ZN(_08927_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17801_ (.A1(_08926_),
    .A2(_08927_),
    .A3(net20718),
    .ZN(_08928_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17802_ (.A1(_08924_),
    .A2(net20712),
    .A3(_08928_),
    .ZN(_08929_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17803_ (.A1(_08923_),
    .A2(_08929_),
    .B(_08642_),
    .ZN(_08930_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17804_ (.A1(_08918_),
    .A2(_08930_),
    .ZN(_08931_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17805_ (.A1(_08901_),
    .A2(_08931_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17806_ (.A1(net20120),
    .A2(_08694_),
    .A3(net20848),
    .ZN(_08932_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17807_ (.I(_08919_),
    .ZN(_08933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17808_ (.A1(net20821),
    .A2(net20830),
    .ZN(_08934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17809_ (.A1(_08587_),
    .A2(_08934_),
    .ZN(_08935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17810_ (.A1(_08935_),
    .A2(net20736),
    .ZN(_08936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17811_ (.A1(_08933_),
    .A2(_08936_),
    .A3(net20720),
    .ZN(_08937_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17812_ (.A1(_08932_),
    .A2(_08937_),
    .A3(_08595_),
    .ZN(_08938_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17813_ (.A1(net20721),
    .A2(net20622),
    .Z(_08939_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17814_ (.A1(_08939_),
    .A2(net20319),
    .B(net20848),
    .ZN(_08940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17815_ (.A1(_08940_),
    .A2(net20712),
    .ZN(_08941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17816_ (.A1(_08681_),
    .A2(_08587_),
    .ZN(_08942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17817_ (.A1(_08676_),
    .A2(_08942_),
    .Z(_08943_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17818_ (.A1(_08943_),
    .A2(_08941_),
    .Z(_08944_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17819_ (.A1(_08944_),
    .A2(net20508),
    .A3(_08938_),
    .ZN(_08945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17820_ (.A1(net20329),
    .A2(net20333),
    .ZN(_08946_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17821_ (.A1(_08740_),
    .A2(net20719),
    .ZN(_08947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17822_ (.A1(_08946_),
    .A2(_08947_),
    .B(net20712),
    .ZN(_08948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17823_ (.A1(_08753_),
    .A2(_07639_),
    .Z(_08949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17824_ (.A1(_08949_),
    .A2(_08769_),
    .A3(net20127),
    .ZN(_08950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17825_ (.A1(_08948_),
    .A2(_08950_),
    .ZN(_08951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17826_ (.A1(_08734_),
    .A2(net20505),
    .ZN(_08952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17827_ (.A1(_08581_),
    .A2(_08952_),
    .A3(net20853),
    .ZN(_08953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17828_ (.A1(_08759_),
    .A2(net20719),
    .Z(_08954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17829_ (.A1(_08954_),
    .A2(net19902),
    .B(_08595_),
    .ZN(_08955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17830_ (.A1(_08953_),
    .A2(_08955_),
    .ZN(_08956_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17831_ (.A1(_08951_),
    .A2(_08956_),
    .A3(net20711),
    .ZN(_08957_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17832_ (.A1(_08667_),
    .A2(_08957_),
    .A3(_08945_),
    .ZN(_08958_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17833_ (.A1(net20340),
    .A2(net20107),
    .B(_08826_),
    .C(net20716),
    .ZN(_08959_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17834_ (.A1(_08782_),
    .A2(net20848),
    .Z(_08960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17835_ (.A1(_08740_),
    .A2(net20828),
    .ZN(_08961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17836_ (.A1(_08960_),
    .A2(_08731_),
    .A3(_08961_),
    .ZN(_08962_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17837_ (.A1(_08959_),
    .A2(_08595_),
    .A3(_08962_),
    .ZN(_08963_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17838_ (.A1(_08701_),
    .A2(net20578),
    .B(_07639_),
    .ZN(_08964_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17839_ (.I(_08964_),
    .ZN(_08965_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17840_ (.A1(net20319),
    .A2(net20112),
    .ZN(_08966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17841_ (.A1(_08965_),
    .A2(_08966_),
    .B(_08595_),
    .ZN(_08967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17842_ (.A1(_08592_),
    .A2(net20729),
    .ZN(_08968_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17843_ (.A1(_08968_),
    .A2(_08661_),
    .Z(_08969_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17844_ (.A1(net20848),
    .A2(_08683_),
    .A3(_08969_),
    .ZN(_08970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17845_ (.A1(_08967_),
    .A2(_08970_),
    .B(net20711),
    .ZN(_08971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17846_ (.A1(_08971_),
    .A2(_08963_),
    .ZN(_08972_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17847_ (.A1(net20506),
    .A2(net20118),
    .A3(net20591),
    .ZN(_08973_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17848_ (.A1(_08936_),
    .A2(net20720),
    .A3(_08973_),
    .Z(_08974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17849_ (.A1(_08770_),
    .A2(_08840_),
    .B(net20720),
    .ZN(_08975_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17850_ (.A1(_08974_),
    .A2(_08975_),
    .B(_08595_),
    .ZN(_08976_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17851_ (.A1(net20327),
    .A2(net20378),
    .B(net20590),
    .ZN(_08977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17852_ (.A1(_08772_),
    .A2(_08977_),
    .A3(net20852),
    .ZN(_08978_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17853_ (.A1(net20338),
    .A2(net20852),
    .ZN(_08979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17854_ (.A1(_08979_),
    .A2(net19905),
    .B(_08595_),
    .ZN(_08980_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17855_ (.A1(_08978_),
    .A2(_08980_),
    .B(_08642_),
    .ZN(_08981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17856_ (.A1(_08976_),
    .A2(_08981_),
    .ZN(_08982_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17857_ (.A1(_08972_),
    .A2(_08982_),
    .A3(net20847),
    .ZN(_08983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17858_ (.A1(_08983_),
    .A2(_08958_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17859_ (.A1(_08965_),
    .A2(net20123),
    .B(net20709),
    .ZN(_08984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17860_ (.A1(net20510),
    .A2(net20580),
    .ZN(_08985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17861_ (.A1(_08985_),
    .A2(net20106),
    .ZN(_08986_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17862_ (.A1(_08789_),
    .A2(_08986_),
    .Z(_08987_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17863_ (.A1(_08984_),
    .A2(_08987_),
    .B(net20847),
    .ZN(_08988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17864_ (.A1(_08610_),
    .A2(net20331),
    .ZN(_08989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17865_ (.A1(_08888_),
    .A2(_08587_),
    .ZN(_08990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17866_ (.A1(_08989_),
    .A2(_08990_),
    .B(net20854),
    .ZN(_08991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17867_ (.A1(_07630_),
    .A2(net20821),
    .ZN(_08992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17868_ (.A1(_08624_),
    .A2(_08992_),
    .B(net20715),
    .ZN(_08993_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17869_ (.A1(_08991_),
    .A2(_08993_),
    .B(net20710),
    .ZN(_08994_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17870_ (.A1(_08988_),
    .A2(_08994_),
    .B(_08595_),
    .ZN(_08995_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17871_ (.A1(_08601_),
    .A2(net20121),
    .Z(_08996_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17872_ (.A1(_08996_),
    .A2(_08571_),
    .B(net20854),
    .ZN(_08997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17873_ (.A1(_08751_),
    .A2(net20510),
    .Z(_08998_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17874_ (.A1(_08682_),
    .A2(net20114),
    .A3(net20727),
    .Z(_08999_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17875_ (.A1(_08998_),
    .A2(_08999_),
    .B(net20715),
    .ZN(_09000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17876_ (.A1(_08997_),
    .A2(_09000_),
    .A3(net20709),
    .ZN(_09001_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17877_ (.A1(_08579_),
    .A2(_08645_),
    .A3(net20725),
    .Z(_09002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17878_ (.A1(_08616_),
    .A2(net20663),
    .ZN(_09003_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17879_ (.A1(_09002_),
    .A2(_09003_),
    .A3(net20715),
    .ZN(_09004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17880_ (.A1(net20725),
    .A2(net20821),
    .ZN(_09005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17881_ (.A1(_09005_),
    .A2(net20830),
    .ZN(_09006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17882_ (.A1(net20127),
    .A2(_09006_),
    .ZN(_09007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17883_ (.A1(_09007_),
    .A2(net20853),
    .ZN(_09008_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17884_ (.A1(_09004_),
    .A2(_08642_),
    .A3(_09008_),
    .ZN(_09009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17885_ (.A1(_09001_),
    .A2(_09009_),
    .ZN(_09010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17886_ (.A1(_09010_),
    .A2(net20847),
    .ZN(_09011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17887_ (.A1(_08995_),
    .A2(_09011_),
    .ZN(_09012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17888_ (.A1(_07639_),
    .A2(_08894_),
    .ZN(_09013_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17889_ (.A1(_08734_),
    .A2(_09013_),
    .Z(_09014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17890_ (.A1(_09014_),
    .A2(net20708),
    .Z(_09015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17891_ (.A1(_08603_),
    .A2(net20724),
    .ZN(_09016_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17892_ (.A1(_08926_),
    .A2(net20855),
    .A3(_09016_),
    .ZN(_09017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17893_ (.A1(_09015_),
    .A2(_09017_),
    .B(_08667_),
    .ZN(_09018_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17894_ (.A1(_08654_),
    .A2(net20586),
    .Z(_09019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17895_ (.A1(_09019_),
    .A2(_08648_),
    .ZN(_09020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17896_ (.A1(_08814_),
    .A2(net20728),
    .ZN(_09021_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17897_ (.A1(_09020_),
    .A2(net20849),
    .A3(_09021_),
    .ZN(_09022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17898_ (.A1(_08796_),
    .A2(net20506),
    .ZN(_09023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17899_ (.A1(_08842_),
    .A2(_09023_),
    .ZN(_09024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17900_ (.A1(_09022_),
    .A2(_09024_),
    .A3(_08642_),
    .ZN(_09025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17901_ (.A1(_09025_),
    .A2(_09018_),
    .B(net20712),
    .ZN(_09026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17902_ (.A1(_08746_),
    .A2(net20110),
    .ZN(_09027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17903_ (.A1(_09027_),
    .A2(_08581_),
    .A3(net20853),
    .ZN(_09028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17904_ (.A1(net19907),
    .A2(net20581),
    .ZN(_09029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17905_ (.A1(_08815_),
    .A2(net19903),
    .A3(_09029_),
    .ZN(_09030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17906_ (.A1(_09028_),
    .A2(net20711),
    .A3(_09030_),
    .ZN(_09031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17907_ (.A1(_08736_),
    .A2(_08690_),
    .ZN(_09032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17908_ (.I(net20318),
    .ZN(_09033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17909_ (.A1(_09032_),
    .A2(_08815_),
    .A3(_09033_),
    .ZN(_09034_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17910_ (.A1(net20824),
    .A2(net20518),
    .B(net20721),
    .ZN(_09035_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17911_ (.A1(net20384),
    .A2(net20735),
    .B(_09035_),
    .C(net20848),
    .ZN(_09036_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17912_ (.A1(_09034_),
    .A2(_09036_),
    .A3(_08642_),
    .ZN(_09037_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17913_ (.A1(_09031_),
    .A2(_09037_),
    .A3(_08667_),
    .ZN(_09038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17914_ (.A1(_09026_),
    .A2(_09038_),
    .ZN(_09039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17915_ (.A1(_09012_),
    .A2(_09039_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17916_ (.I(_08654_),
    .ZN(_09040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17917_ (.A1(_09040_),
    .A2(net20724),
    .ZN(_09041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17918_ (.A1(_08926_),
    .A2(net20855),
    .A3(_09041_),
    .ZN(_09042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17919_ (.A1(_08725_),
    .A2(_08607_),
    .ZN(_09043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17920_ (.A1(_09042_),
    .A2(_09043_),
    .ZN(_09044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17921_ (.A1(_09044_),
    .A2(_08595_),
    .ZN(_09045_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17922_ (.A1(_08576_),
    .A2(net20727),
    .A3(net20665),
    .Z(_09046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17923_ (.A1(net20514),
    .A2(_08894_),
    .A3(net20727),
    .ZN(_09047_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17924_ (.A1(_09046_),
    .A2(net20848),
    .A3(_09047_),
    .ZN(_09048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17925_ (.A1(_08623_),
    .A2(_07630_),
    .ZN(_09049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17926_ (.A1(_09049_),
    .A2(_08968_),
    .ZN(_09050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17927_ (.A1(_07639_),
    .A2(net20666),
    .Z(_09051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17928_ (.A1(_09050_),
    .A2(_09051_),
    .B(_08595_),
    .ZN(_09052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17929_ (.A1(_09048_),
    .A2(_09052_),
    .ZN(_09053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17930_ (.A1(_09045_),
    .A2(_09053_),
    .A3(net20710),
    .ZN(_09054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17931_ (.A1(_08690_),
    .A2(net20725),
    .ZN(_09055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17932_ (.A1(_08942_),
    .A2(_09055_),
    .ZN(_09056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17933_ (.A1(_09056_),
    .A2(net20715),
    .ZN(_09057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17934_ (.A1(_08823_),
    .A2(_08595_),
    .Z(_09058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17935_ (.A1(_09057_),
    .A2(_09058_),
    .B(net20709),
    .ZN(_09059_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17936_ (.A1(net20317),
    .A2(net20123),
    .B(_08749_),
    .ZN(_09060_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17937_ (.A1(net20722),
    .A2(_15593_[0]),
    .Z(_09061_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17938_ (.A1(_08990_),
    .A2(net20854),
    .A3(_09061_),
    .ZN(_09062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17939_ (.A1(_09060_),
    .A2(_09062_),
    .ZN(_09063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17940_ (.A1(_09063_),
    .A2(net20713),
    .ZN(_09064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17941_ (.A1(_09059_),
    .A2(_09064_),
    .ZN(_09065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17942_ (.A1(_09054_),
    .A2(_09065_),
    .ZN(_09066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17943_ (.A1(_09066_),
    .A2(_08667_),
    .ZN(_09067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17944_ (.A1(_08888_),
    .A2(_08592_),
    .ZN(_09068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17945_ (.A1(net20824),
    .A2(net20517),
    .ZN(_09069_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17946_ (.A1(_09069_),
    .A2(net20721),
    .ZN(_09070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17947_ (.I(_09070_),
    .ZN(_09071_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17948_ (.A1(_09068_),
    .A2(net20849),
    .A3(_08670_),
    .A4(_09071_),
    .Z(_09072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17949_ (.A1(net20328),
    .A2(net20504),
    .ZN(_09073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17950_ (.A1(_09073_),
    .A2(net20718),
    .A3(_08926_),
    .ZN(_09074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17951_ (.A1(_09074_),
    .A2(_08595_),
    .ZN(_09075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17952_ (.A1(_08833_),
    .A2(net20579),
    .ZN(_09076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17953_ (.A1(_08949_),
    .A2(_08915_),
    .A3(_09076_),
    .ZN(_09077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17954_ (.A1(_08935_),
    .A2(net20579),
    .ZN(_09078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17955_ (.A1(net20742),
    .A2(net20721),
    .ZN(_09079_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17956_ (.A1(_09079_),
    .A2(net20848),
    .Z(_09080_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17957_ (.A1(_09078_),
    .A2(_09080_),
    .B(_08595_),
    .ZN(_09081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17958_ (.A1(_09077_),
    .A2(_09081_),
    .ZN(_09082_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17959_ (.A1(_09072_),
    .A2(_09075_),
    .B(net20708),
    .C(_09082_),
    .ZN(_09083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17960_ (.A1(_08586_),
    .A2(net20331),
    .ZN(_09084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17961_ (.A1(_08855_),
    .A2(_07639_),
    .ZN(_09085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17962_ (.I(_09085_),
    .ZN(_09086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17963_ (.A1(_09084_),
    .A2(_09086_),
    .B(_08595_),
    .ZN(_09087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17964_ (.A1(_08610_),
    .A2(net20515),
    .ZN(_09088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17965_ (.A1(_08796_),
    .A2(net20507),
    .ZN(_09089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17966_ (.A1(_09088_),
    .A2(_09089_),
    .A3(net20855),
    .ZN(_09090_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17967_ (.A1(_09087_),
    .A2(_09090_),
    .B(net20710),
    .ZN(_09091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17968_ (.A1(_08672_),
    .A2(_07639_),
    .Z(_09092_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17969_ (.I(_08849_),
    .ZN(_09093_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17970_ (.A1(_09093_),
    .A2(net20664),
    .ZN(_09094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17971_ (.A1(_09092_),
    .A2(_09094_),
    .B(net20712),
    .ZN(_09095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17972_ (.A1(_09093_),
    .A2(net20666),
    .ZN(_09096_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17973_ (.A1(_09073_),
    .A2(_09096_),
    .A3(net20848),
    .ZN(_09097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17974_ (.A1(_09095_),
    .A2(_09097_),
    .ZN(_09098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17975_ (.A1(_09091_),
    .A2(_09098_),
    .B(_08667_),
    .ZN(_09099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17976_ (.A1(_09083_),
    .A2(_09099_),
    .ZN(_09100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17977_ (.A1(_09067_),
    .A2(_09100_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17978_ (.A1(_08637_),
    .A2(net20731),
    .ZN(_09101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17979_ (.A1(_08849_),
    .A2(_09101_),
    .ZN(_09102_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17980_ (.A1(_09102_),
    .A2(net20718),
    .A3(_09041_),
    .Z(_09103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17981_ (.A1(net20337),
    .A2(net20588),
    .ZN(_09104_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17982_ (.A1(_09016_),
    .A2(_09104_),
    .A3(net20848),
    .Z(_09105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17983_ (.A1(_09103_),
    .A2(_09105_),
    .B(_08595_),
    .ZN(_09106_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17984_ (.A1(_08985_),
    .A2(net20339),
    .B(net20716),
    .C(_09005_),
    .ZN(_09107_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17985_ (.A1(net20516),
    .A2(net20509),
    .A3(net20737),
    .ZN(_09108_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17986_ (.A1(_08840_),
    .A2(_09108_),
    .A3(net20852),
    .ZN(_09109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17987_ (.A1(_09107_),
    .A2(_09109_),
    .A3(net20712),
    .ZN(_09110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17988_ (.A1(_09106_),
    .A2(_08667_),
    .A3(_09110_),
    .ZN(_09111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17989_ (.I(_08817_),
    .ZN(_09112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17990_ (.A1(net20590),
    .A2(_15603_[0]),
    .ZN(_09113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17991_ (.A1(_09113_),
    .A2(net20848),
    .ZN(_09114_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17992_ (.A1(_09112_),
    .A2(_09114_),
    .ZN(_09115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17993_ (.A1(net20115),
    .A2(net20730),
    .ZN(_09116_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17994_ (.A1(_09115_),
    .A2(_09116_),
    .B(net20712),
    .ZN(_09117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17995_ (.A1(_09019_),
    .A2(net20325),
    .ZN(_09118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17996_ (.A1(_08749_),
    .A2(_09118_),
    .A3(_08851_),
    .ZN(_09119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17997_ (.A1(_09117_),
    .A2(_09119_),
    .ZN(_09120_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17998_ (.A1(_08832_),
    .A2(net20579),
    .B(net20848),
    .ZN(_09121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17999_ (.A1(net20579),
    .A2(net20517),
    .Z(_09122_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18000_ (.A1(_09121_),
    .A2(_09122_),
    .Z(_09123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18001_ (.A1(_09123_),
    .A2(net20712),
    .Z(_09124_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18002_ (.A1(_08769_),
    .A2(_08676_),
    .A3(net20127),
    .ZN(_09125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18003_ (.A1(_09124_),
    .A2(_09125_),
    .ZN(_09126_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18004_ (.A1(_09120_),
    .A2(_09126_),
    .A3(net20847),
    .ZN(_09127_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18005_ (.A1(_09111_),
    .A2(_09127_),
    .A3(net20508),
    .ZN(_09128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18006_ (.A1(net20322),
    .A2(_08637_),
    .ZN(_09129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18007_ (.A1(_08933_),
    .A2(_09129_),
    .A3(net20720),
    .ZN(_09130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18008_ (.A1(_09019_),
    .A2(_08690_),
    .ZN(_09131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18009_ (.A1(net20740),
    .A2(net20326),
    .ZN(_09132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18010_ (.A1(_09132_),
    .A2(net20316),
    .ZN(_09133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18011_ (.A1(_09133_),
    .A2(net20736),
    .ZN(_09134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18012_ (.A1(_09131_),
    .A2(net20852),
    .A3(_09134_),
    .ZN(_09135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18013_ (.A1(_09130_),
    .A2(_09135_),
    .A3(net20712),
    .ZN(_09136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18014_ (.A1(net20734),
    .A2(net20385),
    .ZN(_09137_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18015_ (.A1(_09078_),
    .A2(net20719),
    .A3(_09137_),
    .ZN(_09138_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18016_ (.A1(net20519),
    .A2(net20735),
    .B(_09132_),
    .ZN(_09139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18017_ (.A1(_09139_),
    .A2(_09121_),
    .Z(_09140_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18018_ (.A1(_09138_),
    .A2(_09140_),
    .A3(_08595_),
    .ZN(_09141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18019_ (.A1(_09136_),
    .A2(_09141_),
    .A3(net20847),
    .ZN(_09142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18020_ (.A1(_08968_),
    .A2(net20848),
    .Z(_09143_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18021_ (.A1(_09143_),
    .A2(_08942_),
    .B(_08595_),
    .ZN(_09144_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18022_ (.A1(_08616_),
    .A2(_09070_),
    .B(net20323),
    .ZN(_09145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18023_ (.A1(_09145_),
    .A2(_08878_),
    .ZN(_09146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18024_ (.A1(_09144_),
    .A2(_09146_),
    .B(net20847),
    .ZN(_09147_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18025_ (.A1(_08847_),
    .A2(_09068_),
    .A3(net20849),
    .ZN(_09148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18026_ (.A1(net20716),
    .A2(_08730_),
    .A3(_08913_),
    .ZN(_09149_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18027_ (.A1(_09148_),
    .A2(_08595_),
    .A3(_09149_),
    .ZN(_09150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18028_ (.A1(_09150_),
    .A2(_09147_),
    .ZN(_09151_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18029_ (.A1(_09142_),
    .A2(_09151_),
    .A3(net20711),
    .ZN(_09152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18030_ (.A1(_09152_),
    .A2(_09128_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18031_ (.A1(net21527),
    .A2(_07550_),
    .B(_07553_),
    .ZN(_15605_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18032_ (.A1(net20922),
    .A2(net21519),
    .B(_07561_),
    .ZN(_09153_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17626 (.I(_06876_),
    .Z(net17626));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17655 (.I(_05725_),
    .Z(net17655));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18035_ (.A1(_07541_),
    .A2(net21526),
    .B(_07545_),
    .ZN(_15606_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18036_ (.A1(net20775),
    .A2(net20814),
    .ZN(_09155_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18037_ (.I(_09155_),
    .ZN(_09156_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17659 (.I(_05571_),
    .Z(net17659));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17622 (.I(_06902_),
    .Z(net17622));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18040_ (.A1(_09156_),
    .A2(net20762),
    .ZN(_09159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18041_ (.I(_15608_[0]),
    .ZN(_09160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18042_ (.A1(_09160_),
    .A2(net20771),
    .ZN(_09161_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18043_ (.I(_09161_),
    .ZN(_09162_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17620 (.I(_06945_),
    .Z(net17620));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18045_ (.A1(_09162_),
    .A2(net20757),
    .ZN(_09164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18046_ (.A1(net20814),
    .A2(_09160_),
    .ZN(_09165_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17619 (.I(_06962_),
    .Z(net17619));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17618 (.I(_06984_),
    .Z(net17618));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18049_ (.A1(net20312),
    .A2(net20597),
    .ZN(_09168_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18050_ (.A1(net20105),
    .A2(_09164_),
    .A3(_09168_),
    .ZN(_09169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18051_ (.A1(_09169_),
    .A2(net20859),
    .ZN(_09170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18052_ (.I(_15621_[0]),
    .ZN(_09171_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18053_ (.A1(net20771),
    .A2(_09171_),
    .Z(_09172_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18054_ (.I(_15617_[0]),
    .ZN(_09173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18055_ (.A1(net20814),
    .A2(_09173_),
    .ZN(_09174_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18056_ (.I(_09174_),
    .ZN(_09175_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17617 (.I(_06996_),
    .Z(net17617));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18058_ (.A1(_09172_),
    .A2(_09175_),
    .B(net20766),
    .ZN(_09177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18059_ (.A1(_07571_),
    .A2(_09161_),
    .ZN(_09178_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18060_ (.I(_09178_),
    .ZN(_09179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18061_ (.A1(net20816),
    .A2(net20372),
    .ZN(_09180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18062_ (.A1(_09179_),
    .A2(_09180_),
    .ZN(_09181_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18063_ (.I(_07578_),
    .ZN(_09182_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17824 (.I(net17820),
    .Z(net17824));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17623 (.I(_06896_),
    .Z(net17623));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18066_ (.A1(_09177_),
    .A2(_09181_),
    .A3(net20654),
    .ZN(_09185_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _18067_ (.I(_07586_),
    .ZN(_09186_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17614 (.I(_07053_),
    .Z(net17614));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18069_ (.A1(_09170_),
    .A2(_09185_),
    .A3(net20499),
    .ZN(_09188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18070_ (.A1(net20771),
    .A2(_09173_),
    .ZN(_09189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18071_ (.I(_09189_),
    .ZN(_09190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18072_ (.A1(net20816),
    .A2(_09171_),
    .ZN(_09191_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18073_ (.I(_09191_),
    .ZN(_09192_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18074_ (.A1(_09190_),
    .A2(net19898),
    .B(net20597),
    .ZN(_09193_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18075_ (.A1(_09161_),
    .A2(net20763),
    .Z(_09194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18076_ (.A1(net20813),
    .A2(net20617),
    .ZN(_09195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18077_ (.A1(_09194_),
    .A2(net20491),
    .ZN(_09196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18078_ (.A1(_09193_),
    .A2(_09196_),
    .A3(net20656),
    .ZN(_09197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18079_ (.A1(net20771),
    .A2(net20812),
    .ZN(_09198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18080_ (.A1(_09198_),
    .A2(net20757),
    .ZN(_09199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _18081_ (.I(_09199_),
    .ZN(_09200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18082_ (.A1(net20776),
    .A2(net20773),
    .ZN(_09201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18083_ (.A1(_09200_),
    .A2(_09201_),
    .ZN(_09202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18084_ (.A1(net20813),
    .A2(net20811),
    .ZN(_09203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18085_ (.A1(net20776),
    .A2(net20819),
    .ZN(_09204_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17657 (.I(_05635_),
    .Z(net17657));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18087_ (.A1(_09203_),
    .A2(_09204_),
    .A3(net20597),
    .ZN(_09206_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17613 (.I(_07134_),
    .Z(net17613));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18089_ (.A1(_09202_),
    .A2(_09206_),
    .A3(net20861),
    .ZN(_09208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18090_ (.A1(_09197_),
    .A2(_09208_),
    .A3(net20754),
    .ZN(_09209_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _18091_ (.I(_00403_),
    .ZN(_09210_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17624 (.I(_06896_),
    .Z(net17624));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18093_ (.A1(_09188_),
    .A2(_09209_),
    .A3(_09210_),
    .ZN(_09212_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _18094_ (.I(_00404_),
    .ZN(_09213_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17610 (.I(_15739_[0]),
    .Z(net17610));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18096_ (.A1(net20776),
    .A2(net20813),
    .ZN(_09215_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18097_ (.A1(net20486),
    .A2(net20763),
    .Z(_09216_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17621 (.I(_06908_),
    .Z(net17621));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18099_ (.A1(_09216_),
    .A2(net20861),
    .ZN(_09218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18100_ (.A1(net20814),
    .A2(net20377),
    .ZN(_09219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18101_ (.A1(_09219_),
    .A2(net20594),
    .ZN(_09220_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18102_ (.I(_09220_),
    .ZN(_09221_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17611 (.I(_07294_),
    .Z(net17611));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18104_ (.I(_15614_[0]),
    .ZN(_09223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18105_ (.A1(net20767),
    .A2(_09223_),
    .ZN(_09224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18106_ (.A1(_09221_),
    .A2(net20100),
    .ZN(_09225_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17612 (.I(_07155_),
    .Z(net17612));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18108_ (.A1(_09218_),
    .A2(_09225_),
    .B(net20495),
    .ZN(_09227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18109_ (.A1(net20776),
    .A2(net20767),
    .B(net20594),
    .ZN(_09228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18110_ (.A1(_09228_),
    .A2(net20310),
    .ZN(_09229_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18111_ (.I(_15609_[0]),
    .ZN(_09230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18112_ (.A1(net20814),
    .A2(_09230_),
    .ZN(_09231_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18113_ (.A1(_09231_),
    .A2(net20594),
    .ZN(_09232_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18114_ (.I(_09232_),
    .ZN(_09233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18115_ (.A1(_09233_),
    .A2(net20314),
    .ZN(_09234_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18241 (.I(net18240),
    .Z(net18241));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18117_ (.A1(_09229_),
    .A2(_09234_),
    .A3(net20861),
    .ZN(_09236_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17606 (.I(_15753_[0]),
    .Z(net17606));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18119_ (.A1(_09227_),
    .A2(_09236_),
    .B(_09210_),
    .ZN(_09238_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18120_ (.A1(net20771),
    .A2(_15623_[0]),
    .Z(_09239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18121_ (.A1(_09239_),
    .A2(net20766),
    .ZN(_09240_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18122_ (.A1(_09159_),
    .A2(_09240_),
    .Z(_09241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18123_ (.A1(net20599),
    .A2(net20811),
    .Z(_09242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18124_ (.A1(_09242_),
    .A2(net20813),
    .ZN(_09243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18125_ (.I(_15607_[0]),
    .ZN(_09244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18126_ (.A1(net20770),
    .A2(_09244_),
    .ZN(_09245_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18127_ (.I(_09245_),
    .ZN(_09246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18128_ (.A1(_09246_),
    .A2(net20594),
    .B(net20859),
    .ZN(_09247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18129_ (.A1(_09241_),
    .A2(_09243_),
    .A3(_09247_),
    .ZN(_09248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18130_ (.A1(net20775),
    .A2(net20771),
    .ZN(_09249_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18131_ (.A1(_09249_),
    .A2(net20760),
    .Z(_09250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18132_ (.A1(_09250_),
    .A2(net20310),
    .ZN(_09251_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18242 (.I(net18240),
    .Z(net18242));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18134_ (.A1(net20487),
    .A2(net20594),
    .Z(_09253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18135_ (.A1(net20769),
    .A2(_09230_),
    .ZN(_09254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18136_ (.A1(_09253_),
    .A2(net20303),
    .ZN(_09255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18137_ (.A1(_09251_),
    .A2(_09255_),
    .A3(net20861),
    .ZN(_09256_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17605 (.I(_15867_[0]),
    .Z(net17605));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18139_ (.A1(_09248_),
    .A2(_09256_),
    .A3(net20496),
    .ZN(_09258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18140_ (.A1(_09238_),
    .A2(_09258_),
    .ZN(_09259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18141_ (.A1(_09212_),
    .A2(_09213_),
    .A3(_09259_),
    .ZN(_09260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18142_ (.A1(net20813),
    .A2(net20375),
    .ZN(_09261_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18143_ (.A1(_09261_),
    .A2(_07571_),
    .Z(_09262_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18144_ (.A1(_09247_),
    .A2(_09243_),
    .A3(_09262_),
    .ZN(_09263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18145_ (.A1(_09262_),
    .A2(net20859),
    .Z(_09264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18146_ (.A1(net20771),
    .A2(net20373),
    .ZN(_09265_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18147_ (.I(_09265_),
    .ZN(_09266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18148_ (.A1(_09266_),
    .A2(net20763),
    .ZN(_09267_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18149_ (.A1(_09267_),
    .A2(net20101),
    .Z(_09268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18150_ (.A1(_09264_),
    .A2(_09268_),
    .ZN(_09269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18151_ (.A1(_09263_),
    .A2(_09269_),
    .A3(_09186_),
    .ZN(_09270_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17604 (.I(_15868_[0]),
    .Z(net17604));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18153_ (.A1(net20305),
    .A2(_09192_),
    .B(net20766),
    .ZN(_09272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18154_ (.A1(_09224_),
    .A2(net20596),
    .ZN(_09273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18155_ (.A1(_09272_),
    .A2(net20859),
    .A3(net19897),
    .ZN(_09274_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18156_ (.A1(net20776),
    .A2(net20767),
    .ZN(_09275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18157_ (.A1(net20815),
    .A2(net20374),
    .ZN(_09276_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18158_ (.A1(net20482),
    .A2(_09276_),
    .A3(net20596),
    .ZN(_09277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18159_ (.A1(net20767),
    .A2(net20818),
    .ZN(_09278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18160_ (.A1(_15608_[0]),
    .A2(net20814),
    .ZN(_09279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _18161_ (.A1(net20481),
    .A2(net20478),
    .A3(net20761),
    .ZN(_09280_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17607 (.I(_15744_[0]),
    .Z(net17607));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18163_ (.A1(_09277_),
    .A2(_09280_),
    .A3(net20654),
    .ZN(_09282_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17678 (.I(_05048_),
    .Z(net17678));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18165_ (.A1(_09274_),
    .A2(_09282_),
    .A3(net20753),
    .ZN(_09284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18166_ (.A1(_09270_),
    .A2(_09284_),
    .A3(net20858),
    .ZN(_09285_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18167_ (.I(_15619_[0]),
    .ZN(_09286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18168_ (.A1(net20814),
    .A2(_09286_),
    .ZN(_09287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18169_ (.A1(_09287_),
    .A2(_07571_),
    .ZN(_09288_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18170_ (.I(_09288_),
    .ZN(_09289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18171_ (.A1(net20769),
    .A2(net20377),
    .ZN(_09290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18172_ (.A1(net19441),
    .A2(net20301),
    .ZN(_09291_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18173_ (.A1(_09291_),
    .A2(net20658),
    .A3(_09240_),
    .ZN(_09292_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18174_ (.I(_15612_[0]),
    .ZN(_09293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18175_ (.A1(_07563_),
    .A2(_09293_),
    .ZN(_09294_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18176_ (.A1(_09294_),
    .A2(_07571_),
    .Z(_09295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18177_ (.A1(_09295_),
    .A2(net20859),
    .Z(_09296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18178_ (.A1(_09239_),
    .A2(net20597),
    .ZN(_09297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18179_ (.A1(_09175_),
    .A2(net20761),
    .ZN(_09298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18180_ (.A1(_09297_),
    .A2(_09298_),
    .Z(_09299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18181_ (.A1(net19440),
    .A2(_09299_),
    .ZN(_09300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18182_ (.A1(_09292_),
    .A2(_09300_),
    .A3(net20755),
    .ZN(_09301_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18183_ (.A1(_09203_),
    .A2(net20301),
    .A3(net20764),
    .Z(_09302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18184_ (.A1(_09172_),
    .A2(net20600),
    .B(net20859),
    .ZN(_09303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18185_ (.A1(_09303_),
    .A2(_09243_),
    .ZN(_09304_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18186_ (.I(_09279_),
    .ZN(_09305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18187_ (.A1(net20299),
    .A2(net20764),
    .ZN(_09306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18188_ (.I(_15633_[0]),
    .ZN(_09307_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18189_ (.A1(net20764),
    .A2(_09307_),
    .B(net20859),
    .ZN(_09308_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18190_ (.I(_09308_),
    .ZN(_09309_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17609 (.I(_15740_[0]),
    .Z(net17609));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18192_ (.A1(_09306_),
    .A2(_09309_),
    .B(net20748),
    .ZN(_09311_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18193_ (.A1(_09302_),
    .A2(_09304_),
    .B(_09311_),
    .ZN(_09312_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18194_ (.A1(_09301_),
    .A2(_09210_),
    .A3(_09312_),
    .ZN(_09313_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18195_ (.A1(_09285_),
    .A2(_09313_),
    .A3(net20857),
    .ZN(_09314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18196_ (.A1(_09260_),
    .A2(_09314_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18197_ (.A1(net19895),
    .A2(_09262_),
    .Z(_09315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18198_ (.A1(_09254_),
    .A2(net20312),
    .A3(net20598),
    .ZN(_09316_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17600 (.I(_15881_[0]),
    .Z(net17600));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18200_ (.A1(_09315_),
    .A2(_09316_),
    .A3(net20660),
    .ZN(_09318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18201_ (.A1(_09278_),
    .A2(net20757),
    .Z(_09319_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _18202_ (.A1(net20862),
    .A2(_09223_),
    .A3(net21123),
    .ZN(_09320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18203_ (.A1(_09319_),
    .A2(net20094),
    .ZN(_09321_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18204_ (.A1(net20758),
    .A2(_15626_[0]),
    .Z(_09322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18205_ (.A1(_09322_),
    .A2(net20859),
    .ZN(_09323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18206_ (.I(_09323_),
    .ZN(_09324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18207_ (.A1(_09321_),
    .A2(_09324_),
    .B(net20750),
    .ZN(_09325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18208_ (.A1(_09318_),
    .A2(_09325_),
    .B(net20858),
    .ZN(_09326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18209_ (.A1(_09224_),
    .A2(net20757),
    .ZN(_09327_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18210_ (.I(_09327_),
    .ZN(_09328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18211_ (.A1(_09328_),
    .A2(net20652),
    .ZN(_09329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18212_ (.A1(net19899),
    .A2(net20487),
    .ZN(_09330_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18213_ (.A1(_09329_),
    .A2(_09330_),
    .A3(net20859),
    .ZN(_09331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18214_ (.A1(_09319_),
    .A2(_09201_),
    .ZN(_09332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18215_ (.A1(net20814),
    .A2(net20300),
    .ZN(_09333_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17756 (.I(_02437_),
    .Z(net17756));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18217_ (.A1(_09333_),
    .A2(net20760),
    .Z(_09335_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18218_ (.A1(_09332_),
    .A2(net20657),
    .A3(_09335_),
    .ZN(_09336_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18219_ (.A1(_09331_),
    .A2(_09336_),
    .A3(net20751),
    .ZN(_09337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18220_ (.A1(_09326_),
    .A2(_09337_),
    .ZN(_09338_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18221_ (.A1(net20767),
    .A2(net20376),
    .Z(_09339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18222_ (.A1(_09339_),
    .A2(net20758),
    .B(net20861),
    .ZN(_09340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18223_ (.A1(_09195_),
    .A2(net20593),
    .ZN(_09341_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18224_ (.I(_09341_),
    .ZN(_09342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18225_ (.A1(net20771),
    .A2(net20616),
    .ZN(_09343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18226_ (.A1(_09342_),
    .A2(net20477),
    .ZN(_09344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18227_ (.A1(_09340_),
    .A2(_09344_),
    .B(net20492),
    .ZN(_09345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18228_ (.A1(_09233_),
    .A2(_09249_),
    .ZN(_09346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18229_ (.A1(_09246_),
    .A2(net20760),
    .ZN(_09347_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18230_ (.A1(_09346_),
    .A2(net20861),
    .A3(net19892),
    .ZN(_09348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18231_ (.A1(_09345_),
    .A2(_09348_),
    .B(_09210_),
    .ZN(_09349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18232_ (.A1(_09228_),
    .A2(net20478),
    .ZN(_09350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18233_ (.A1(net20773),
    .A2(net20811),
    .ZN(_09351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18234_ (.A1(_09253_),
    .A2(_09351_),
    .ZN(_09352_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18235_ (.A1(_09350_),
    .A2(_09352_),
    .A3(net20657),
    .ZN(_09353_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18236_ (.I(_09203_),
    .ZN(_09354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18237_ (.A1(_09354_),
    .A2(net20764),
    .B(net20654),
    .ZN(_09355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18238_ (.A1(_09320_),
    .A2(net20594),
    .ZN(_09356_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18239_ (.I(_09343_),
    .ZN(_09357_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18240_ (.A1(_09356_),
    .A2(_09357_),
    .Z(_09358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18241_ (.A1(net20103),
    .A2(net20759),
    .ZN(_09359_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18242_ (.A1(_09355_),
    .A2(_09358_),
    .A3(_09359_),
    .ZN(_09360_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18243_ (.A1(_09353_),
    .A2(_09360_),
    .A3(net20492),
    .ZN(_09361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18244_ (.A1(_09349_),
    .A2(_09361_),
    .ZN(_09362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18245_ (.A1(_09338_),
    .A2(_09362_),
    .A3(net20857),
    .ZN(_09363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18246_ (.A1(_09246_),
    .A2(net20594),
    .ZN(_09364_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18247_ (.A1(_09364_),
    .A2(net20748),
    .Z(_09365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18248_ (.A1(_09228_),
    .A2(_09180_),
    .ZN(_09366_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18249_ (.A1(_09365_),
    .A2(_09366_),
    .A3(_09335_),
    .ZN(_09367_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18250_ (.A1(_09273_),
    .A2(_09156_),
    .Z(_09368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18251_ (.A1(net20813),
    .A2(net20818),
    .ZN(_09369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18252_ (.A1(_09200_),
    .A2(net20650),
    .ZN(_09370_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18253_ (.A1(_09368_),
    .A2(_09370_),
    .A3(net20493),
    .ZN(_09371_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18254_ (.A1(_09367_),
    .A2(_09371_),
    .A3(net20859),
    .ZN(_09372_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18255_ (.A1(_09245_),
    .A2(_09174_),
    .B(_07571_),
    .ZN(_09373_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18256_ (.A1(net20748),
    .A2(_15635_[0]),
    .A3(net20758),
    .ZN(_09374_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18257_ (.A1(_09373_),
    .A2(_09374_),
    .Z(_09375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18258_ (.A1(_09375_),
    .A2(net20660),
    .B(net20858),
    .ZN(_09376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18259_ (.A1(_09372_),
    .A2(_09376_),
    .B(net20857),
    .ZN(_09377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18260_ (.A1(_09172_),
    .A2(net20597),
    .ZN(_09378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18261_ (.A1(_07571_),
    .A2(_09305_),
    .ZN(_09379_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _18262_ (.A1(net19890),
    .A2(_09355_),
    .A3(_09240_),
    .A4(net20091),
    .ZN(_09380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18263_ (.A1(_09200_),
    .A2(_09180_),
    .ZN(_09381_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18264_ (.A1(_09368_),
    .A2(_09381_),
    .A3(net20657),
    .ZN(_09382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18265_ (.A1(_09380_),
    .A2(net20750),
    .A3(_09382_),
    .ZN(_09383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18266_ (.A1(_09347_),
    .A2(net20654),
    .Z(_09384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18267_ (.A1(net20101),
    .A2(_09203_),
    .Z(_09385_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18268_ (.A1(_09384_),
    .A2(_09385_),
    .B(net20752),
    .ZN(_09386_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18269_ (.A1(net20771),
    .A2(net20371),
    .B(net20757),
    .ZN(_09387_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18270_ (.I(_09387_),
    .ZN(_09388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18271_ (.A1(_09388_),
    .A2(net20303),
    .ZN(_09389_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18272_ (.A1(_09389_),
    .A2(_09344_),
    .A3(net20861),
    .ZN(_09390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18273_ (.A1(_09386_),
    .A2(_09390_),
    .B(_09210_),
    .ZN(_09391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18274_ (.A1(_09383_),
    .A2(_09391_),
    .ZN(_09392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18275_ (.A1(_09377_),
    .A2(_09392_),
    .ZN(_09393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18276_ (.A1(_09363_),
    .A2(_09393_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _18277_ (.A1(_09278_),
    .A2(_09219_),
    .A3(_07571_),
    .Z(_09394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18278_ (.I(_09231_),
    .ZN(_09395_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18279_ (.A1(_09327_),
    .A2(_09395_),
    .ZN(_09396_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18280_ (.A1(_09394_),
    .A2(_09396_),
    .B(net20859),
    .ZN(_09397_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18281_ (.A1(net20096),
    .A2(net20302),
    .A3(_07571_),
    .ZN(_09398_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17601 (.I(_15877_[0]),
    .Z(net17601));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18283_ (.A1(_09280_),
    .A2(_09398_),
    .A3(net20654),
    .ZN(_09400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18284_ (.A1(_09397_),
    .A2(net20498),
    .A3(_09400_),
    .ZN(_09401_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18285_ (.A1(_09254_),
    .A2(net20491),
    .A3(net20593),
    .ZN(_09402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18286_ (.A1(_09219_),
    .A2(net20758),
    .ZN(_09403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18287_ (.A1(_09402_),
    .A2(_09403_),
    .ZN(_09404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18288_ (.A1(_09404_),
    .A2(net20654),
    .ZN(_09405_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18289_ (.A1(net20502),
    .A2(_09343_),
    .A3(net20763),
    .ZN(_09406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18290_ (.A1(net20815),
    .A2(net20371),
    .ZN(_09407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18291_ (.A1(net20489),
    .A2(_09407_),
    .A3(net20598),
    .ZN(_09408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18292_ (.A1(_09406_),
    .A2(_09408_),
    .A3(net20859),
    .ZN(_09409_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18293_ (.A1(_09405_),
    .A2(_09409_),
    .A3(net20748),
    .ZN(_09410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18294_ (.A1(_09401_),
    .A2(_09410_),
    .A3(_09210_),
    .ZN(_09411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18295_ (.A1(_09262_),
    .A2(_09356_),
    .ZN(_09412_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18296_ (.A1(_09249_),
    .A2(net20654),
    .Z(_09413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18297_ (.A1(_09267_),
    .A2(_09186_),
    .ZN(_09414_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18298_ (.A1(_09412_),
    .A2(_09413_),
    .B(_09414_),
    .ZN(_09415_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18299_ (.A1(_09275_),
    .A2(net20596),
    .A3(_09320_),
    .Z(_09416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18300_ (.A1(net20814),
    .A2(net20615),
    .ZN(_09417_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18301_ (.I(_09417_),
    .ZN(_09418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18302_ (.A1(_09418_),
    .A2(net20765),
    .ZN(_09419_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18303_ (.I(_09419_),
    .ZN(_09420_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18304_ (.A1(_09416_),
    .A2(_09420_),
    .B(net20859),
    .ZN(_09421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18305_ (.A1(_09415_),
    .A2(_09421_),
    .B(_09210_),
    .ZN(_09422_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18306_ (.A1(_09179_),
    .A2(net20478),
    .Z(_09423_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18307_ (.A1(_09275_),
    .A2(net20763),
    .A3(net20097),
    .Z(_09424_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18308_ (.A1(_09423_),
    .A2(_09424_),
    .B(net20656),
    .ZN(_09425_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18309_ (.A1(_09199_),
    .A2(_09418_),
    .B(net20859),
    .ZN(_09426_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18310_ (.A1(_09155_),
    .A2(_09265_),
    .A3(net20597),
    .Z(_09427_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18311_ (.A1(_09426_),
    .A2(_09427_),
    .Z(_09428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18312_ (.A1(_09425_),
    .A2(_09428_),
    .A3(net20753),
    .ZN(_09429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18313_ (.A1(_09429_),
    .A2(_09422_),
    .ZN(_09430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18314_ (.A1(_09411_),
    .A2(_09430_),
    .ZN(_09431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18315_ (.A1(_09431_),
    .A2(_09213_),
    .ZN(_09432_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18316_ (.A1(net20757),
    .A2(_15631_[0]),
    .Z(_09433_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18317_ (.A1(_09403_),
    .A2(net20659),
    .A3(_09433_),
    .Z(_09434_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18318_ (.A1(_09434_),
    .A2(net20749),
    .ZN(_09435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18319_ (.A1(net20765),
    .A2(_15628_[0]),
    .ZN(_09436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18320_ (.A1(_09436_),
    .A2(net20859),
    .ZN(_09437_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18321_ (.A1(_09394_),
    .A2(_09437_),
    .Z(_09438_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18322_ (.A1(_09435_),
    .A2(_09438_),
    .B(net20858),
    .ZN(_09439_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18323_ (.A1(_09342_),
    .A2(net20489),
    .Z(_09440_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18324_ (.A1(_09440_),
    .A2(net20659),
    .A3(_09373_),
    .Z(_09441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18325_ (.A1(_09179_),
    .A2(net20093),
    .ZN(_09442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18326_ (.A1(_09172_),
    .A2(net20761),
    .B(net20859),
    .ZN(_09443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18327_ (.A1(_09442_),
    .A2(_09443_),
    .B(_09186_),
    .ZN(_09444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18328_ (.A1(_09441_),
    .A2(_09444_),
    .ZN(_09445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18329_ (.A1(_09439_),
    .A2(_09445_),
    .B(_09213_),
    .ZN(_09446_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18330_ (.A1(_09201_),
    .A2(net20479),
    .A3(net20595),
    .ZN(_09447_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18331_ (.A1(net20369),
    .A2(net20593),
    .B(_09447_),
    .C(net20661),
    .ZN(_09448_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18332_ (.A1(net20092),
    .A2(net20859),
    .Z(_09449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18333_ (.A1(_09250_),
    .A2(_09180_),
    .ZN(_09450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18334_ (.A1(_09190_),
    .A2(net20597),
    .ZN(_09451_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18335_ (.A1(_09449_),
    .A2(_09450_),
    .A3(_09451_),
    .ZN(_09452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18336_ (.A1(_09448_),
    .A2(_09452_),
    .A3(_09186_),
    .ZN(_09453_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18337_ (.A1(_09290_),
    .A2(net20601),
    .Z(_09454_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18338_ (.I(_09454_),
    .ZN(_09455_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18339_ (.I(_09165_),
    .ZN(_09456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18340_ (.A1(net20764),
    .A2(net20370),
    .ZN(_09457_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18341_ (.A1(_09455_),
    .A2(net20089),
    .B(net20654),
    .C(_09457_),
    .ZN(_09458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18342_ (.I(_09198_),
    .ZN(_09459_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18343_ (.A1(net20296),
    .A2(_15628_[0]),
    .B(net20598),
    .ZN(_09460_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18344_ (.A1(_09460_),
    .A2(net20859),
    .A3(_09280_),
    .ZN(_09461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18345_ (.A1(_09458_),
    .A2(net20755),
    .A3(_09461_),
    .ZN(_09462_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18346_ (.A1(_09453_),
    .A2(_09462_),
    .A3(net20858),
    .ZN(_09463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18347_ (.A1(_09446_),
    .A2(_09463_),
    .ZN(_09464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18348_ (.A1(_09432_),
    .A2(_09464_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18349_ (.A1(_09200_),
    .A2(net20488),
    .ZN(_09465_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18350_ (.A1(net20503),
    .A2(net20314),
    .A3(net20597),
    .ZN(_09466_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18351_ (.A1(_09465_),
    .A2(net20656),
    .A3(_09466_),
    .ZN(_09467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18352_ (.I(_15628_[0]),
    .ZN(_09468_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18353_ (.A1(net20490),
    .A2(_09468_),
    .A3(net20766),
    .ZN(_09469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18354_ (.A1(_09456_),
    .A2(net20597),
    .ZN(_09470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18355_ (.A1(_09469_),
    .A2(_09470_),
    .ZN(_09471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18356_ (.A1(_09471_),
    .A2(net20861),
    .ZN(_09472_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18357_ (.A1(_09467_),
    .A2(net20500),
    .A3(_09472_),
    .ZN(_09473_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18358_ (.A1(net20653),
    .A2(_09189_),
    .A3(net20766),
    .ZN(_09474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18359_ (.A1(_09474_),
    .A2(_09168_),
    .ZN(_09475_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18360_ (.A1(_09378_),
    .A2(net20859),
    .Z(_09476_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18361_ (.A1(_09475_),
    .A2(_09476_),
    .ZN(_09477_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18362_ (.A1(_09254_),
    .A2(net20095),
    .A3(net20597),
    .ZN(_09478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18363_ (.A1(_09406_),
    .A2(_09478_),
    .A3(net20654),
    .ZN(_09479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18364_ (.A1(_09477_),
    .A2(net20754),
    .A3(_09479_),
    .ZN(_09480_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18365_ (.A1(_09473_),
    .A2(_09480_),
    .A3(_09210_),
    .ZN(_09481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18366_ (.A1(_09220_),
    .A2(net20654),
    .Z(_09482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18367_ (.A1(_09465_),
    .A2(_09482_),
    .B(net20754),
    .ZN(_09483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18368_ (.A1(net20097),
    .A2(net20757),
    .ZN(_09484_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18369_ (.I(_09484_),
    .ZN(_09485_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18370_ (.A1(_09485_),
    .A2(net20476),
    .ZN(_09486_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18371_ (.A1(_09346_),
    .A2(_09486_),
    .A3(net20861),
    .ZN(_09487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18372_ (.A1(_09483_),
    .A2(_09487_),
    .B(_09210_),
    .ZN(_09488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18373_ (.A1(_09189_),
    .A2(_09333_),
    .B(net20766),
    .ZN(_09489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18374_ (.A1(_09245_),
    .A2(net20478),
    .B(net20597),
    .ZN(_09490_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18375_ (.A1(_09489_),
    .A2(_09490_),
    .B(net20654),
    .ZN(_09491_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18376_ (.A1(net20314),
    .A2(net20102),
    .A3(net20766),
    .ZN(_09492_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18377_ (.A1(_09206_),
    .A2(_09492_),
    .A3(net20861),
    .ZN(_09493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18378_ (.A1(_09491_),
    .A2(_09493_),
    .ZN(_09494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18379_ (.A1(_09494_),
    .A2(net20754),
    .ZN(_09495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18380_ (.A1(_09488_),
    .A2(_09495_),
    .ZN(_09496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18381_ (.A1(_09481_),
    .A2(_09496_),
    .B(_09213_),
    .ZN(_09497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18382_ (.A1(_09194_),
    .A2(_09215_),
    .ZN(_09498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18383_ (.A1(_09233_),
    .A2(net20490),
    .ZN(_09499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18384_ (.A1(_09498_),
    .A2(_09499_),
    .A3(net20495),
    .ZN(_09500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18385_ (.A1(_09266_),
    .A2(net20597),
    .ZN(_09501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18386_ (.A1(_09501_),
    .A2(net20748),
    .ZN(_09502_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18387_ (.A1(_09424_),
    .A2(_09502_),
    .Z(_09503_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18388_ (.A1(_09500_),
    .A2(_09503_),
    .B(net20861),
    .ZN(_09504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18389_ (.A1(_09249_),
    .A2(net20102),
    .B(net20597),
    .ZN(_09505_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18390_ (.I(_09470_),
    .ZN(_09506_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18391_ (.A1(_09505_),
    .A2(_09506_),
    .B(net20499),
    .ZN(_09507_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18392_ (.A1(_09164_),
    .A2(_09186_),
    .ZN(_09508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18393_ (.A1(_09297_),
    .A2(net20859),
    .ZN(_09509_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18394_ (.A1(_09508_),
    .A2(_09509_),
    .ZN(_09510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18395_ (.A1(_09507_),
    .A2(_09510_),
    .ZN(_09511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18396_ (.A1(_09511_),
    .A2(_09210_),
    .ZN(_09512_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18397_ (.A1(_09504_),
    .A2(_09512_),
    .B(_09213_),
    .ZN(_09513_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18398_ (.A1(_09288_),
    .A2(_09459_),
    .ZN(_09514_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18399_ (.A1(_09514_),
    .A2(_09373_),
    .B(net20654),
    .ZN(_09515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18400_ (.A1(_09515_),
    .A2(_09426_),
    .ZN(_09516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18401_ (.A1(_09516_),
    .A2(net20500),
    .ZN(_09517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18402_ (.A1(_09332_),
    .A2(_09303_),
    .A3(_09243_),
    .ZN(_09518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18403_ (.A1(_09194_),
    .A2(net20306),
    .ZN(_09519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18404_ (.A1(_09215_),
    .A2(_09265_),
    .ZN(_09520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18405_ (.A1(_09520_),
    .A2(net20597),
    .ZN(_09521_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18406_ (.A1(_09519_),
    .A2(net20861),
    .A3(_09521_),
    .ZN(_09522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18407_ (.A1(_09518_),
    .A2(_09522_),
    .A3(net20752),
    .ZN(_09523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18408_ (.A1(_09517_),
    .A2(_09523_),
    .B(_09210_),
    .ZN(_09524_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18409_ (.A1(_09513_),
    .A2(_09524_),
    .ZN(_09525_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18410_ (.A1(_09497_),
    .A2(_09525_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18411_ (.A1(_09396_),
    .A2(net20654),
    .ZN(_09526_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18412_ (.A1(net20315),
    .A2(_09455_),
    .B(_09526_),
    .ZN(_09527_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18413_ (.A1(_09369_),
    .A2(net20759),
    .Z(_09528_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18414_ (.A1(_09315_),
    .A2(_09303_),
    .A3(_09528_),
    .ZN(_09529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18415_ (.A1(_09527_),
    .A2(_09529_),
    .A3(net20498),
    .ZN(_09530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18416_ (.A1(_09379_),
    .A2(_09265_),
    .Z(_09531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18417_ (.A1(_09264_),
    .A2(_09531_),
    .B(_09186_),
    .ZN(_09532_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18418_ (.A1(_09254_),
    .A2(net20762),
    .Z(_09533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18419_ (.A1(_09533_),
    .A2(net20313),
    .ZN(_09534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18420_ (.A1(_09534_),
    .A2(_09291_),
    .A3(net20658),
    .ZN(_09535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18421_ (.A1(_09532_),
    .A2(_09535_),
    .B(_09213_),
    .ZN(_09536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18422_ (.A1(_09530_),
    .A2(_09536_),
    .ZN(_09537_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18423_ (.I(_09514_),
    .ZN(_09538_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18424_ (.A1(net20502),
    .A2(_09204_),
    .Z(_09539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18425_ (.A1(_09539_),
    .A2(net20762),
    .ZN(_09540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18426_ (.A1(_09538_),
    .A2(_09540_),
    .A3(net20859),
    .ZN(_09541_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18427_ (.A1(_09272_),
    .A2(net20658),
    .A3(_09206_),
    .ZN(_09542_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18428_ (.A1(_09541_),
    .A2(_09542_),
    .A3(_09186_),
    .ZN(_09543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18429_ (.A1(_09289_),
    .A2(_09249_),
    .ZN(_09544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18430_ (.A1(_09296_),
    .A2(_09544_),
    .Z(_09545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18431_ (.A1(net20757),
    .A2(net20617),
    .ZN(_09546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18432_ (.A1(_09379_),
    .A2(_09546_),
    .ZN(_09547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18433_ (.A1(_09547_),
    .A2(net20654),
    .ZN(_09548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18434_ (.A1(_09548_),
    .A2(net20748),
    .ZN(_09549_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18435_ (.A1(_09545_),
    .A2(_09549_),
    .Z(_09550_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18436_ (.A1(_09543_),
    .A2(_09550_),
    .A3(_09213_),
    .ZN(_09551_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18437_ (.A1(_09537_),
    .A2(_09551_),
    .A3(_09210_),
    .ZN(_09552_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18438_ (.A1(net20484),
    .A2(_09180_),
    .A3(net20595),
    .ZN(_09553_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18439_ (.A1(net20595),
    .A2(_09539_),
    .B(_09553_),
    .C(net20859),
    .ZN(_09554_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18440_ (.A1(_09370_),
    .A2(net20660),
    .A3(_09447_),
    .ZN(_09555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18441_ (.A1(_09554_),
    .A2(_09555_),
    .A3(net20492),
    .ZN(_09556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18442_ (.A1(net20597),
    .A2(_15637_[0]),
    .ZN(_09557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18443_ (.A1(_09557_),
    .A2(net20654),
    .ZN(_09558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18444_ (.A1(net20767),
    .A2(_09242_),
    .B(_09558_),
    .ZN(_09559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18445_ (.A1(_09559_),
    .A2(_09366_),
    .ZN(_09560_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18446_ (.A1(net20305),
    .A2(net20654),
    .ZN(_09561_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18447_ (.A1(_09561_),
    .A2(net19896),
    .B(_09186_),
    .ZN(_09562_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18448_ (.A1(_09560_),
    .A2(_09562_),
    .B(_09213_),
    .ZN(_09563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18449_ (.A1(_09556_),
    .A2(_09563_),
    .ZN(_09564_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18450_ (.A1(_09159_),
    .A2(net20859),
    .Z(_09565_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18451_ (.A1(_09565_),
    .A2(_09359_),
    .A3(_09368_),
    .ZN(_09566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18452_ (.A1(_09200_),
    .A2(net20307),
    .ZN(_09567_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18453_ (.A1(net20595),
    .A2(net20813),
    .B(net20859),
    .ZN(_09568_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18454_ (.A1(_09567_),
    .A2(_09568_),
    .B(net20750),
    .ZN(_09569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18455_ (.A1(_09566_),
    .A2(_09569_),
    .ZN(_09570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18456_ (.A1(_09341_),
    .A2(net20859),
    .Z(_09571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18457_ (.A1(_09571_),
    .A2(net20297),
    .B(_09186_),
    .ZN(_09572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18458_ (.A1(_09328_),
    .A2(net20478),
    .ZN(_09573_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18459_ (.A1(_09573_),
    .A2(_09247_),
    .A3(_09243_),
    .ZN(_09574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18460_ (.A1(_09572_),
    .A2(_09574_),
    .ZN(_09575_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18461_ (.A1(_09570_),
    .A2(_09575_),
    .A3(_09213_),
    .ZN(_09576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18462_ (.A1(_09564_),
    .A2(_09576_),
    .A3(net20858),
    .ZN(_09577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18463_ (.A1(_09552_),
    .A2(_09577_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18464_ (.A1(net20490),
    .A2(net20594),
    .ZN(_09578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18465_ (.A1(_09384_),
    .A2(_09333_),
    .A3(net20295),
    .ZN(_09579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18466_ (.A1(_09264_),
    .A2(net20099),
    .ZN(_09580_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18467_ (.A1(_09579_),
    .A2(net20752),
    .A3(_09580_),
    .ZN(_09581_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18468_ (.A1(_09164_),
    .A2(_09419_),
    .A3(net20859),
    .Z(_09582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18469_ (.A1(net19900),
    .A2(_09276_),
    .ZN(_09583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18470_ (.A1(_09582_),
    .A2(_09583_),
    .ZN(_09584_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18471_ (.A1(net20475),
    .A2(net20815),
    .B1(net20311),
    .B2(net20757),
    .ZN(_09585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18472_ (.A1(_09585_),
    .A2(net20654),
    .B(net20748),
    .ZN(_09586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18473_ (.A1(_09584_),
    .A2(_09586_),
    .ZN(_09587_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18474_ (.A1(_09581_),
    .A2(_09587_),
    .A3(_09210_),
    .ZN(_09588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18475_ (.A1(_09347_),
    .A2(_09419_),
    .Z(_09589_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18476_ (.A1(_09175_),
    .A2(net20594),
    .B(net20654),
    .ZN(_09590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18477_ (.A1(_09589_),
    .A2(_09590_),
    .B(net20752),
    .ZN(_09591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18478_ (.A1(net20309),
    .A2(net20094),
    .ZN(_09592_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18479_ (.A1(_09592_),
    .A2(_09247_),
    .A3(_09243_),
    .ZN(_09593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18480_ (.A1(_09591_),
    .A2(_09593_),
    .B(_09210_),
    .ZN(_09594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18481_ (.A1(_09221_),
    .A2(net20314),
    .ZN(_09595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18482_ (.A1(_09485_),
    .A2(_09249_),
    .ZN(_09596_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18483_ (.A1(_09595_),
    .A2(_09596_),
    .A3(net20861),
    .ZN(_09597_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18484_ (.I(net20304),
    .ZN(_09598_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18485_ (.A1(_09202_),
    .A2(net20657),
    .A3(_09598_),
    .ZN(_09599_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18486_ (.A1(_09597_),
    .A2(_09599_),
    .A3(net20752),
    .ZN(_09600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18487_ (.A1(_09594_),
    .A2(_09600_),
    .ZN(_09601_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18488_ (.A1(_09588_),
    .A2(_09601_),
    .A3(_09213_),
    .ZN(_09602_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18489_ (.A1(net19893),
    .A2(_09333_),
    .Z(_09603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18490_ (.A1(_09603_),
    .A2(net20861),
    .B(net20752),
    .ZN(_09604_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18491_ (.I(_09194_),
    .ZN(_09605_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18492_ (.A1(_09521_),
    .A2(_09605_),
    .A3(net20655),
    .ZN(_09606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18493_ (.A1(_09604_),
    .A2(_09606_),
    .B(_09210_),
    .ZN(_09607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18494_ (.A1(_09233_),
    .A2(net20100),
    .ZN(_09608_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18495_ (.A1(_09241_),
    .A2(net20655),
    .A3(_09608_),
    .ZN(_09609_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18496_ (.I(_09578_),
    .ZN(_09610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18497_ (.A1(_09610_),
    .A2(net20095),
    .ZN(_09611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18498_ (.A1(_09485_),
    .A2(net20301),
    .ZN(_09612_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18499_ (.A1(_09611_),
    .A2(_09612_),
    .A3(net20861),
    .ZN(_09613_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18500_ (.A1(_09609_),
    .A2(_09613_),
    .A3(net20752),
    .ZN(_09614_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18501_ (.A1(_09607_),
    .A2(_09614_),
    .B(_09213_),
    .ZN(_09615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18502_ (.A1(net20759),
    .A2(net20811),
    .ZN(_09616_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18503_ (.A1(net20315),
    .A2(net20759),
    .B1(_09616_),
    .B2(net20818),
    .ZN(_09617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18504_ (.A1(_09617_),
    .A2(net20655),
    .ZN(_09618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18505_ (.A1(net20308),
    .A2(_09351_),
    .ZN(_09619_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18506_ (.A1(_09619_),
    .A2(_09590_),
    .A3(net19891),
    .ZN(_09620_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18507_ (.A1(_09618_),
    .A2(_09620_),
    .A3(net20752),
    .ZN(_09621_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18508_ (.A1(_09343_),
    .A2(net20598),
    .Z(_09622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18509_ (.A1(_09622_),
    .A2(_09180_),
    .ZN(_09623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18510_ (.A1(_09623_),
    .A2(net20654),
    .A3(_09419_),
    .ZN(_09624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18511_ (.A1(_09388_),
    .A2(net20480),
    .ZN(_09625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18512_ (.A1(_09449_),
    .A2(_09625_),
    .ZN(_09626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18513_ (.A1(_09624_),
    .A2(_09626_),
    .A3(net20494),
    .ZN(_09627_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18514_ (.A1(_09621_),
    .A2(_09627_),
    .A3(_09210_),
    .ZN(_09628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18515_ (.A1(_09615_),
    .A2(_09628_),
    .ZN(_09629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18516_ (.A1(_09602_),
    .A2(_09629_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18517_ (.A1(_09200_),
    .A2(net20478),
    .ZN(_09630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18518_ (.A1(_09454_),
    .A2(net20652),
    .ZN(_09631_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18519_ (.A1(_09630_),
    .A2(_09631_),
    .A3(net20662),
    .ZN(_09632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18520_ (.A1(_09454_),
    .A2(net20651),
    .ZN(_09633_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18521_ (.A1(_09633_),
    .A2(net20860),
    .A3(net19439),
    .ZN(_09634_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18522_ (.A1(_09632_),
    .A2(_09634_),
    .A3(net20497),
    .ZN(_09635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18523_ (.A1(_09388_),
    .A2(net20477),
    .ZN(_09636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18524_ (.A1(_09221_),
    .A2(net20483),
    .ZN(_09637_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18525_ (.A1(_09636_),
    .A2(_09637_),
    .A3(net20654),
    .ZN(_09638_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18526_ (.A1(net20090),
    .A2(net20104),
    .B(net20860),
    .C(_09433_),
    .ZN(_09639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18527_ (.A1(_09638_),
    .A2(net20749),
    .A3(_09639_),
    .ZN(_09640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18528_ (.A1(_09635_),
    .A2(_09640_),
    .A3(net20857),
    .ZN(_09641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18529_ (.A1(_09276_),
    .A2(net20761),
    .ZN(_09642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18530_ (.A1(net18949),
    .A2(_09642_),
    .B(net20654),
    .ZN(_09643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18531_ (.A1(_09398_),
    .A2(net20654),
    .ZN(_09644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18532_ (.A1(_09644_),
    .A2(net20498),
    .ZN(_09645_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18533_ (.A1(_09643_),
    .A2(_09645_),
    .ZN(_09646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18534_ (.A1(_09622_),
    .A2(net20307),
    .ZN(_09647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18535_ (.A1(_09355_),
    .A2(_09647_),
    .ZN(_09648_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18536_ (.A1(_15627_[0]),
    .A2(net20758),
    .B(net20659),
    .ZN(_09649_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18537_ (.I(_09649_),
    .ZN(_09650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18538_ (.A1(_09596_),
    .A2(_09650_),
    .ZN(_09651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18539_ (.A1(_09648_),
    .A2(_09651_),
    .B(net20494),
    .ZN(_09652_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18540_ (.A1(_09646_),
    .A2(_09652_),
    .B(_09213_),
    .ZN(_09653_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18541_ (.A1(_09641_),
    .A2(_09653_),
    .A3(_09210_),
    .ZN(_09654_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18542_ (.I(_09407_),
    .ZN(_09655_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18543_ (.A1(net20098),
    .A2(_09655_),
    .B(net20601),
    .ZN(_09656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18544_ (.A1(_09172_),
    .A2(net20764),
    .B(net20654),
    .ZN(_09657_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18545_ (.A1(_09656_),
    .A2(_09657_),
    .B(_09186_),
    .ZN(_09658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18546_ (.A1(_09539_),
    .A2(net20600),
    .ZN(_09659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18547_ (.A1(net20773),
    .A2(net20764),
    .ZN(_09660_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18548_ (.A1(_09659_),
    .A2(net20654),
    .A3(_09660_),
    .ZN(_09661_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18549_ (.A1(_09658_),
    .A2(_09661_),
    .B(_09213_),
    .ZN(_09662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18550_ (.A1(_09297_),
    .A2(net20654),
    .Z(_09663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18551_ (.A1(_09485_),
    .A2(_09254_),
    .ZN(_09664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18552_ (.A1(net20601),
    .A2(net20485),
    .ZN(_09665_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18553_ (.A1(_09665_),
    .A2(net20772),
    .Z(_09666_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18554_ (.A1(_09663_),
    .A2(_09664_),
    .A3(_09666_),
    .ZN(_09667_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18555_ (.A1(_09630_),
    .A2(_09521_),
    .A3(net20860),
    .ZN(_09668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18556_ (.A1(_09667_),
    .A2(_09668_),
    .A3(net20501),
    .ZN(_09669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18557_ (.A1(_09662_),
    .A2(_09669_),
    .B(_09210_),
    .ZN(_09670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18558_ (.A1(_09250_),
    .A2(_09333_),
    .ZN(_09671_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18559_ (.A1(_09201_),
    .A2(net20652),
    .A3(_07571_),
    .ZN(_09672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18560_ (.A1(_09671_),
    .A2(_09672_),
    .ZN(_09673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18561_ (.A1(_09673_),
    .A2(net20661),
    .ZN(_09674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18562_ (.A1(_09533_),
    .A2(_09203_),
    .ZN(_09675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18563_ (.A1(_09675_),
    .A2(net20859),
    .A3(_09672_),
    .ZN(_09676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18564_ (.A1(_09674_),
    .A2(_09676_),
    .A3(net20749),
    .ZN(_09677_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18565_ (.A1(_09229_),
    .A2(net20859),
    .A3(_09322_),
    .ZN(_09678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18566_ (.A1(_09357_),
    .A2(net20759),
    .ZN(_09679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18567_ (.A1(_09521_),
    .A2(net20657),
    .A3(_09679_),
    .ZN(_09680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18568_ (.A1(_09678_),
    .A2(net20492),
    .A3(_09680_),
    .ZN(_09681_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18569_ (.A1(_09677_),
    .A2(_09681_),
    .A3(_09213_),
    .ZN(_09682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18570_ (.A1(_09670_),
    .A2(_09682_),
    .ZN(_09683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18571_ (.A1(_09654_),
    .A2(_09683_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18572_ (.A1(net20764),
    .A2(_09655_),
    .B(_09172_),
    .ZN(_09684_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18573_ (.A1(net20315),
    .A2(net20595),
    .ZN(_09685_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18574_ (.A1(_09684_),
    .A2(net20662),
    .A3(_09685_),
    .ZN(_09686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18575_ (.A1(net20764),
    .A2(net20376),
    .ZN(_09687_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18576_ (.A1(_09659_),
    .A2(net20859),
    .A3(_09687_),
    .ZN(_09688_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18577_ (.A1(_09686_),
    .A2(_09688_),
    .A3(net20497),
    .ZN(_09689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18578_ (.A1(net20298),
    .A2(net20491),
    .ZN(_09690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18579_ (.A1(_09538_),
    .A2(_09690_),
    .A3(net20860),
    .ZN(_09691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18580_ (.A1(net20477),
    .A2(_09276_),
    .A3(_07571_),
    .ZN(_09692_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18581_ (.A1(_07571_),
    .A2(net20617),
    .A3(net20767),
    .Z(_09693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18582_ (.A1(_09443_),
    .A2(_09692_),
    .A3(_09693_),
    .ZN(_09694_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18583_ (.A1(_09691_),
    .A2(_09694_),
    .A3(net20749),
    .ZN(_09695_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18584_ (.A1(_09689_),
    .A2(_09695_),
    .A3(net20858),
    .ZN(_09696_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18585_ (.I(_09267_),
    .ZN(_09697_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18586_ (.A1(_09697_),
    .A2(_09558_),
    .ZN(_09698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18587_ (.A1(net20089),
    .A2(net20765),
    .ZN(_09699_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18588_ (.A1(_09698_),
    .A2(_09699_),
    .B(net20755),
    .ZN(_09700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18589_ (.A1(_09622_),
    .A2(net20313),
    .ZN(_09701_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18590_ (.A1(_09355_),
    .A2(_09701_),
    .A3(_09457_),
    .ZN(_09702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18591_ (.A1(_09700_),
    .A2(_09702_),
    .ZN(_09703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18592_ (.A1(_09565_),
    .A2(net19894),
    .A3(_09368_),
    .ZN(_09704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18593_ (.A1(_09665_),
    .A2(net20654),
    .ZN(_09705_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18594_ (.I(_09705_),
    .ZN(_09706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18595_ (.A1(_09655_),
    .A2(net20764),
    .ZN(_09707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18596_ (.A1(_09706_),
    .A2(_09707_),
    .B(_09186_),
    .ZN(_09708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18597_ (.A1(_09704_),
    .A2(_09708_),
    .ZN(_09709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18598_ (.A1(_09703_),
    .A2(_09210_),
    .A3(_09709_),
    .ZN(_09710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18599_ (.A1(_09696_),
    .A2(_09710_),
    .A3(net20857),
    .ZN(_09711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18600_ (.A1(_09216_),
    .A2(net20301),
    .ZN(_09712_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18601_ (.A1(_09476_),
    .A2(_09666_),
    .A3(_09712_),
    .ZN(_09713_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18602_ (.A1(_09533_),
    .A2(net20859),
    .ZN(_09714_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18603_ (.A1(_09714_),
    .A2(net18949),
    .B(_09186_),
    .ZN(_09715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18604_ (.A1(_09713_),
    .A2(_09715_),
    .B(_09210_),
    .ZN(_09716_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18605_ (.A1(_09460_),
    .A2(_09664_),
    .A3(net20654),
    .ZN(_09717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18606_ (.A1(_09498_),
    .A2(net20859),
    .A3(_09316_),
    .ZN(_09718_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18607_ (.A1(_09717_),
    .A2(_09718_),
    .A3(net20501),
    .ZN(_09719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18608_ (.A1(_09716_),
    .A2(_09719_),
    .ZN(_09720_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18609_ (.A1(net20477),
    .A2(net20491),
    .A3(net20761),
    .ZN(_09721_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18610_ (.A1(_09455_),
    .A2(_09721_),
    .A3(net20860),
    .ZN(_09722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18611_ (.A1(_09247_),
    .A2(net19901),
    .ZN(_09723_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18612_ (.A1(_09722_),
    .A2(_09723_),
    .A3(net20497),
    .ZN(_09724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18613_ (.A1(_09610_),
    .A2(net20503),
    .ZN(_09725_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18614_ (.A1(_09616_),
    .A2(net20859),
    .Z(_09726_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18615_ (.A1(_09725_),
    .A2(_09726_),
    .B(net20494),
    .ZN(_09727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18616_ (.A1(_09250_),
    .A2(net20491),
    .ZN(_09728_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18617_ (.A1(_09728_),
    .A2(net20661),
    .A3(_09447_),
    .ZN(_09729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18618_ (.A1(_09727_),
    .A2(_09729_),
    .ZN(_09730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18619_ (.A1(_09724_),
    .A2(_09730_),
    .A3(_09210_),
    .ZN(_09731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18620_ (.A1(_09720_),
    .A2(_09731_),
    .A3(_09213_),
    .ZN(_09732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18621_ (.A1(_09711_),
    .A2(_09732_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18622_ (.I(_15650_[0]),
    .ZN(_15639_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18623_ (.A1(net21540),
    .A2(net47),
    .ZN(_09733_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _18624_ (.A1(_07694_),
    .A2(net21540),
    .B(_09733_),
    .ZN(_09734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17594 (.I(_10623_),
    .Z(net17594));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18626_ (.A1(_07679_),
    .A2(net21526),
    .ZN(_09735_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18627_ (.I(_07680_),
    .ZN(_09736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18628_ (.A1(_09736_),
    .A2(_09735_),
    .ZN(_15640_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18629_ (.A1(_07706_),
    .A2(net20697),
    .ZN(_09737_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18630_ (.I(_09737_),
    .ZN(_09738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18631_ (.A1(_09738_),
    .A2(net664),
    .Z(_09739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18632_ (.I(_15641_[0]),
    .ZN(_09740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18633_ (.A1(net20810),
    .A2(_09740_),
    .ZN(_09741_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _18634_ (.I(_07706_),
    .ZN(_09742_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18635_ (.A1(_09741_),
    .A2(_09742_),
    .B(net20669),
    .ZN(_09743_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18636_ (.A1(_09739_),
    .A2(_09743_),
    .ZN(_09744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18637_ (.I(_09744_),
    .ZN(_09745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18638_ (.A1(net20810),
    .A2(net20152),
    .ZN(_09746_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18639_ (.I(_09746_),
    .ZN(_09747_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17603 (.I(_15869_[0]),
    .Z(net17603));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18641_ (.A1(_09747_),
    .A2(net20464),
    .ZN(_09749_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17593 (.I(_10652_),
    .Z(net17593));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18643_ (.I(_15642_[0]),
    .ZN(_09751_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _18644_ (.A1(_09751_),
    .A2(net21110),
    .A3(net20843),
    .ZN(_09752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18645_ (.A1(_09752_),
    .A2(_07706_),
    .ZN(_09753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18646_ (.A1(_09749_),
    .A2(_07717_),
    .A3(net19437),
    .ZN(_09754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18647_ (.A1(_09745_),
    .A2(_09754_),
    .ZN(_09755_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17599 (.I(_10500_),
    .Z(net17599));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18649_ (.A1(net20701),
    .A2(net20154),
    .ZN(_09757_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18650_ (.I(_09757_),
    .ZN(_09758_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17602 (.I(net423),
    .Z(net17602));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18652_ (.A1(_09758_),
    .A2(net20465),
    .ZN(_09760_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18653_ (.A1(_09760_),
    .A2(net20668),
    .Z(_09761_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _18654_ (.I(net20837),
    .ZN(_09762_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17825 (.I(net17820),
    .Z(net17825));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18656_ (.A1(_09755_),
    .A2(_09761_),
    .B(_09762_),
    .ZN(_09764_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18657_ (.I(_15655_[0]),
    .ZN(_09765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18658_ (.A1(net20697),
    .A2(_09765_),
    .ZN(_09766_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18659_ (.I(_09766_),
    .ZN(_09767_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18660_ (.A1(net20810),
    .A2(_15657_[0]),
    .Z(_09768_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17592 (.I(_10767_),
    .Z(net17592));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18662_ (.A1(_09767_),
    .A2(_09768_),
    .B(net20461),
    .ZN(_09770_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18663_ (.I(_15648_[0]),
    .ZN(_09771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18664_ (.A1(net20810),
    .A2(_09771_),
    .ZN(_09772_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17596 (.I(_10562_),
    .Z(net17596));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18666_ (.A1(_09772_),
    .A2(net20685),
    .ZN(_09774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18667_ (.A1(_09770_),
    .A2(net19436),
    .ZN(_09775_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17597 (.I(_10562_),
    .Z(net17597));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18669_ (.A1(_09775_),
    .A2(_07717_),
    .ZN(_09777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18670_ (.A1(net20474),
    .A2(net20810),
    .ZN(_09778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18671_ (.A1(net20156),
    .A2(net20697),
    .ZN(_09779_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18672_ (.A1(_09778_),
    .A2(net20082),
    .A3(net20461),
    .ZN(_09780_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18673_ (.I(_09780_),
    .ZN(_09781_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18674_ (.I(_15651_[0]),
    .ZN(_09782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18675_ (.A1(net20697),
    .A2(_09782_),
    .ZN(_09783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18676_ (.A1(net20472),
    .A2(net20810),
    .ZN(_09784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18677_ (.A1(net19885),
    .A2(net20291),
    .B(net20462),
    .ZN(_09785_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17585 (.I(_11293_),
    .Z(net17585));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17590 (.I(_11245_),
    .Z(net17590));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18680_ (.A1(_09781_),
    .A2(_09785_),
    .B(net20672),
    .ZN(_09788_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17584 (.I(_11327_),
    .Z(net17584));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18682_ (.A1(_09777_),
    .A2(_09788_),
    .A3(_07727_),
    .ZN(_09790_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18683_ (.A1(_09764_),
    .A2(_09790_),
    .ZN(_09791_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18684_ (.I(_15653_[0]),
    .ZN(_09792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18685_ (.A1(_09792_),
    .A2(net20697),
    .ZN(_09793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18686_ (.A1(net20810),
    .A2(_15646_[0]),
    .ZN(_09794_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17582 (.I(_11370_),
    .Z(net17582));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18688_ (.A1(net534),
    .A2(_09794_),
    .A3(net20685),
    .ZN(_09796_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17580 (.I(_11420_),
    .Z(net17580));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18690_ (.A1(_09768_),
    .A2(net20461),
    .ZN(_09798_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18691_ (.A1(_09796_),
    .A2(net20672),
    .A3(_09798_),
    .ZN(_09799_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18692_ (.I(_09783_),
    .ZN(_09800_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18693_ (.I(_15646_[0]),
    .ZN(_09801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18694_ (.A1(net20810),
    .A2(_09801_),
    .ZN(_09802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18695_ (.I(_09802_),
    .ZN(_09803_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18696_ (.A1(_09800_),
    .A2(_09803_),
    .B(net20463),
    .ZN(_09804_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18697_ (.A1(_09768_),
    .A2(net20688),
    .B(net20669),
    .ZN(_09805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18698_ (.A1(_09804_),
    .A2(_09805_),
    .ZN(_09806_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17579 (.I(_11455_),
    .Z(net17579));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18700_ (.A1(_09799_),
    .A2(_09806_),
    .A3(_07727_),
    .ZN(_09808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18701_ (.A1(net20810),
    .A2(_09765_),
    .ZN(_09809_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17578 (.I(_11458_),
    .Z(net17578));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18703_ (.A1(_09809_),
    .A2(net20461),
    .B(net20669),
    .ZN(_09811_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18704_ (.A1(_09739_),
    .A2(_09811_),
    .ZN(_09812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18705_ (.A1(net20697),
    .A2(net20472),
    .ZN(_09813_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18706_ (.A1(net20289),
    .A2(net20461),
    .Z(_09814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18707_ (.A1(_09814_),
    .A2(net20078),
    .ZN(_09815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18708_ (.A1(_09812_),
    .A2(_09815_),
    .ZN(_09816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18709_ (.I(_09779_),
    .ZN(_09817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18710_ (.A1(_09817_),
    .A2(net20461),
    .ZN(_09818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18711_ (.A1(net20685),
    .A2(_15662_[0]),
    .B(net20669),
    .ZN(_09819_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18712_ (.A1(_09818_),
    .A2(_09819_),
    .B(_07727_),
    .ZN(_09820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18713_ (.A1(_09816_),
    .A2(_09820_),
    .ZN(_09821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18714_ (.A1(_09808_),
    .A2(_09821_),
    .ZN(_09822_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17577 (.I(_11462_),
    .Z(net17577));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18716_ (.A1(_09822_),
    .A2(_09762_),
    .ZN(_09824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18717_ (.A1(_09791_),
    .A2(_09824_),
    .ZN(_09825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18718_ (.A1(_09825_),
    .A2(_00399_),
    .ZN(_09826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18719_ (.A1(net20697),
    .A2(net20705),
    .ZN(_09827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18720_ (.A1(_09827_),
    .A2(net20465),
    .Z(_09828_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17581 (.I(_11395_),
    .Z(net17581));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18722_ (.A1(_09828_),
    .A2(_07717_),
    .ZN(_09830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18723_ (.A1(net20698),
    .A2(_15646_[0]),
    .ZN(_09831_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17575 (.I(_11473_),
    .Z(net17575));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18725_ (.A1(net20074),
    .A2(net19886),
    .A3(net20693),
    .ZN(_09833_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17574 (.I(_11481_),
    .Z(net17574));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18727_ (.A1(_09830_),
    .A2(_09833_),
    .B(net20668),
    .ZN(_09835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18728_ (.A1(_09831_),
    .A2(net20465),
    .ZN(_09836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18729_ (.I(_09836_),
    .ZN(_09837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18730_ (.A1(net20810),
    .A2(net666),
    .ZN(_09838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18731_ (.A1(_09837_),
    .A2(_09838_),
    .ZN(_09839_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _18732_ (.I(_09753_),
    .ZN(_09840_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18733_ (.I(_15643_[0]),
    .ZN(_09841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18734_ (.A1(net20700),
    .A2(_09841_),
    .ZN(_09842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18735_ (.A1(net18945),
    .A2(net19879),
    .ZN(_09843_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17583 (.I(_11369_),
    .Z(net17583));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18737_ (.A1(_09839_),
    .A2(_09843_),
    .A3(net20576),
    .ZN(_09845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18738_ (.A1(_09835_),
    .A2(_09845_),
    .B(_09762_),
    .ZN(_09846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18739_ (.A1(net20810),
    .A2(net20704),
    .ZN(_09847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18740_ (.A1(_09837_),
    .A2(net20450),
    .ZN(_09848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18741_ (.A1(_09841_),
    .A2(net20810),
    .ZN(_09849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18742_ (.A1(_09849_),
    .A2(net20685),
    .ZN(_09850_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18743_ (.I(_09850_),
    .ZN(_09851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18744_ (.A1(net18944),
    .A2(net20454),
    .ZN(_09852_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18745_ (.A1(_09848_),
    .A2(_09852_),
    .A3(net20576),
    .ZN(_09853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18746_ (.A1(net20697),
    .A2(net20704),
    .ZN(_09854_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18747_ (.I(_09854_),
    .ZN(_09855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18748_ (.A1(_09855_),
    .A2(net20461),
    .ZN(_09856_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18749_ (.A1(_09856_),
    .A2(_09798_),
    .Z(_09857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18750_ (.A1(net18948),
    .A2(_09857_),
    .ZN(_09858_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17576 (.I(_11468_),
    .Z(net17576));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18752_ (.A1(_09853_),
    .A2(_09858_),
    .A3(net20668),
    .ZN(_09860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18753_ (.A1(_09846_),
    .A2(_09860_),
    .B(_00399_),
    .ZN(_09861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18754_ (.A1(_09856_),
    .A2(_07717_),
    .ZN(_09862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18755_ (.A1(net20697),
    .A2(net20087),
    .ZN(_09863_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18756_ (.A1(_09863_),
    .A2(net20696),
    .Z(_09864_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18757_ (.A1(net19889),
    .A2(net20696),
    .ZN(_09865_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18758_ (.A1(_09862_),
    .A2(_09864_),
    .A3(net19435),
    .ZN(_09866_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _18759_ (.I(_09809_),
    .ZN(_09867_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17586 (.I(_11293_),
    .Z(net17586));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18761_ (.A1(_09800_),
    .A2(_09867_),
    .B(net20462),
    .ZN(_09869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18762_ (.A1(net20697),
    .A2(net20368),
    .ZN(_09870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18763_ (.A1(net18945),
    .A2(net20286),
    .ZN(_09871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18764_ (.A1(_09871_),
    .A2(_09869_),
    .B(net20575),
    .ZN(_09872_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18765_ (.A1(_09872_),
    .A2(_09866_),
    .B(net20668),
    .ZN(_09873_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18766_ (.A1(_09784_),
    .A2(net20461),
    .Z(_09874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18767_ (.A1(net20705),
    .A2(net20704),
    .ZN(_09875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18768_ (.A1(_09874_),
    .A2(net20447),
    .ZN(_09876_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18769_ (.I(_09784_),
    .ZN(_09877_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18770_ (.I(_09875_),
    .ZN(_09878_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17591 (.I(_10906_),
    .Z(net17591));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _18772_ (.A1(_09877_),
    .A2(_09878_),
    .B(net20685),
    .ZN(_09880_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18773_ (.A1(_09876_),
    .A2(net19876),
    .A3(net20575),
    .ZN(_09881_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18774_ (.A1(_09767_),
    .A2(net20688),
    .B(_07717_),
    .ZN(_09882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18775_ (.A1(net20460),
    .A2(net19888),
    .ZN(_09883_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _18776_ (.I(_09883_),
    .ZN(_09884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18777_ (.A1(net20700),
    .A2(net20157),
    .ZN(_09885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18778_ (.A1(net662),
    .A2(net20072),
    .ZN(_09886_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18779_ (.A1(net20810),
    .A2(_09782_),
    .Z(_09887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18780_ (.A1(_09887_),
    .A2(net20687),
    .ZN(_09888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18781_ (.A1(_09882_),
    .A2(_09886_),
    .A3(net19433),
    .ZN(_09889_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18782_ (.A1(_09881_),
    .A2(_09889_),
    .A3(net20557),
    .ZN(_09890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18783_ (.A1(_09762_),
    .A2(_09890_),
    .A3(_09873_),
    .ZN(_09891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18784_ (.A1(_09861_),
    .A2(_09891_),
    .ZN(_09892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18785_ (.A1(_09826_),
    .A2(_09892_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18786_ (.A1(_09774_),
    .A2(_09855_),
    .Z(_09893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18787_ (.A1(_09874_),
    .A2(net20286),
    .ZN(_09894_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17567 (.I(_11638_),
    .Z(net17567));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18789_ (.A1(_09893_),
    .A2(_09894_),
    .A3(net20670),
    .ZN(_09896_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18790_ (.A1(net20076),
    .A2(net20463),
    .B(_07717_),
    .ZN(_09897_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18791_ (.I(_09798_),
    .ZN(_09898_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18792_ (.A1(_09897_),
    .A2(_09898_),
    .ZN(_09899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18793_ (.I(_09813_),
    .ZN(_09900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18794_ (.A1(_09900_),
    .A2(net20461),
    .ZN(_09901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18795_ (.A1(_09817_),
    .A2(net20685),
    .ZN(_09902_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18796_ (.A1(_09901_),
    .A2(_09902_),
    .Z(_09903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18797_ (.A1(_09899_),
    .A2(_09903_),
    .ZN(_09904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18798_ (.A1(_09896_),
    .A2(_09904_),
    .A3(net20557),
    .ZN(_09905_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18799_ (.A1(_09741_),
    .A2(net20685),
    .Z(_09906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18800_ (.A1(_09906_),
    .A2(_09901_),
    .Z(_09907_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17568 (.I(_11544_),
    .Z(net17568));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18802_ (.A1(net19437),
    .A2(net20676),
    .Z(_09909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18803_ (.A1(_09909_),
    .A2(_09907_),
    .B(net20561),
    .ZN(_09910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18804_ (.A1(_09885_),
    .A2(net20685),
    .Z(_09911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18805_ (.A1(net20810),
    .A2(net20156),
    .ZN(_09912_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18806_ (.A1(_09911_),
    .A2(net20070),
    .ZN(_09913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18807_ (.A1(_09849_),
    .A2(net20465),
    .ZN(_09914_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18808_ (.I(_09914_),
    .ZN(_09915_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18809_ (.I(_15657_[0]),
    .ZN(_09916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18810_ (.A1(net20698),
    .A2(_09916_),
    .ZN(_09917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18811_ (.A1(_09915_),
    .A2(_09917_),
    .ZN(_09918_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18812_ (.A1(_09913_),
    .A2(_09918_),
    .A3(net20567),
    .ZN(_09919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18813_ (.A1(_09919_),
    .A2(_09910_),
    .ZN(_09920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18814_ (.A1(_09905_),
    .A2(net20839),
    .A3(_09920_),
    .ZN(_09921_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18815_ (.A1(_09870_),
    .A2(_09838_),
    .A3(net20459),
    .ZN(_09922_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18816_ (.A1(net20810),
    .A2(net20157),
    .ZN(_09923_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17572 (.I(_11494_),
    .Z(net17572));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18818_ (.A1(net20074),
    .A2(net20069),
    .A3(net20693),
    .ZN(_09925_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18819_ (.A1(_09922_),
    .A2(_09925_),
    .A3(net20558),
    .ZN(_09926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18820_ (.A1(_09926_),
    .A2(net20576),
    .ZN(_09927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18821_ (.A1(net20697),
    .A2(net20474),
    .ZN(_09928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18822_ (.A1(_09874_),
    .A2(_09928_),
    .ZN(_09929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18823_ (.A1(_09893_),
    .A2(_09929_),
    .ZN(_09930_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18824_ (.A1(_09930_),
    .A2(_07727_),
    .ZN(_09931_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18825_ (.A1(net20455),
    .A2(_15669_[0]),
    .A3(_07727_),
    .Z(_09932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18826_ (.A1(_09783_),
    .A2(_09741_),
    .ZN(_09933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18827_ (.A1(_09933_),
    .A2(net20465),
    .ZN(_09934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18828_ (.A1(_09932_),
    .A2(net18943),
    .ZN(_09935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18829_ (.A1(_09935_),
    .A2(net20677),
    .ZN(_09936_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18830_ (.A1(_09927_),
    .A2(_09931_),
    .B(net20646),
    .C(_09936_),
    .ZN(_09937_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17573 (.I(_11491_),
    .Z(net17573));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18832_ (.A1(_07744_),
    .A2(_09937_),
    .A3(_09921_),
    .ZN(_09939_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17616 (.I(_07015_),
    .Z(net17616));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18834_ (.A1(_09758_),
    .A2(net20465),
    .B(net20669),
    .ZN(_09941_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _18835_ (.I(_09847_),
    .ZN(_09942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18836_ (.A1(net20842),
    .A2(net21514),
    .B(_15665_[0]),
    .ZN(_09943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18837_ (.A1(_09942_),
    .A2(net20457),
    .B(_09943_),
    .ZN(_09944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18838_ (.A1(_09941_),
    .A2(_09944_),
    .B(net20558),
    .ZN(_09945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18839_ (.A1(_09851_),
    .A2(_09863_),
    .ZN(_09946_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17589 (.I(_11247_),
    .Z(net17589));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18841_ (.A1(net20086),
    .A2(_09802_),
    .ZN(_09948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18842_ (.A1(_09948_),
    .A2(net20466),
    .ZN(_09949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18843_ (.A1(_09946_),
    .A2(net20677),
    .A3(_09949_),
    .ZN(_09950_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17564 (.I(_12054_),
    .Z(net17564));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18845_ (.A1(_09945_),
    .A2(_09950_),
    .B(net20839),
    .ZN(_09952_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18846_ (.A1(_09772_),
    .A2(net20461),
    .ZN(_09953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18847_ (.I(_09953_),
    .ZN(_09954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18848_ (.A1(_09954_),
    .A2(net20288),
    .ZN(_09955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18849_ (.A1(net18946),
    .A2(net20454),
    .ZN(_09956_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18850_ (.A1(_09955_),
    .A2(_09956_),
    .A3(net20575),
    .ZN(_09957_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18851_ (.A1(_09778_),
    .A2(net20459),
    .A3(net20447),
    .ZN(_09958_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18852_ (.A1(net20698),
    .A2(_09801_),
    .Z(_09959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18853_ (.A1(_09959_),
    .A2(net20690),
    .ZN(_09960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18854_ (.A1(_09958_),
    .A2(_09960_),
    .A3(net20673),
    .ZN(_09961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18855_ (.A1(_09957_),
    .A2(net20559),
    .A3(_09961_),
    .ZN(_09962_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18856_ (.A1(_09962_),
    .A2(_09952_),
    .B(_07744_),
    .ZN(_09963_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18857_ (.A1(net20082),
    .A2(_09838_),
    .A3(net20461),
    .Z(_09964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18858_ (.A1(net20474),
    .A2(net20472),
    .ZN(_09965_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18859_ (.A1(net20283),
    .A2(_09838_),
    .B(net20461),
    .ZN(_09966_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18860_ (.A1(_09964_),
    .A2(_09966_),
    .B(net20676),
    .ZN(_09967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18861_ (.A1(_09814_),
    .A2(net20076),
    .ZN(_09968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18862_ (.A1(_09840_),
    .A2(net20085),
    .ZN(_09969_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18863_ (.A1(_09968_),
    .A2(_09969_),
    .A3(net20564),
    .ZN(_09970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18864_ (.A1(_09967_),
    .A2(_09970_),
    .ZN(_09971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18865_ (.A1(_09971_),
    .A2(net20668),
    .ZN(_09972_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18866_ (.A1(_09842_),
    .A2(net20691),
    .Z(_09973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18867_ (.A1(_09973_),
    .A2(net20451),
    .ZN(_09974_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18868_ (.A1(_09974_),
    .A2(net20564),
    .A3(_09906_),
    .ZN(_09975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18869_ (.A1(net20465),
    .A2(net20154),
    .ZN(_09976_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18870_ (.A1(_09976_),
    .A2(net20697),
    .Z(_09977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18871_ (.A1(_09913_),
    .A2(net20675),
    .A3(_09977_),
    .ZN(_09978_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18872_ (.A1(_09975_),
    .A2(_09978_),
    .A3(net20560),
    .ZN(_09979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18873_ (.A1(net20840),
    .A2(_09979_),
    .A3(_09972_),
    .ZN(_09980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18874_ (.A1(_09963_),
    .A2(_09980_),
    .ZN(_09981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18875_ (.A1(_09981_),
    .A2(_09939_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18876_ (.A1(_09757_),
    .A2(_09802_),
    .A3(net20685),
    .ZN(_09982_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18877_ (.A1(_09780_),
    .A2(_09982_),
    .A3(net20678),
    .Z(_09983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18878_ (.A1(_09778_),
    .A2(_09831_),
    .A3(net20681),
    .ZN(_09984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18879_ (.A1(_09842_),
    .A2(net19886),
    .A3(net20465),
    .ZN(_09985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18880_ (.A1(_09984_),
    .A2(_09985_),
    .B(net20678),
    .ZN(_09986_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18881_ (.A1(_09983_),
    .A2(_09986_),
    .B(net20648),
    .ZN(_09987_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17561 (.I(_12216_),
    .Z(net17561));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18883_ (.A1(_09747_),
    .A2(net20465),
    .B(net20675),
    .ZN(_09989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18884_ (.A1(net20702),
    .A2(net20084),
    .ZN(_09990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18885_ (.A1(_09990_),
    .A2(_09838_),
    .A3(net20694),
    .ZN(_09991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18886_ (.A1(net20700),
    .A2(net20155),
    .ZN(_09992_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18887_ (.A1(_09992_),
    .A2(net20694),
    .Z(_09993_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18888_ (.A1(_09989_),
    .A2(_09991_),
    .A3(_09993_),
    .ZN(_09994_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18889_ (.A1(_09746_),
    .A2(net20683),
    .B(net20680),
    .ZN(_09995_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18890_ (.I(_09995_),
    .ZN(_09996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18891_ (.A1(_09990_),
    .A2(net20451),
    .A3(net20685),
    .ZN(_09997_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18892_ (.A1(_09996_),
    .A2(_09760_),
    .A3(_09997_),
    .ZN(_09998_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18893_ (.A1(_09994_),
    .A2(_09998_),
    .A3(net20839),
    .ZN(_09999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18894_ (.A1(_09987_),
    .A2(_09999_),
    .A3(net20668),
    .ZN(_10000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18895_ (.A1(_09992_),
    .A2(net20465),
    .ZN(_10001_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18896_ (.A1(_10001_),
    .A2(net20073),
    .B(net20568),
    .ZN(_10002_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18897_ (.A1(net20448),
    .A2(_09746_),
    .A3(net20690),
    .Z(_10003_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18898_ (.A1(_10002_),
    .A2(_10003_),
    .ZN(_10004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18899_ (.A1(net19884),
    .A2(_09838_),
    .A3(net20466),
    .ZN(_10005_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18900_ (.A1(net20083),
    .A2(net19887),
    .A3(net20686),
    .ZN(_10006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18901_ (.A1(_10005_),
    .A2(_10006_),
    .B(net20570),
    .ZN(_10007_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18902_ (.A1(_10004_),
    .A2(_10007_),
    .B(net20839),
    .ZN(_10008_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18903_ (.A1(_09836_),
    .A2(net20678),
    .Z(_10009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18904_ (.A1(_09911_),
    .A2(_09849_),
    .ZN(_10010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18905_ (.A1(_10009_),
    .A2(_10010_),
    .B(net20837),
    .ZN(_10011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18906_ (.A1(net20697),
    .A2(net20367),
    .ZN(_10012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18907_ (.I(_10012_),
    .ZN(_10013_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18908_ (.A1(_10013_),
    .A2(net20073),
    .B(net20686),
    .ZN(_10014_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18909_ (.A1(net20284),
    .A2(net20466),
    .A3(net19887),
    .ZN(_10015_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18910_ (.A1(_10014_),
    .A2(net20570),
    .A3(_10015_),
    .ZN(_10016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18911_ (.A1(_10011_),
    .A2(_10016_),
    .ZN(_10017_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18912_ (.A1(_10008_),
    .A2(net20562),
    .A3(_10017_),
    .ZN(_10018_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18913_ (.A1(_10000_),
    .A2(_10018_),
    .A3(_07744_),
    .ZN(_10019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18914_ (.A1(_09867_),
    .A2(net20468),
    .B(_07717_),
    .ZN(_10020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18915_ (.A1(_09840_),
    .A2(_09990_),
    .ZN(_10021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18916_ (.A1(_10020_),
    .A2(_10021_),
    .B(net20668),
    .ZN(_10022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18917_ (.A1(_09784_),
    .A2(net20685),
    .Z(_10023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18918_ (.A1(_10023_),
    .A2(_09885_),
    .ZN(_10024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18919_ (.A1(_10024_),
    .A2(_07717_),
    .A3(_09934_),
    .ZN(_10025_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18920_ (.A1(_10022_),
    .A2(_10025_),
    .ZN(_10026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18921_ (.A1(net20455),
    .A2(_15667_[0]),
    .ZN(_10027_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18922_ (.A1(_10027_),
    .A2(_07717_),
    .ZN(_10028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18923_ (.I(_10028_),
    .ZN(_10029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18924_ (.A1(_10029_),
    .A2(_09984_),
    .ZN(_10030_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18925_ (.A1(net20455),
    .A2(_15660_[0]),
    .Z(_10031_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18926_ (.A1(_10031_),
    .A2(net19881),
    .A3(net20678),
    .ZN(_10032_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18927_ (.A1(_10030_),
    .A2(_10032_),
    .A3(net20668),
    .ZN(_10033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18928_ (.A1(_10026_),
    .A2(net20646),
    .A3(_10033_),
    .ZN(_10034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18929_ (.A1(_10034_),
    .A2(_00399_),
    .ZN(_10035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18930_ (.I(_10035_),
    .ZN(_10036_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18931_ (.A1(net19882),
    .A2(_09887_),
    .B(net20687),
    .ZN(_10037_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18932_ (.A1(net20286),
    .A2(net20450),
    .A3(net20459),
    .ZN(_10038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18933_ (.A1(_10037_),
    .A2(_10038_),
    .B(net20677),
    .ZN(_10039_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18934_ (.A1(_09778_),
    .A2(net20685),
    .A3(net20446),
    .ZN(_10040_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18935_ (.A1(net20681),
    .A2(_15669_[0]),
    .Z(_10041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18936_ (.A1(net20067),
    .A2(_10041_),
    .B(net20576),
    .ZN(_10042_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18937_ (.A1(_10039_),
    .A2(_10042_),
    .B(net20668),
    .ZN(_10043_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18938_ (.A1(net20448),
    .A2(net20452),
    .A3(net20681),
    .ZN(_10044_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18939_ (.A1(_09780_),
    .A2(_10044_),
    .A3(net20572),
    .ZN(_10045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18940_ (.A1(_09794_),
    .A2(net20685),
    .ZN(_10046_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _18941_ (.I(_09863_),
    .ZN(_10047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18942_ (.A1(net20465),
    .A2(_15662_[0]),
    .ZN(_10048_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18943_ (.A1(net19874),
    .A2(_10047_),
    .B(_10048_),
    .C(net20679),
    .ZN(_10049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18944_ (.A1(_10045_),
    .A2(_10049_),
    .A3(net20562),
    .ZN(_10050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18945_ (.A1(_10043_),
    .A2(net20838),
    .A3(_10050_),
    .ZN(_10051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18946_ (.A1(_10036_),
    .A2(_10051_),
    .ZN(_10052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18947_ (.A1(_10019_),
    .A2(_10052_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18948_ (.A1(_09851_),
    .A2(_09990_),
    .Z(_10053_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18949_ (.A1(net20448),
    .A2(net20070),
    .A3(net20461),
    .Z(_10054_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18950_ (.A1(_10053_),
    .A2(_10054_),
    .B(net20676),
    .ZN(_10055_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18951_ (.I(_09887_),
    .ZN(_10056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18952_ (.A1(_09814_),
    .A2(_10056_),
    .ZN(_10057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18953_ (.A1(_09864_),
    .A2(net20076),
    .ZN(_10058_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18954_ (.A1(_10057_),
    .A2(_10058_),
    .A3(_07717_),
    .ZN(_10059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18955_ (.A1(_10055_),
    .A2(_10059_),
    .A3(_09762_),
    .ZN(_10060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18956_ (.A1(_09923_),
    .A2(net20461),
    .ZN(_10061_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18957_ (.I(_10061_),
    .ZN(_10062_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18958_ (.A1(_10062_),
    .A2(_09863_),
    .Z(_10063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18959_ (.A1(_09960_),
    .A2(_09888_),
    .ZN(_10064_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18960_ (.A1(_10063_),
    .A2(_10064_),
    .B(net20672),
    .ZN(_10065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18961_ (.A1(net19885),
    .A2(_09884_),
    .ZN(_10066_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18962_ (.A1(_09880_),
    .A2(_10066_),
    .A3(_07717_),
    .ZN(_10067_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18963_ (.A1(_10065_),
    .A2(net20837),
    .A3(_10067_),
    .ZN(_10068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18964_ (.A1(_10060_),
    .A2(_10068_),
    .ZN(_10069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18965_ (.A1(_10069_),
    .A2(net20561),
    .ZN(_10070_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18966_ (.A1(net20071),
    .A2(net20285),
    .B(net20461),
    .ZN(_10071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18967_ (.A1(net18946),
    .A2(net20448),
    .ZN(_10072_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18968_ (.A1(_10071_),
    .A2(_10072_),
    .A3(net20674),
    .ZN(_10073_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18969_ (.A1(_09863_),
    .A2(net20691),
    .B(net20676),
    .ZN(_10074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18970_ (.A1(net20448),
    .A2(net20453),
    .A3(net20464),
    .ZN(_10075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18971_ (.A1(_10074_),
    .A2(_10075_),
    .B(net20837),
    .ZN(_10076_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18972_ (.A1(_10073_),
    .A2(_10076_),
    .B(net20561),
    .ZN(_10077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18973_ (.A1(_09793_),
    .A2(net20465),
    .Z(_10078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18974_ (.A1(_10078_),
    .A2(net20070),
    .ZN(_10079_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18975_ (.A1(_09974_),
    .A2(_10079_),
    .A3(net20565),
    .ZN(_10080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18976_ (.A1(_09831_),
    .A2(net20681),
    .ZN(_10081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18977_ (.A1(_10071_),
    .A2(net20674),
    .A3(net19873),
    .ZN(_10082_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18978_ (.A1(_10080_),
    .A2(_10082_),
    .A3(net20840),
    .ZN(_10083_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18979_ (.A1(_10077_),
    .A2(_10083_),
    .B(_07744_),
    .ZN(_10084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18980_ (.A1(_10070_),
    .A2(_10084_),
    .ZN(_10085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18981_ (.A1(_09793_),
    .A2(_09784_),
    .A3(net20690),
    .ZN(_10086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18982_ (.A1(net18943),
    .A2(_10086_),
    .B(net20570),
    .ZN(_10087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18983_ (.I(_10002_),
    .ZN(_10088_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18984_ (.A1(_10087_),
    .A2(_10088_),
    .B(net20668),
    .ZN(_10089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18985_ (.A1(_09812_),
    .A2(_09958_),
    .ZN(_10090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18986_ (.A1(net662),
    .A2(net19879),
    .ZN(_10091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18987_ (.A1(_09827_),
    .A2(_09746_),
    .ZN(_10092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18988_ (.A1(_10092_),
    .A2(net20689),
    .ZN(_10093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18989_ (.A1(_10091_),
    .A2(_10093_),
    .A3(net20575),
    .ZN(_10094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18990_ (.A1(_10090_),
    .A2(_10094_),
    .A3(net20559),
    .ZN(_10095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18991_ (.A1(_10089_),
    .A2(_10095_),
    .A3(net20839),
    .ZN(_10096_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18992_ (.A1(net19879),
    .A2(net20290),
    .A3(net20690),
    .ZN(_10097_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18993_ (.A1(_09827_),
    .A2(net20466),
    .A3(net659),
    .ZN(_10098_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18994_ (.A1(_10097_),
    .A2(_10098_),
    .A3(net20668),
    .ZN(_10099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18995_ (.A1(_09747_),
    .A2(net20693),
    .ZN(_10100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18996_ (.A1(_10005_),
    .A2(net20560),
    .A3(_10100_),
    .ZN(_10101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18997_ (.A1(_10099_),
    .A2(_10101_),
    .B(net20569),
    .ZN(_10102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18998_ (.A1(net20699),
    .A2(net20153),
    .ZN(_10103_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18999_ (.A1(net20292),
    .A2(_10103_),
    .A3(net20467),
    .ZN(_10104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19000_ (.A1(_10047_),
    .A2(net20695),
    .ZN(_10105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19001_ (.A1(_10104_),
    .A2(_10105_),
    .ZN(_10106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19002_ (.A1(_09865_),
    .A2(_07727_),
    .ZN(_10107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19003_ (.A1(_09805_),
    .A2(_10107_),
    .ZN(_10108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19004_ (.A1(net20668),
    .A2(_10106_),
    .B(_10108_),
    .ZN(_10109_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19005_ (.A1(_10102_),
    .A2(_10109_),
    .B(_09762_),
    .ZN(_10110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19006_ (.A1(_10096_),
    .A2(_10110_),
    .A3(_07744_),
    .ZN(_10111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19007_ (.A1(_10111_),
    .A2(_10085_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19008_ (.A1(net20696),
    .A2(net20076),
    .B(_09893_),
    .ZN(_10112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19009_ (.A1(_09874_),
    .A2(net19879),
    .ZN(_10113_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19010_ (.A1(net20470),
    .A2(net20670),
    .Z(_10114_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19011_ (.A1(_10113_),
    .A2(_10114_),
    .B(_07727_),
    .ZN(_10115_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19012_ (.A1(_10112_),
    .A2(net19878),
    .B(_10115_),
    .ZN(_10116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19013_ (.A1(_09954_),
    .A2(net20083),
    .ZN(_10117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19014_ (.A1(net18948),
    .A2(_10117_),
    .ZN(_10118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19015_ (.A1(net20072),
    .A2(net20681),
    .B(net20678),
    .ZN(_10119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19016_ (.A1(_09917_),
    .A2(net20455),
    .ZN(_10120_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19017_ (.A1(_10119_),
    .A2(net19872),
    .B(net20668),
    .ZN(_10121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19018_ (.A1(_10118_),
    .A2(_10121_),
    .B(_09762_),
    .ZN(_10122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19019_ (.A1(_10116_),
    .A2(_10122_),
    .ZN(_10123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19020_ (.A1(_09793_),
    .A2(net20681),
    .ZN(_10124_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19021_ (.A1(_10124_),
    .A2(_09942_),
    .Z(_10125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19022_ (.A1(_09803_),
    .A2(net20461),
    .ZN(_10126_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19023_ (.A1(_10125_),
    .A2(_07717_),
    .A3(_10126_),
    .ZN(_10127_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19024_ (.A1(net20682),
    .A2(net20157),
    .B(net20678),
    .ZN(_10128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19025_ (.I(_10128_),
    .ZN(_10129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19026_ (.A1(net20081),
    .A2(net20682),
    .ZN(_10130_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19027_ (.A1(_10129_),
    .A2(_10130_),
    .B(net20668),
    .ZN(_10131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19028_ (.A1(_10127_),
    .A2(_10131_),
    .B(net20841),
    .ZN(_10132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19029_ (.A1(_09770_),
    .A2(net19875),
    .A3(net20671),
    .ZN(_10133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19030_ (.A1(_09965_),
    .A2(_09847_),
    .ZN(_10134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19031_ (.A1(_10134_),
    .A2(net20465),
    .ZN(_10135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19032_ (.A1(net19871),
    .A2(_10086_),
    .A3(net20570),
    .ZN(_10136_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19033_ (.A1(_10133_),
    .A2(_10136_),
    .A3(net20668),
    .ZN(_10137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19034_ (.A1(_10132_),
    .A2(_10137_),
    .ZN(_10138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19035_ (.A1(_10123_),
    .A2(_10138_),
    .B(_00399_),
    .ZN(_10139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19036_ (.A1(_09929_),
    .A2(_10040_),
    .ZN(_10140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19037_ (.A1(_10140_),
    .A2(net20668),
    .ZN(_10141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19038_ (.A1(_09928_),
    .A2(_09838_),
    .A3(net20685),
    .ZN(_10142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19039_ (.A1(_10142_),
    .A2(_09922_),
    .ZN(_10143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19040_ (.A1(_10143_),
    .A2(_07727_),
    .ZN(_10144_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19041_ (.A1(_10141_),
    .A2(net20677),
    .A3(_10144_),
    .ZN(_10145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19042_ (.I(_09768_),
    .ZN(_10146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19043_ (.A1(_10124_),
    .A2(_10146_),
    .ZN(_10147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19044_ (.A1(_10147_),
    .A2(net20562),
    .B(net20679),
    .ZN(_10148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19045_ (.A1(_09778_),
    .A2(_09766_),
    .A3(net20681),
    .ZN(_10149_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19046_ (.A1(_10135_),
    .A2(_10149_),
    .A3(net20668),
    .ZN(_10150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19047_ (.A1(_10148_),
    .A2(_10150_),
    .B(_09762_),
    .ZN(_10151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19048_ (.A1(_10145_),
    .A2(_10151_),
    .ZN(_10152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19049_ (.A1(_10152_),
    .A2(_00399_),
    .ZN(_10153_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19050_ (.I(_10046_),
    .ZN(_10154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19051_ (.A1(_10154_),
    .A2(net20448),
    .ZN(_10155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19052_ (.A1(_10155_),
    .A2(net20571),
    .A3(_09985_),
    .ZN(_10156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19053_ (.I(net19883),
    .ZN(_10157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19054_ (.A1(net20294),
    .A2(net20474),
    .ZN(_10158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19055_ (.A1(_10157_),
    .A2(_09949_),
    .A3(_10158_),
    .ZN(_10159_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19056_ (.A1(_10156_),
    .A2(_10159_),
    .A3(net20668),
    .ZN(_10160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19057_ (.A1(net683),
    .A2(_09863_),
    .ZN(_10161_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19058_ (.A1(_10161_),
    .A2(net20674),
    .A3(_09796_),
    .ZN(_10162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19059_ (.A1(_09902_),
    .A2(_07717_),
    .Z(_10163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19060_ (.A1(_09760_),
    .A2(_09746_),
    .Z(_10164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19061_ (.A1(_10163_),
    .A2(_10164_),
    .ZN(_10165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19062_ (.A1(_10162_),
    .A2(_10165_),
    .A3(net20560),
    .ZN(_10166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19063_ (.A1(_10166_),
    .A2(_10160_),
    .B(net20839),
    .ZN(_10167_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19064_ (.A1(_10167_),
    .A2(_10153_),
    .ZN(_10168_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19065_ (.A1(_10139_),
    .A2(_10168_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19066_ (.A1(_09840_),
    .A2(_09831_),
    .Z(_10169_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19067_ (.A1(_09793_),
    .A2(_09847_),
    .A3(net20465),
    .Z(_10170_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19068_ (.A1(_10169_),
    .A2(_10170_),
    .A3(net20675),
    .Z(_10171_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19069_ (.A1(net20690),
    .A2(net664),
    .B(_07717_),
    .ZN(_10172_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19070_ (.A1(_09876_),
    .A2(_10172_),
    .B(_09762_),
    .ZN(_10173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19071_ (.A1(_10171_),
    .A2(_10173_),
    .ZN(_10174_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19072_ (.A1(net20074),
    .A2(net20069),
    .A3(net20465),
    .ZN(_10175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19073_ (.I(_10023_),
    .ZN(_10176_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19074_ (.A1(_10175_),
    .A2(_10176_),
    .A3(net20675),
    .ZN(_10177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19075_ (.I(_09973_),
    .ZN(_10178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19076_ (.A1(_09941_),
    .A2(_10178_),
    .ZN(_10179_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19077_ (.A1(_10177_),
    .A2(_10179_),
    .A3(net20647),
    .ZN(_10180_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19078_ (.A1(_10174_),
    .A2(net20560),
    .A3(_10180_),
    .ZN(_10181_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19079_ (.A1(_09990_),
    .A2(_09838_),
    .A3(net20461),
    .Z(_10182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19080_ (.A1(_09800_),
    .A2(net20692),
    .B(net20676),
    .ZN(_10183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19081_ (.A1(_10062_),
    .A2(net19880),
    .ZN(_10184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19082_ (.A1(_10183_),
    .A2(_10184_),
    .ZN(_10185_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _19083_ (.A1(_09745_),
    .A2(_10182_),
    .B(_10185_),
    .C(net20840),
    .ZN(_10186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19084_ (.A1(net20692),
    .A2(net20080),
    .ZN(_10187_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19085_ (.A1(_10061_),
    .A2(net20676),
    .A3(_10187_),
    .Z(_10188_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19086_ (.A1(_10188_),
    .A2(net20840),
    .ZN(_10189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19087_ (.A1(net18947),
    .A2(_10103_),
    .ZN(_10190_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19088_ (.A1(net19880),
    .A2(net20070),
    .A3(net20461),
    .ZN(_10191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19089_ (.A1(_10190_),
    .A2(_10191_),
    .A3(net20564),
    .ZN(_10192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19090_ (.A1(_10189_),
    .A2(_10192_),
    .B(net20560),
    .ZN(_10193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19091_ (.A1(_10186_),
    .A2(_10193_),
    .ZN(_10194_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19092_ (.A1(_10181_),
    .A2(_10194_),
    .A3(_07744_),
    .ZN(_10195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19093_ (.A1(_10001_),
    .A2(net19437),
    .ZN(_10196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19094_ (.A1(_09882_),
    .A2(_10196_),
    .B(net20837),
    .ZN(_10197_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19095_ (.A1(net20292),
    .A2(_09917_),
    .A3(net20467),
    .ZN(_10198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19096_ (.A1(_10163_),
    .A2(_10198_),
    .ZN(_10199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19097_ (.A1(_10197_),
    .A2(_10199_),
    .B(net20560),
    .ZN(_10200_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19098_ (.A1(_09954_),
    .A2(net20673),
    .A3(_09959_),
    .Z(_10201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19099_ (.A1(_10093_),
    .A2(net20669),
    .A3(net19434),
    .ZN(_10202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19100_ (.A1(_10201_),
    .A2(_10202_),
    .A3(net20837),
    .ZN(_10203_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19101_ (.A1(_10200_),
    .A2(_10203_),
    .B(_07744_),
    .ZN(_10204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19102_ (.A1(net20695),
    .A2(net20704),
    .ZN(_10205_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19103_ (.A1(_10135_),
    .A2(net20669),
    .A3(_10205_),
    .Z(_10206_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19104_ (.A1(_09933_),
    .A2(net20465),
    .B(_07717_),
    .ZN(_10207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19105_ (.A1(_09828_),
    .A2(net20283),
    .Z(_10208_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19106_ (.A1(_10207_),
    .A2(_10208_),
    .ZN(_10209_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19107_ (.A1(_10206_),
    .A2(_10209_),
    .B(net20647),
    .ZN(_10210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19108_ (.A1(_09973_),
    .A2(net19886),
    .ZN(_10211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19109_ (.A1(_09857_),
    .A2(net20674),
    .A3(_10211_),
    .ZN(_10212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19110_ (.A1(_10078_),
    .A2(net20078),
    .ZN(_10213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19111_ (.A1(_10023_),
    .A2(_09990_),
    .ZN(_10214_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19112_ (.A1(_10213_),
    .A2(_10214_),
    .A3(net20565),
    .ZN(_10215_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19113_ (.A1(_10212_),
    .A2(_10215_),
    .A3(net20840),
    .ZN(_10216_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19114_ (.A1(_10210_),
    .A2(_10216_),
    .A3(net20560),
    .ZN(_10217_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19115_ (.A1(_10204_),
    .A2(_10217_),
    .ZN(_10218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19116_ (.A1(_10195_),
    .A2(_10218_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19117_ (.A1(net20081),
    .A2(net20290),
    .A3(net20456),
    .ZN(_10219_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19118_ (.A1(_10093_),
    .A2(_10219_),
    .A3(net20573),
    .ZN(_10220_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19119_ (.A1(net20810),
    .A2(net20158),
    .ZN(_10221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19120_ (.A1(_10221_),
    .A2(net20683),
    .B(_07717_),
    .ZN(_10222_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19121_ (.A1(_09793_),
    .A2(net535),
    .A3(net20468),
    .ZN(_10223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19122_ (.A1(net20293),
    .A2(net20683),
    .ZN(_10224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19123_ (.A1(_10222_),
    .A2(_10223_),
    .A3(_10224_),
    .ZN(_10225_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19124_ (.A1(_10220_),
    .A2(_10225_),
    .A3(net20841),
    .ZN(_10226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19125_ (.A1(net20288),
    .A2(net20079),
    .A3(net20695),
    .ZN(_10227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19126_ (.A1(_10219_),
    .A2(_10227_),
    .A3(net20679),
    .ZN(_10228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19127_ (.A1(_09800_),
    .A2(net20461),
    .B(net20671),
    .ZN(_10229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19128_ (.A1(_10154_),
    .A2(net20284),
    .ZN(_10230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19129_ (.A1(_10229_),
    .A2(_10230_),
    .ZN(_10231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19130_ (.A1(_10228_),
    .A2(_10231_),
    .A3(_09762_),
    .ZN(_10232_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19131_ (.A1(_10226_),
    .A2(_10232_),
    .A3(net20668),
    .ZN(_10233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19132_ (.A1(_09867_),
    .A2(net20469),
    .B(net20680),
    .ZN(_10234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19133_ (.A1(_10012_),
    .A2(_09746_),
    .ZN(_10235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19134_ (.A1(_10235_),
    .A2(net20683),
    .ZN(_10236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19135_ (.A1(_10234_),
    .A2(_10236_),
    .B(_09762_),
    .ZN(_10237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19136_ (.A1(net20065),
    .A2(net20683),
    .ZN(_10238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19137_ (.A1(net20469),
    .A2(net20703),
    .B(_07717_),
    .ZN(_10239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19138_ (.A1(_10238_),
    .A2(_10239_),
    .ZN(_10240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19139_ (.A1(_10237_),
    .A2(_10240_),
    .B(net20668),
    .ZN(_10241_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19140_ (.I(_09912_),
    .ZN(_10242_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19141_ (.A1(_10120_),
    .A2(_10242_),
    .ZN(_10243_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19142_ (.A1(_10081_),
    .A2(_09942_),
    .ZN(_10244_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19143_ (.A1(_10243_),
    .A2(_10244_),
    .B(net20678),
    .ZN(_10245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19144_ (.A1(net662),
    .A2(net20075),
    .ZN(_10246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19145_ (.A1(_10246_),
    .A2(_10031_),
    .ZN(_10247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19146_ (.A1(_10247_),
    .A2(net20577),
    .ZN(_10248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19147_ (.A1(_10248_),
    .A2(_10245_),
    .ZN(_10249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19148_ (.A1(_10249_),
    .A2(_09762_),
    .ZN(_10250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19149_ (.A1(_10250_),
    .A2(_10241_),
    .ZN(_10251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19150_ (.A1(_10251_),
    .A2(_10233_),
    .B(_07744_),
    .ZN(_10252_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19151_ (.A1(_09959_),
    .A2(_09942_),
    .A3(net20681),
    .Z(_10253_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _19152_ (.A1(net20071),
    .A2(net20461),
    .A3(_09878_),
    .Z(_10254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19153_ (.A1(_10253_),
    .A2(_10254_),
    .A3(net20679),
    .ZN(_10255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19154_ (.A1(_10255_),
    .A2(net20841),
    .ZN(_10256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19155_ (.A1(_09915_),
    .A2(net20288),
    .ZN(_10257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19156_ (.A1(_10254_),
    .A2(_10257_),
    .B(net20679),
    .ZN(_10258_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19157_ (.A1(_10256_),
    .A2(_10258_),
    .ZN(_10259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19158_ (.A1(_09912_),
    .A2(net20681),
    .ZN(_10260_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19159_ (.I(_10260_),
    .ZN(_10261_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19160_ (.A1(_10261_),
    .A2(_09842_),
    .Z(_10262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19161_ (.A1(_09901_),
    .A2(_07717_),
    .ZN(_10263_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19162_ (.A1(_10262_),
    .A2(_10263_),
    .ZN(_10264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19163_ (.A1(net20681),
    .A2(_15661_[0]),
    .ZN(_10265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19164_ (.A1(_10265_),
    .A2(net20678),
    .ZN(_10266_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19165_ (.A1(_10170_),
    .A2(_10266_),
    .ZN(_10267_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19166_ (.A1(_10264_),
    .A2(_10267_),
    .B(_09762_),
    .ZN(_10268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19167_ (.A1(_10268_),
    .A2(net20563),
    .ZN(_10269_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19168_ (.A1(_10259_),
    .A2(_10269_),
    .ZN(_10270_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19169_ (.I(_09943_),
    .ZN(_10271_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19170_ (.A1(_09839_),
    .A2(net20577),
    .A3(_10271_),
    .ZN(_10272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19171_ (.A1(_10242_),
    .A2(net20458),
    .ZN(_10273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19172_ (.A1(_10093_),
    .A2(net20678),
    .A3(_10273_),
    .ZN(_10274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19173_ (.A1(_10272_),
    .A2(_10274_),
    .B(_09762_),
    .ZN(_10275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19174_ (.A1(_10103_),
    .A2(net20469),
    .ZN(_10276_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19175_ (.A1(_10124_),
    .A2(_09942_),
    .B(_10276_),
    .ZN(_10277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19176_ (.A1(_10277_),
    .A2(net20572),
    .ZN(_10278_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19177_ (.A1(_09982_),
    .A2(net20679),
    .B(net20837),
    .ZN(_10279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19178_ (.A1(_10278_),
    .A2(_10279_),
    .ZN(_10280_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19179_ (.A1(_10280_),
    .A2(net20668),
    .ZN(_10281_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19180_ (.A1(_10275_),
    .A2(_10281_),
    .B(_07744_),
    .ZN(_10282_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19181_ (.A1(_10270_),
    .A2(_10282_),
    .ZN(_10283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19182_ (.A1(_10283_),
    .A2(_10252_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19183_ (.A1(_10098_),
    .A2(net20570),
    .A3(_09946_),
    .ZN(_10284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19184_ (.A1(_10044_),
    .A2(_10223_),
    .A3(net20679),
    .ZN(_10285_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19185_ (.A1(_10284_),
    .A2(_10285_),
    .A3(net20668),
    .ZN(_10286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19186_ (.A1(_09914_),
    .A2(net20679),
    .Z(_10287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19187_ (.A1(_10125_),
    .A2(_10287_),
    .B(net20668),
    .ZN(_10288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19188_ (.A1(_09828_),
    .A2(net20079),
    .ZN(_10289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19189_ (.A1(_09867_),
    .A2(net20684),
    .ZN(_10290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19190_ (.A1(_10221_),
    .A2(net20683),
    .B(net20679),
    .ZN(_10291_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19191_ (.A1(_10289_),
    .A2(_10290_),
    .A3(_10291_),
    .ZN(_10292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19192_ (.A1(_10288_),
    .A2(_10292_),
    .ZN(_10293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19193_ (.A1(_10293_),
    .A2(_10286_),
    .B(net20649),
    .ZN(_10294_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19194_ (.A1(_09885_),
    .A2(_09912_),
    .A3(net20455),
    .Z(_10295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19195_ (.A1(_10046_),
    .A2(_07717_),
    .ZN(_10296_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19196_ (.A1(_10295_),
    .A2(_10296_),
    .ZN(_10297_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19197_ (.A1(_09865_),
    .A2(net19438),
    .ZN(_10298_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19198_ (.A1(_10297_),
    .A2(_10298_),
    .B(net20668),
    .ZN(_10299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19199_ (.A1(_10299_),
    .A2(net20646),
    .ZN(_10300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19200_ (.A1(_09885_),
    .A2(net20449),
    .A3(net20465),
    .ZN(_10301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19201_ (.A1(_10301_),
    .A2(_10040_),
    .ZN(_10302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19202_ (.A1(_10302_),
    .A2(net20677),
    .ZN(_10303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19203_ (.A1(net20465),
    .A2(net20705),
    .ZN(_10304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19204_ (.A1(_10142_),
    .A2(_07717_),
    .A3(_10304_),
    .ZN(_10305_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19205_ (.A1(_10303_),
    .A2(net20562),
    .A3(_10305_),
    .Z(_10306_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19206_ (.A1(_10300_),
    .A2(_10306_),
    .ZN(_10307_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19207_ (.A1(_10294_),
    .A2(_10307_),
    .B(_07744_),
    .ZN(_10308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19208_ (.A1(net20681),
    .A2(_15671_[0]),
    .Z(_10309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19209_ (.A1(net20469),
    .A2(_10047_),
    .B(_10309_),
    .ZN(_10310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19210_ (.A1(_10310_),
    .A2(_09996_),
    .B(net20562),
    .ZN(_10311_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19211_ (.I(_10263_),
    .ZN(_10312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19212_ (.A1(net19432),
    .A2(net19877),
    .ZN(_10313_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19213_ (.A1(_10312_),
    .A2(_10048_),
    .A3(_10313_),
    .ZN(_10314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19214_ (.A1(_10311_),
    .A2(_10314_),
    .ZN(_10315_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19215_ (.I(_09862_),
    .ZN(_10316_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19216_ (.A1(_10316_),
    .A2(_10126_),
    .A3(_09893_),
    .ZN(_10317_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19217_ (.A1(_10012_),
    .A2(net20683),
    .ZN(_10318_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19218_ (.I(_10318_),
    .ZN(_10319_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19219_ (.A1(net20683),
    .A2(net20088),
    .B(net20574),
    .ZN(_10320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19220_ (.A1(_10319_),
    .A2(_10320_),
    .B(net20668),
    .ZN(_10321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19221_ (.A1(_10317_),
    .A2(_10321_),
    .ZN(_10322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19222_ (.A1(_10315_),
    .A2(_10322_),
    .A3(_09762_),
    .ZN(_10323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19223_ (.A1(net20077),
    .A2(net20680),
    .ZN(_10324_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19224_ (.A1(_10318_),
    .A2(_10324_),
    .ZN(_10325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19225_ (.A1(net20287),
    .A2(net20683),
    .ZN(_10326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19226_ (.A1(_10325_),
    .A2(_10326_),
    .B(net20562),
    .ZN(_10327_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19227_ (.A1(_10238_),
    .A2(net20566),
    .A3(net20068),
    .ZN(_10328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19228_ (.A1(_10327_),
    .A2(_10328_),
    .B(_09762_),
    .ZN(_10329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19229_ (.A1(net19432),
    .A2(net20066),
    .ZN(_10330_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19230_ (.A1(_09867_),
    .A2(_10221_),
    .B(net20469),
    .ZN(_10331_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19231_ (.A1(_10330_),
    .A2(_10331_),
    .A3(net20680),
    .ZN(_10332_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19232_ (.A1(net20292),
    .A2(_09885_),
    .A3(net20467),
    .ZN(_10333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19233_ (.A1(_10333_),
    .A2(_10086_),
    .A3(net20571),
    .ZN(_10334_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19234_ (.A1(_10332_),
    .A2(net20563),
    .A3(_10334_),
    .ZN(_10335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19235_ (.A1(_10329_),
    .A2(_10335_),
    .ZN(_10336_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19236_ (.A1(_10323_),
    .A2(_10336_),
    .A3(_00399_),
    .ZN(_10337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19237_ (.A1(_10308_),
    .A2(_10337_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _19238_ (.I(\sa00_sr[7] ),
    .ZN(_10338_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19239_ (.I(\sa00_sr[0] ),
    .ZN(_10339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19240_ (.A1(_10339_),
    .A2(_10338_),
    .ZN(_10340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19241_ (.A1(net21471),
    .A2(net21481),
    .ZN(_10341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19242_ (.A1(_10341_),
    .A2(_10340_),
    .ZN(_10342_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _19243_ (.I(\sa30_sr[1] ),
    .ZN(_10343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19244_ (.A1(_10343_),
    .A2(\sa20_sr[1] ),
    .ZN(_10344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19245_ (.I(\sa20_sr[1] ),
    .ZN(_10345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19246_ (.A1(_10345_),
    .A2(net21310),
    .ZN(_10346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19247_ (.A1(_10346_),
    .A2(_10344_),
    .ZN(_10347_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19248_ (.A1(_10342_),
    .A2(net20919),
    .ZN(_10348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19249_ (.A1(net21471),
    .A2(_10339_),
    .ZN(_10349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19250_ (.A1(_10338_),
    .A2(net21481),
    .ZN(_10350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19251_ (.A1(_10350_),
    .A2(_10349_),
    .ZN(_10351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19252_ (.A1(_10345_),
    .A2(_10343_),
    .ZN(_10352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19253_ (.A1(\sa20_sr[1] ),
    .A2(net21310),
    .ZN(_10353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19254_ (.A1(_10353_),
    .A2(_10352_),
    .ZN(_10354_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19255_ (.A1(_10351_),
    .A2(net20918),
    .ZN(_10355_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19256_ (.A1(_10348_),
    .A2(_10355_),
    .ZN(_10356_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19257_ (.I(\sa10_sr[0] ),
    .ZN(_10357_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17608 (.I(_15741_[0]),
    .Z(net17608));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19259_ (.A1(net21415),
    .A2(_10357_),
    .ZN(_10359_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19260_ (.I(\sa10_sr[7] ),
    .ZN(_10360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19261_ (.A1(_10360_),
    .A2(net21430),
    .ZN(_10361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19262_ (.A1(_10361_),
    .A2(_10359_),
    .ZN(_10362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19263_ (.A1(net20917),
    .A2(net21429),
    .ZN(_10363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19264_ (.A1(_10357_),
    .A2(_10360_),
    .ZN(_10364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19265_ (.A1(net21415),
    .A2(net21432),
    .ZN(_10365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19266_ (.A1(_10364_),
    .A2(_10365_),
    .ZN(_10366_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19267_ (.I(\sa10_sr[1] ),
    .ZN(_10367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19268_ (.A1(net21096),
    .A2(net20916),
    .ZN(_10368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19269_ (.A1(_10363_),
    .A2(_10368_),
    .ZN(_10369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19270_ (.A1(_10369_),
    .A2(_10356_),
    .ZN(_10370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19271_ (.A1(_10351_),
    .A2(net20918),
    .ZN(_10371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19272_ (.A1(_10342_),
    .A2(net20919),
    .ZN(_10372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19273_ (.A1(_10371_),
    .A2(_10372_),
    .ZN(_10373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19274_ (.A1(net20916),
    .A2(net21429),
    .ZN(_10374_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19275_ (.A1(net20917),
    .A2(net21096),
    .ZN(_10375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19276_ (.A1(_10374_),
    .A2(_10375_),
    .ZN(_10376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19277_ (.A1(_10376_),
    .A2(_10373_),
    .ZN(_10377_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _19278_ (.I(net21490),
    .ZN(_10378_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17588 (.I(_11247_),
    .Z(net17588));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19280_ (.A1(_10370_),
    .A2(_10377_),
    .A3(_10378_),
    .ZN(_10380_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17559 (.I(net654),
    .Z(net17559));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19282_ (.A1(\text_in_r[121] ),
    .A2(net21500),
    .ZN(_10382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19283_ (.A1(_10382_),
    .A2(_10380_),
    .ZN(_10383_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19284_ (.I(net21222),
    .ZN(_10384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19285_ (.A1(net20064),
    .A2(_10384_),
    .ZN(_10385_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19286_ (.A1(net20282),
    .A2(net21222),
    .A3(net21063),
    .ZN(_10386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19287_ (.A1(_10385_),
    .A2(_10386_),
    .ZN(_15679_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19288_ (.A1(net21102),
    .A2(net21097),
    .ZN(_10387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19289_ (.A1(net21470),
    .A2(net21413),
    .ZN(_10388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19290_ (.A1(_10387_),
    .A2(_10388_),
    .ZN(_10389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19291_ (.A1(net21312),
    .A2(_10389_),
    .ZN(_10390_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19292_ (.I(\sa30_sr[0] ),
    .ZN(_10391_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19293_ (.A1(_10387_),
    .A2(net21062),
    .A3(_10388_),
    .ZN(_10392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19294_ (.A1(_10390_),
    .A2(_10392_),
    .ZN(_10393_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19295_ (.I(\sa20_sr[0] ),
    .ZN(_10394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19296_ (.A1(net21061),
    .A2(net21098),
    .ZN(_10395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19297_ (.A1(net21432),
    .A2(net21372),
    .ZN(_10396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19298_ (.A1(net21060),
    .A2(net20959),
    .ZN(_10397_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19299_ (.I(_10397_),
    .ZN(_10398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19300_ (.A1(_10398_),
    .A2(_10393_),
    .ZN(_10399_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19301_ (.A1(_10397_),
    .A2(_10392_),
    .A3(_10390_),
    .ZN(_10400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19302_ (.A1(_10400_),
    .A2(_10399_),
    .ZN(_10401_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17565 (.I(_11855_),
    .Z(net17565));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17625 (.I(_06888_),
    .Z(net17625));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19305_ (.A1(net21074),
    .A2(_10401_),
    .ZN(_10404_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17552 (.I(_12289_),
    .Z(net17552));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19307_ (.A1(net21074),
    .A2(\text_in_r[120] ),
    .Z(_10406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19308_ (.A1(_10404_),
    .A2(net21114),
    .A3(_10406_),
    .ZN(_10407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19309_ (.A1(net21066),
    .A2(_10400_),
    .A3(_10399_),
    .ZN(_10408_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17560 (.I(_12218_),
    .Z(net17560));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17555 (.I(net17554),
    .Z(net17555));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17548 (.I(_13047_),
    .Z(net17548));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19313_ (.A1(net21500),
    .A2(\text_in_r[120] ),
    .ZN(_10412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19314_ (.A1(_10408_),
    .A2(net21223),
    .A3(_10412_),
    .ZN(_10413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19315_ (.A1(_10413_),
    .A2(_10407_),
    .ZN(_15682_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19316_ (.I(\sa00_sr[1] ),
    .ZN(_10414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19317_ (.A1(_10414_),
    .A2(net21428),
    .ZN(_10415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19318_ (.A1(_10367_),
    .A2(net21477),
    .ZN(_10416_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19319_ (.I(net21367),
    .ZN(_10417_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19320_ (.A1(net20958),
    .A2(net20957),
    .A3(net21058),
    .ZN(_10418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19321_ (.A1(_10367_),
    .A2(_10414_),
    .ZN(_10419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19322_ (.A1(net21427),
    .A2(net21477),
    .ZN(_10420_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19323_ (.A1(net20956),
    .A2(net21367),
    .A3(net21057),
    .ZN(_10421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19324_ (.A1(_10418_),
    .A2(_10421_),
    .ZN(_10422_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _19325_ (.I(\sa30_sr[2] ),
    .ZN(_10423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19326_ (.A1(_10423_),
    .A2(net21423),
    .ZN(_10424_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19327_ (.I(\sa10_sr[2] ),
    .ZN(_10425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19328_ (.A1(_10425_),
    .A2(\sa30_sr[2] ),
    .ZN(_10426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19329_ (.A1(_10424_),
    .A2(_10426_),
    .ZN(_10427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19330_ (.I(net20914),
    .ZN(_10428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19331_ (.A1(_10422_),
    .A2(_10428_),
    .ZN(_10429_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19332_ (.A1(_10418_),
    .A2(_10421_),
    .A3(_10427_),
    .ZN(_10430_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17546 (.I(_13096_),
    .Z(net17546));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19334_ (.A1(_10429_),
    .A2(_10430_),
    .B(net21502),
    .ZN(_10432_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19335_ (.I(\text_in_r[122] ),
    .ZN(_10433_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19336_ (.A1(_10433_),
    .A2(net21502),
    .Z(_10434_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19337_ (.A1(_10432_),
    .A2(_10434_),
    .B(net21112),
    .ZN(_10435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19338_ (.A1(_10429_),
    .A2(_10430_),
    .ZN(_10436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19339_ (.A1(_10436_),
    .A2(net21074),
    .ZN(_10437_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19340_ (.I(_10434_),
    .ZN(_10438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19341_ (.A1(_10437_),
    .A2(net21221),
    .A3(_10438_),
    .ZN(_10439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19342_ (.A1(_10435_),
    .A2(_10439_),
    .ZN(_10440_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17629 (.I(_06824_),
    .Z(net17629));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19344_ (.A1(_10406_),
    .A2(net21223),
    .A3(_10404_),
    .ZN(_10441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19345_ (.A1(net21114),
    .A2(_10408_),
    .A3(_10412_),
    .ZN(_10442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19346_ (.A1(_10441_),
    .A2(_10442_),
    .ZN(_15673_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19347_ (.A1(_10432_),
    .A2(_10434_),
    .B(net21221),
    .ZN(_10443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19348_ (.A1(_10437_),
    .A2(net21112),
    .A3(_10438_),
    .ZN(_10444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19349_ (.A1(_10443_),
    .A2(_10444_),
    .ZN(_10445_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17595 (.I(_10604_),
    .Z(net17595));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19351_ (.A1(net19429),
    .A2(_10445_),
    .ZN(_10446_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19352_ (.I(_10446_),
    .ZN(_10447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19353_ (.A1(_10447_),
    .A2(net19425),
    .ZN(_10448_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19354_ (.A1(\sa20_sr[3] ),
    .A2(\sa30_sr[3] ),
    .Z(_10449_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19355_ (.I(\sa00_sr[2] ),
    .ZN(_10450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19356_ (.A1(net21103),
    .A2(_10450_),
    .ZN(_10451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19357_ (.A1(net21470),
    .A2(\sa00_sr[2] ),
    .ZN(_10452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19358_ (.A1(_10451_),
    .A2(_10452_),
    .ZN(_10453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19359_ (.A1(_10449_),
    .A2(_10453_),
    .ZN(_10454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19360_ (.A1(_10450_),
    .A2(net21470),
    .ZN(_10455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19361_ (.A1(net21103),
    .A2(\sa00_sr[2] ),
    .ZN(_10456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19362_ (.A1(_10455_),
    .A2(_10456_),
    .ZN(_10457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19363_ (.I(\sa20_sr[3] ),
    .ZN(_10458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19364_ (.I(\sa30_sr[3] ),
    .ZN(_10459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19365_ (.A1(_10458_),
    .A2(_10459_),
    .ZN(_10460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19366_ (.A1(net21365),
    .A2(net21304),
    .ZN(_10461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19367_ (.A1(_10460_),
    .A2(_10461_),
    .ZN(_10462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19368_ (.A1(_10457_),
    .A2(_10462_),
    .ZN(_10463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19369_ (.A1(_10454_),
    .A2(_10463_),
    .ZN(_10464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19370_ (.I(_10464_),
    .ZN(_10465_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19371_ (.I(\sa10_sr[3] ),
    .ZN(_10466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19372_ (.A1(_10466_),
    .A2(net21413),
    .ZN(_10467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19373_ (.A1(net504),
    .A2(net21421),
    .ZN(_10468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19374_ (.A1(_10467_),
    .A2(_10468_),
    .ZN(_10469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19375_ (.A1(_10469_),
    .A2(net21425),
    .ZN(_10470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19376_ (.A1(net504),
    .A2(_10466_),
    .ZN(_10471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19377_ (.A1(net21414),
    .A2(net21421),
    .ZN(_10472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19378_ (.A1(_10471_),
    .A2(_10472_),
    .ZN(_10473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19379_ (.A1(_10473_),
    .A2(net21056),
    .ZN(_10474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19380_ (.A1(_10470_),
    .A2(_10474_),
    .ZN(_10475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19381_ (.A1(_10465_),
    .A2(net20645),
    .ZN(_10476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19382_ (.I(_10475_),
    .ZN(_10477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19383_ (.A1(_10477_),
    .A2(_10464_),
    .ZN(_10478_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17823 (.I(net17820),
    .Z(net17823));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19385_ (.A1(_10476_),
    .A2(_10478_),
    .A3(net21080),
    .ZN(_10480_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19386_ (.I(net21220),
    .ZN(_10481_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17570 (.I(net17569),
    .Z(net17570));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17539 (.I(_13258_),
    .Z(net17539));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19389_ (.A1(net21501),
    .A2(\text_in_r[123] ),
    .ZN(_10484_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19390_ (.A1(_10480_),
    .A2(_10481_),
    .A3(_10484_),
    .ZN(_10485_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19391_ (.A1(_10465_),
    .A2(_10477_),
    .ZN(_10486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19392_ (.A1(_10464_),
    .A2(_10475_),
    .ZN(_10487_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19393_ (.A1(_10486_),
    .A2(net21080),
    .A3(_10487_),
    .ZN(_10488_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17536 (.I(_13765_),
    .Z(net17536));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19395_ (.A1(net21080),
    .A2(\text_in_r[123] ),
    .Z(_10490_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19396_ (.A1(_10488_),
    .A2(net21220),
    .A3(_10490_),
    .ZN(_10491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19397_ (.A1(_10485_),
    .A2(_10491_),
    .ZN(_10492_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17571 (.I(_11502_),
    .Z(net17571));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19399_ (.I(_15680_[0]),
    .ZN(_10494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19400_ (.A1(net19869),
    .A2(_10494_),
    .ZN(_10495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19401_ (.A1(_10448_),
    .A2(net19413),
    .A3(net17970),
    .ZN(_10496_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19402_ (.A1(net19869),
    .A2(net19428),
    .ZN(_10497_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19403_ (.I(_15675_[0]),
    .ZN(_10498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19404_ (.A1(net19866),
    .A2(_10498_),
    .ZN(_10499_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19405_ (.A1(_10497_),
    .A2(_10499_),
    .ZN(_10500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19406_ (.A1(_10480_),
    .A2(net21220),
    .A3(_10484_),
    .ZN(_10501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19407_ (.A1(_10488_),
    .A2(_10481_),
    .A3(_10490_),
    .ZN(_10502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19408_ (.A1(_10501_),
    .A2(_10502_),
    .ZN(_10503_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17598 (.I(_10539_),
    .Z(net17598));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17920 (.I(_12145_),
    .Z(net17920));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19411_ (.A1(_10500_),
    .A2(net19402),
    .ZN(_10506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19412_ (.A1(net20280),
    .A2(net20062),
    .A3(_15677_[0]),
    .ZN(_10507_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19413_ (.I(_10507_),
    .ZN(_10508_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17535 (.I(_13783_),
    .Z(net17535));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19415_ (.A1(_10508_),
    .A2(net19413),
    .ZN(_10510_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19416_ (.A1(net21470),
    .A2(\sa00_sr[3] ),
    .Z(_10511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19417_ (.I(\sa20_sr[4] ),
    .ZN(_10512_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19418_ (.A1(_10511_),
    .A2(net21052),
    .Z(_10513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19419_ (.A1(_10511_),
    .A2(net21052),
    .ZN(_10514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19420_ (.A1(_10513_),
    .A2(_10514_),
    .ZN(_10515_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19421_ (.I(_10515_),
    .ZN(_10516_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19422_ (.A1(net21418),
    .A2(net21303),
    .Z(_10517_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19423_ (.A1(_10473_),
    .A2(_10517_),
    .Z(_10518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19424_ (.A1(_10516_),
    .A2(_10518_),
    .ZN(_10519_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19425_ (.A1(_10469_),
    .A2(_10517_),
    .Z(_10520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19426_ (.A1(_10520_),
    .A2(net20913),
    .ZN(_10521_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17534 (.I(_13812_),
    .Z(net17534));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17857 (.I(_14536_),
    .Z(net17857));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19429_ (.A1(_10519_),
    .A2(_10521_),
    .A3(net21065),
    .ZN(_10524_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17849 (.I(_14596_),
    .Z(net17849));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17531 (.I(_13964_),
    .Z(net17531));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19432_ (.A1(net21500),
    .A2(\text_in_r[124] ),
    .ZN(_10527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19433_ (.A1(_10524_),
    .A2(_10527_),
    .ZN(_10528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19434_ (.A1(_10528_),
    .A2(net21219),
    .ZN(_10529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19435_ (.I(net21219),
    .ZN(_10530_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19436_ (.A1(_10524_),
    .A2(_10530_),
    .A3(_10527_),
    .ZN(_10531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19437_ (.A1(_10529_),
    .A2(_10531_),
    .ZN(_10532_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17848 (.I(_14608_),
    .Z(net17848));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19439_ (.A1(_10510_),
    .A2(net19862),
    .Z(_10534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19440_ (.A1(_10496_),
    .A2(_10506_),
    .A3(_10534_),
    .ZN(_10535_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19441_ (.A1(_15676_[0]),
    .A2(net20280),
    .A3(net20062),
    .ZN(_10536_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _19442_ (.I(_10536_),
    .ZN(_10537_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17529 (.I(_14086_),
    .Z(net17529));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _19444_ (.A1(net19413),
    .A2(_10537_),
    .B(_10532_),
    .ZN(_10539_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17846 (.I(_14644_),
    .Z(net17846));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19446_ (.A1(net19402),
    .A2(net18419),
    .ZN(_10541_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19447_ (.A1(\sa10_sr[4] ),
    .A2(\sa00_sr[4] ),
    .Z(_10542_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19448_ (.A1(\sa20_sr[5] ),
    .A2(\sa30_sr[5] ),
    .Z(_10543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19449_ (.A1(\sa20_sr[5] ),
    .A2(\sa30_sr[5] ),
    .ZN(_10544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19450_ (.A1(_10543_),
    .A2(_10544_),
    .ZN(_10545_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19451_ (.A1(net21417),
    .A2(_10545_),
    .Z(_10546_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19452_ (.A1(net21051),
    .A2(_10546_),
    .Z(_10547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19453_ (.A1(_10547_),
    .A2(net21065),
    .ZN(_10548_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17844 (.I(_14680_),
    .Z(net17844));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19455_ (.A1(net21065),
    .A2(\text_in_r[125] ),
    .Z(_10550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19456_ (.A1(_10548_),
    .A2(_10550_),
    .ZN(_10551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19457_ (.I(net21218),
    .ZN(_10552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19458_ (.A1(_10551_),
    .A2(_10552_),
    .ZN(_10553_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19459_ (.A1(_10548_),
    .A2(net21218),
    .A3(_10550_),
    .ZN(_10554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19460_ (.A1(_10553_),
    .A2(_10554_),
    .ZN(_10555_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _19461_ (.I(_10555_),
    .ZN(_10556_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17527 (.I(_14388_),
    .Z(net17527));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19463_ (.A1(net17598),
    .A2(_10541_),
    .B(net19857),
    .ZN(_10558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19464_ (.A1(_10535_),
    .A2(_10558_),
    .ZN(_10559_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19465_ (.I(_15685_[0]),
    .ZN(_10560_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19466_ (.A1(net20280),
    .A2(net20062),
    .A3(_10560_),
    .ZN(_10561_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19467_ (.A1(_10561_),
    .A2(net19400),
    .Z(_10562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19468_ (.A1(_10448_),
    .A2(net17597),
    .ZN(_10563_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17530 (.I(_14073_),
    .Z(net17530));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19470_ (.A1(net19866),
    .A2(_15677_[0]),
    .Z(_10565_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17528 (.I(_14232_),
    .Z(net17528));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19472_ (.A1(_10565_),
    .A2(net19413),
    .ZN(_10567_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19473_ (.A1(_10563_),
    .A2(_10532_),
    .A3(_10567_),
    .ZN(_10568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19474_ (.A1(_10565_),
    .A2(net19401),
    .ZN(_10569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19475_ (.A1(_10528_),
    .A2(_10530_),
    .ZN(_10570_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19476_ (.A1(_10524_),
    .A2(net21219),
    .A3(_10527_),
    .ZN(_10571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19477_ (.A1(_10570_),
    .A2(_10571_),
    .ZN(_10572_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17525 (.I(_14552_),
    .Z(net17525));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19479_ (.A1(_10569_),
    .A2(net19840),
    .Z(_10574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19480_ (.A1(net19869),
    .A2(_15683_[0]),
    .ZN(_10575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19481_ (.A1(_10575_),
    .A2(net19413),
    .Z(_10576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19482_ (.A1(_10448_),
    .A2(_10576_),
    .ZN(_10577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19483_ (.A1(_10574_),
    .A2(_10577_),
    .ZN(_10578_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17830 (.I(_15330_),
    .Z(net17830));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19485_ (.A1(_10568_),
    .A2(_10578_),
    .A3(net19857),
    .ZN(_10580_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _19486_ (.A1(\sa10_sr[5] ),
    .A2(\sa00_sr[5] ),
    .ZN(_10581_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _19487_ (.A1(\sa20_sr[6] ),
    .A2(\sa30_sr[6] ),
    .ZN(_10582_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19488_ (.A1(\sa10_sr[6] ),
    .A2(_10582_),
    .Z(_10583_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19489_ (.A1(_10581_),
    .A2(_10583_),
    .Z(_10584_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17832 (.I(_15322_),
    .Z(net17832));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17522 (.I(_14647_),
    .Z(net17522));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17521 (.I(_14790_),
    .Z(net17521));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19493_ (.A1(net21492),
    .A2(\text_in_r[126] ),
    .Z(_10588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19494_ (.A1(_10584_),
    .A2(net21065),
    .B(_10588_),
    .ZN(_10589_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19495_ (.A1(net21216),
    .A2(_10589_),
    .Z(_10590_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18392 (.I(_15913_[0]),
    .Z(net18392));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19497_ (.A1(_10559_),
    .A2(_10580_),
    .A3(net20643),
    .ZN(_10592_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18535 (.I(net18532),
    .Z(net18535));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17523 (.I(_14588_),
    .Z(net17523));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19500_ (.A1(net19866),
    .A2(net19427),
    .ZN(_10595_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _19501_ (.I(_15683_[0]),
    .ZN(_10596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19502_ (.A1(net19869),
    .A2(_10596_),
    .ZN(_10597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19503_ (.A1(net18940),
    .A2(net17965),
    .Z(_10598_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19504_ (.A1(net18942),
    .A2(net19418),
    .A3(net18350),
    .ZN(_10599_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17520 (.I(_14812_),
    .Z(net17520));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _19506_ (.A1(net19413),
    .A2(_10598_),
    .B(_10599_),
    .C(net19865),
    .ZN(_10601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19507_ (.A1(net19866),
    .A2(_10494_),
    .ZN(_10602_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18518 (.I(_03985_),
    .Z(net18518));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19509_ (.A1(_10602_),
    .A2(net505),
    .Z(_10604_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17524 (.I(net17523),
    .Z(net17524));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19511_ (.A1(net17595),
    .A2(net19865),
    .ZN(_10606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19512_ (.A1(net19869),
    .A2(_10498_),
    .ZN(_10607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19513_ (.I(_10607_),
    .ZN(_10608_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19514_ (.A1(net18348),
    .A2(_10608_),
    .B(net19420),
    .ZN(_10609_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17532 (.I(_13862_),
    .Z(net17532));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19516_ (.A1(_10606_),
    .A2(_10609_),
    .B(net20059),
    .ZN(_10611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19517_ (.A1(_10601_),
    .A2(_10611_),
    .ZN(_10612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19518_ (.A1(_10447_),
    .A2(net19428),
    .ZN(_10613_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17519 (.I(net454),
    .Z(net17519));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19520_ (.A1(net19869),
    .A2(net19425),
    .ZN(_10615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19521_ (.A1(_10613_),
    .A2(net19403),
    .A3(net18938),
    .ZN(_10616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19522_ (.A1(net19869),
    .A2(net18423),
    .ZN(_10617_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19523_ (.I(_10617_),
    .ZN(_10618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19524_ (.A1(_10618_),
    .A2(net19415),
    .B(net19840),
    .ZN(_10619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19525_ (.A1(_10616_),
    .A2(_10619_),
    .ZN(_10620_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19526_ (.I(_15676_[0]),
    .ZN(_10621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19527_ (.A1(_10621_),
    .A2(net19868),
    .ZN(_10622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19528_ (.A1(_10622_),
    .A2(net19411),
    .ZN(_10623_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19529_ (.A1(_10623_),
    .A2(net19840),
    .Z(_10624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19530_ (.A1(net19866),
    .A2(net18422),
    .ZN(_10625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19531_ (.A1(_10617_),
    .A2(_10625_),
    .ZN(_10626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19532_ (.A1(net17957),
    .A2(net19414),
    .ZN(_10627_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17517 (.I(_15213_),
    .Z(net17517));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19534_ (.A1(_10624_),
    .A2(_10627_),
    .B(net19857),
    .ZN(_10629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19535_ (.A1(_10620_),
    .A2(_10629_),
    .ZN(_10630_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _19536_ (.I(_10590_),
    .ZN(_10631_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17508 (.I(_15274_),
    .Z(net17508));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19538_ (.A1(_10612_),
    .A2(_10630_),
    .A3(_10631_),
    .ZN(_10633_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17505 (.I(_15519_),
    .Z(net17505));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17509 (.I(_15254_),
    .Z(net17509));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19541_ (.A1(net21416),
    .A2(\sa00_sr[6] ),
    .Z(_10636_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _19542_ (.A1(net21413),
    .A2(_10636_),
    .Z(_10637_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _19543_ (.A1(net21362),
    .A2(net21298),
    .A3(_10637_),
    .Z(_10638_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17515 (.I(_15221_),
    .Z(net17515));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19545_ (.I0(_10638_),
    .I1(\text_in_r[127] ),
    .S(net21500),
    .Z(_10640_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _19546_ (.A1(net21215),
    .A2(_10640_),
    .ZN(_10641_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17540 (.I(_13210_),
    .Z(net17540));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19548_ (.I(_10641_),
    .ZN(_10643_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19549_ (.A1(_10592_),
    .A2(_10633_),
    .A3(_10643_),
    .ZN(_10644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19550_ (.A1(net19429),
    .A2(net19869),
    .ZN(_10645_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19551_ (.A1(net20281),
    .A2(net20063),
    .A3(_15676_[0]),
    .ZN(_10646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19552_ (.A1(net19412),
    .A2(_10646_),
    .ZN(_10647_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19553_ (.I(_10647_),
    .ZN(_10648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19554_ (.A1(net19869),
    .A2(_10621_),
    .ZN(_10649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19555_ (.A1(_10649_),
    .A2(net19400),
    .Z(_10650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _19556_ (.A1(net18937),
    .A2(_10648_),
    .B(_10650_),
    .C(net19865),
    .ZN(_10651_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19557_ (.I(_10499_),
    .ZN(_10652_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _19558_ (.I(_10597_),
    .ZN(_10653_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17492 (.I(_01135_),
    .Z(net17492));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19560_ (.A1(net17593),
    .A2(_10653_),
    .B(net19421),
    .ZN(_10655_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _19561_ (.I(_10623_),
    .ZN(_10656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19562_ (.A1(net19870),
    .A2(net18425),
    .ZN(_10657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19563_ (.A1(_10656_),
    .A2(_10657_),
    .ZN(_10658_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17545 (.I(_13102_),
    .Z(net17545));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19565_ (.A1(_10655_),
    .A2(_10658_),
    .B(net19845),
    .ZN(_10660_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17497 (.I(_01062_),
    .Z(net17497));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19567_ (.A1(_10651_),
    .A2(_10660_),
    .B(net20059),
    .ZN(_10662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19568_ (.A1(_10595_),
    .A2(net19413),
    .Z(_10663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19569_ (.A1(net21222),
    .A2(_10383_),
    .ZN(_10664_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19570_ (.A1(_10380_),
    .A2(_10384_),
    .A3(_10382_),
    .ZN(_10665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19571_ (.A1(_10664_),
    .A2(_10665_),
    .ZN(_15674_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19572_ (.A1(net19399),
    .A2(net19425),
    .ZN(_10666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19573_ (.A1(_10663_),
    .A2(net18936),
    .ZN(_10667_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17488 (.I(_01231_),
    .Z(net17488));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19575_ (.A1(net19429),
    .A2(net494),
    .ZN(_10669_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19576_ (.A1(_10669_),
    .A2(net19407),
    .A3(_10497_),
    .ZN(_10670_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19577_ (.A1(_10667_),
    .A2(net19847),
    .A3(_10670_),
    .ZN(_10671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19578_ (.A1(net19868),
    .A2(_10596_),
    .ZN(_10672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19579_ (.A1(net17963),
    .A2(net17954),
    .ZN(_10673_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17489 (.I(_01185_),
    .Z(net17489));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19581_ (.A1(_10673_),
    .A2(net19407),
    .B(net19840),
    .ZN(_10675_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19582_ (.A1(_10622_),
    .A2(net19413),
    .Z(_10676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19583_ (.A1(net19431),
    .A2(net19427),
    .A3(net19869),
    .ZN(_10677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19584_ (.A1(_10676_),
    .A2(net18935),
    .ZN(_10678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19585_ (.A1(_10675_),
    .A2(_10678_),
    .ZN(_10679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19586_ (.A1(_10671_),
    .A2(_10679_),
    .A3(net19854),
    .ZN(_10680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19587_ (.A1(_10662_),
    .A2(_10680_),
    .A3(net20643),
    .ZN(_10681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19588_ (.A1(_10615_),
    .A2(net19413),
    .ZN(_10682_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19589_ (.A1(_10682_),
    .A2(net19864),
    .Z(_10683_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19590_ (.A1(net19430),
    .A2(net494),
    .A3(net19869),
    .ZN(_10684_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19591_ (.A1(_10604_),
    .A2(_10684_),
    .ZN(_10685_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17490 (.I(_01165_),
    .Z(net17490));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19593_ (.A1(_10683_),
    .A2(_10685_),
    .B(net20061),
    .ZN(_10687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19594_ (.A1(net19425),
    .A2(net19868),
    .ZN(_10688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19595_ (.A1(net19413),
    .A2(_10688_),
    .Z(_10689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19596_ (.A1(_10689_),
    .A2(_10684_),
    .ZN(_10690_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _19597_ (.I(_15689_[0]),
    .ZN(_10691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19598_ (.A1(net19869),
    .A2(_10691_),
    .ZN(_10692_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19599_ (.A1(_10692_),
    .A2(net19409),
    .Z(_10693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19600_ (.A1(_10693_),
    .A2(net17959),
    .ZN(_10694_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19601_ (.A1(_10690_),
    .A2(_10694_),
    .A3(net19849),
    .ZN(_10695_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17544 (.I(_13124_),
    .Z(net17544));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19603_ (.A1(_10687_),
    .A2(_10695_),
    .B(net20643),
    .ZN(_10697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19604_ (.A1(_10567_),
    .A2(net19863),
    .ZN(_10698_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19605_ (.A1(net19431),
    .A2(net19866),
    .ZN(_10699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19606_ (.A1(_10699_),
    .A2(net19413),
    .Z(_10700_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19607_ (.A1(_10698_),
    .A2(_10700_),
    .ZN(_10701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19608_ (.A1(_10701_),
    .A2(_10616_),
    .ZN(_10702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19609_ (.A1(net19399),
    .A2(net19868),
    .ZN(_10703_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17484 (.I(_01672_),
    .Z(net17484));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19611_ (.A1(_10684_),
    .A2(net19413),
    .A3(net18929),
    .ZN(_10705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19612_ (.A1(net19866),
    .A2(_10691_),
    .ZN(_10706_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19613_ (.A1(net18938),
    .A2(net17951),
    .A3(net19403),
    .ZN(_10707_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19614_ (.A1(_10705_),
    .A2(net19850),
    .A3(_10707_),
    .ZN(_10708_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19615_ (.A1(_10702_),
    .A2(_10708_),
    .A3(net20061),
    .ZN(_10709_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19616_ (.A1(_10697_),
    .A2(_10709_),
    .B(_10643_),
    .ZN(_10710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19617_ (.A1(_10681_),
    .A2(_10710_),
    .ZN(_10711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19618_ (.A1(_10644_),
    .A2(_10711_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _19619_ (.I(_10682_),
    .ZN(_10712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19620_ (.A1(_10613_),
    .A2(_10712_),
    .ZN(_10713_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19621_ (.A1(_10623_),
    .A2(net19864),
    .Z(_10714_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19622_ (.A1(_10713_),
    .A2(_10714_),
    .B(net19857),
    .ZN(_10715_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19623_ (.A1(_10706_),
    .A2(net19412),
    .Z(_10716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19624_ (.I(_15677_[0]),
    .ZN(_10717_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19625_ (.A1(net19869),
    .A2(_10717_),
    .ZN(_10718_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19626_ (.A1(_10716_),
    .A2(net17950),
    .B(net19860),
    .ZN(_10719_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19627_ (.A1(_10677_),
    .A2(net19401),
    .A3(net18343),
    .ZN(_10720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19628_ (.A1(_10719_),
    .A2(_10720_),
    .ZN(_10721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19629_ (.A1(_10715_),
    .A2(_10721_),
    .B(net20643),
    .ZN(_10722_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19630_ (.I(_10497_),
    .ZN(_10723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19631_ (.A1(_10723_),
    .A2(net19413),
    .ZN(_10724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19632_ (.A1(_10724_),
    .A2(_10567_),
    .Z(_10725_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19633_ (.A1(net17593),
    .A2(net500),
    .B(net19403),
    .ZN(_10726_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19634_ (.A1(_10725_),
    .A2(net19850),
    .A3(_10726_),
    .ZN(_10727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19635_ (.A1(_10663_),
    .A2(_10657_),
    .ZN(_10728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19636_ (.A1(net19399),
    .A2(net19869),
    .ZN(_10729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19637_ (.A1(_10604_),
    .A2(net18928),
    .ZN(_10730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19638_ (.A1(_10728_),
    .A2(_10730_),
    .A3(net19864),
    .ZN(_10731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19639_ (.A1(_10727_),
    .A2(_10731_),
    .A3(net19859),
    .ZN(_10732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19640_ (.A1(_10722_),
    .A2(_10732_),
    .B(_10643_),
    .ZN(_10733_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19641_ (.A1(_10613_),
    .A2(net19403),
    .A3(_10684_),
    .ZN(_10734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19642_ (.A1(_10689_),
    .A2(_10657_),
    .B(net20059),
    .ZN(_10735_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19643_ (.A1(_10734_),
    .A2(_10735_),
    .ZN(_10736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19644_ (.A1(_10663_),
    .A2(net18937),
    .ZN(_10737_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19645_ (.A1(_10737_),
    .A2(_10730_),
    .A3(net20059),
    .ZN(_10738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19646_ (.A1(_10736_),
    .A2(_10738_),
    .B(net19864),
    .ZN(_10739_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19647_ (.A1(_10556_),
    .A2(_15699_[0]),
    .A3(net19413),
    .Z(_10740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19648_ (.A1(_10613_),
    .A2(_10576_),
    .ZN(_10741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19649_ (.A1(_10740_),
    .A2(net19861),
    .A3(_10741_),
    .ZN(_10742_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19650_ (.I(_10742_),
    .ZN(_10743_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19651_ (.A1(_10739_),
    .A2(_10743_),
    .B(net20643),
    .ZN(_10744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19652_ (.A1(_10733_),
    .A2(_10744_),
    .ZN(_10745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19653_ (.A1(net19869),
    .A2(net19400),
    .Z(_10746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19654_ (.A1(_10746_),
    .A2(_10669_),
    .ZN(_10747_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19655_ (.A1(_10747_),
    .A2(net19864),
    .Z(_10748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19656_ (.A1(_10446_),
    .A2(net19413),
    .Z(_10749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19657_ (.A1(_10749_),
    .A2(_10666_),
    .ZN(_10750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19658_ (.A1(_10748_),
    .A2(_10750_),
    .ZN(_10751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19659_ (.A1(_10602_),
    .A2(net19413),
    .ZN(_10752_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19660_ (.A1(_10752_),
    .A2(_10723_),
    .Z(_10753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19661_ (.A1(_10656_),
    .A2(net18938),
    .ZN(_10754_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17547 (.I(_13061_),
    .Z(net17547));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19663_ (.A1(_10753_),
    .A2(_10754_),
    .A3(net19850),
    .ZN(_10756_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19664_ (.A1(_10751_),
    .A2(_10756_),
    .A3(net19859),
    .ZN(_10757_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19665_ (.A1(_10650_),
    .A2(net17951),
    .ZN(_10758_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19666_ (.A1(_10758_),
    .A2(net19864),
    .Z(_10759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19667_ (.A1(_10759_),
    .A2(_10496_),
    .ZN(_10760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19668_ (.A1(_10645_),
    .A2(net19400),
    .ZN(_10761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19669_ (.A1(net18342),
    .A2(_10703_),
    .Z(_10762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19670_ (.A1(_10618_),
    .A2(net19413),
    .B(_10532_),
    .ZN(_10763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19671_ (.A1(_10762_),
    .A2(_10763_),
    .B(net19857),
    .ZN(_10764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19672_ (.A1(_10760_),
    .A2(_10764_),
    .ZN(_10765_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19673_ (.A1(_10757_),
    .A2(_10765_),
    .A3(net20643),
    .ZN(_10766_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _19674_ (.I(_10622_),
    .ZN(_10767_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19675_ (.A1(net17592),
    .A2(net17960),
    .B(net19402),
    .ZN(_10768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19676_ (.A1(net17599),
    .A2(net19415),
    .ZN(_10769_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19677_ (.A1(_10768_),
    .A2(net19852),
    .A3(_10769_),
    .ZN(_10770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19678_ (.A1(net19431),
    .A2(net19427),
    .ZN(_10771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19679_ (.A1(net18925),
    .A2(net18933),
    .ZN(_10772_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17491 (.I(_01156_),
    .Z(net17491));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19681_ (.A1(_10772_),
    .A2(net19402),
    .ZN(_10774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19682_ (.A1(_10536_),
    .A2(net19413),
    .Z(_10775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19683_ (.A1(_10775_),
    .A2(net18933),
    .ZN(_10776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19684_ (.A1(_10774_),
    .A2(_10776_),
    .A3(net19862),
    .ZN(_10777_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19685_ (.A1(_10770_),
    .A2(_10777_),
    .A3(net20056),
    .ZN(_10778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19686_ (.A1(_10693_),
    .A2(_10703_),
    .ZN(_10779_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19687_ (.A1(net18925),
    .A2(net19866),
    .A3(net19414),
    .ZN(_10780_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19688_ (.A1(_10779_),
    .A2(_10780_),
    .A3(net19840),
    .ZN(_10781_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19689_ (.A1(net19866),
    .A2(net18424),
    .Z(_10782_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17483 (.I(net472),
    .Z(net17483));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19691_ (.A1(_10782_),
    .A2(net19414),
    .B(net19840),
    .ZN(_10784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19692_ (.A1(_10720_),
    .A2(_10784_),
    .ZN(_10785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19693_ (.A1(_10781_),
    .A2(_10785_),
    .A3(net19858),
    .ZN(_10786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19694_ (.A1(_10778_),
    .A2(_10786_),
    .A3(_10631_),
    .ZN(_10787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19695_ (.A1(_10766_),
    .A2(_10787_),
    .A3(_10643_),
    .ZN(_10788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19696_ (.A1(_10745_),
    .A2(_10788_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19697_ (.A1(_10688_),
    .A2(net17968),
    .ZN(_10789_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19698_ (.A1(_10789_),
    .A2(net19400),
    .A3(_10703_),
    .ZN(_10790_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19699_ (.A1(_10790_),
    .A2(net19860),
    .A3(_10599_),
    .ZN(_10791_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19700_ (.A1(_10669_),
    .A2(_10446_),
    .A3(net19405),
    .ZN(_10792_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19701_ (.A1(_10692_),
    .A2(_10602_),
    .A3(net19413),
    .ZN(_10793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19702_ (.A1(_10792_),
    .A2(_10793_),
    .ZN(_10794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19703_ (.A1(_10794_),
    .A2(net19841),
    .ZN(_10795_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19704_ (.A1(_10791_),
    .A2(_10795_),
    .A3(net20053),
    .ZN(_10796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19705_ (.A1(_10684_),
    .A2(net19423),
    .B(net19840),
    .ZN(_10797_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19706_ (.A1(_10677_),
    .A2(net19401),
    .A3(net17952),
    .ZN(_10798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19707_ (.A1(_10797_),
    .A2(_10798_),
    .ZN(_10799_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19708_ (.A1(_10647_),
    .A2(_10699_),
    .ZN(_10800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19709_ (.A1(_10507_),
    .A2(net19401),
    .ZN(_10801_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19710_ (.I(_10595_),
    .ZN(_10802_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19711_ (.A1(_10801_),
    .A2(_10802_),
    .ZN(_10803_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19712_ (.A1(_10800_),
    .A2(_10803_),
    .B(net19840),
    .ZN(_10804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19713_ (.A1(_10799_),
    .A2(_10804_),
    .ZN(_10805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19714_ (.A1(_10805_),
    .A2(net19857),
    .ZN(_10806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19715_ (.A1(_10796_),
    .A2(_10806_),
    .A3(net20644),
    .ZN(_10807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _19716_ (.A1(net20280),
    .A2(net20062),
    .A3(net18420),
    .ZN(_10808_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19717_ (.A1(net18939),
    .A2(net19412),
    .A3(_10808_),
    .ZN(_10809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19718_ (.A1(_10809_),
    .A2(net19840),
    .ZN(_10810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19719_ (.A1(_10625_),
    .A2(net19404),
    .ZN(_10811_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19720_ (.A1(_10811_),
    .A2(net18931),
    .ZN(_10812_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19721_ (.A1(_10810_),
    .A2(_10812_),
    .ZN(_10813_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19722_ (.A1(_10688_),
    .A2(net19413),
    .A3(net17966),
    .ZN(_10814_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19723_ (.A1(net17958),
    .A2(net18349),
    .A3(net19404),
    .ZN(_10815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19724_ (.A1(_10814_),
    .A2(_10815_),
    .B(net19840),
    .ZN(_10816_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19725_ (.A1(_10813_),
    .A2(_10816_),
    .B(net19857),
    .ZN(_10817_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19726_ (.A1(_10626_),
    .A2(net19413),
    .B(net19840),
    .ZN(_10818_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19727_ (.A1(_10495_),
    .A2(net19401),
    .Z(_10819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19728_ (.A1(_10819_),
    .A2(net18930),
    .ZN(_10820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19729_ (.A1(_10818_),
    .A2(_10820_),
    .ZN(_10821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19730_ (.A1(net18344),
    .A2(_10808_),
    .ZN(_10822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19731_ (.A1(_10822_),
    .A2(net19413),
    .ZN(_10823_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19732_ (.A1(_10688_),
    .A2(net17969),
    .A3(net19400),
    .ZN(_10824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19733_ (.A1(_10823_),
    .A2(_10824_),
    .A3(net19840),
    .ZN(_10825_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19734_ (.A1(_10821_),
    .A2(_10825_),
    .A3(net20053),
    .ZN(_10826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19735_ (.A1(_10817_),
    .A2(_10826_),
    .ZN(_10827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19736_ (.A1(_10827_),
    .A2(_10631_),
    .ZN(_10828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19737_ (.A1(_10807_),
    .A2(_10828_),
    .ZN(_10829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19738_ (.A1(_10829_),
    .A2(net20642),
    .ZN(_10830_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19739_ (.A1(_10749_),
    .A2(_10607_),
    .Z(_10831_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19740_ (.A1(_10672_),
    .A2(net19406),
    .A3(_10536_),
    .Z(_10832_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19741_ (.A1(_10831_),
    .A2(_10832_),
    .B(net19843),
    .ZN(_10833_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19742_ (.A1(_10666_),
    .A2(_10446_),
    .A3(net19407),
    .Z(_10834_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19743_ (.A1(_10834_),
    .A2(net19840),
    .ZN(_10835_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19744_ (.A1(net19406),
    .A2(_15699_[0]),
    .Z(_10836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19745_ (.A1(_10835_),
    .A2(_10836_),
    .ZN(_10837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19746_ (.A1(_10833_),
    .A2(_10837_),
    .A3(net20060),
    .ZN(_10838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19747_ (.A1(_10448_),
    .A2(_10650_),
    .ZN(_10839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19748_ (.A1(_15696_[0]),
    .A2(net19414),
    .B(net19840),
    .ZN(_10840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19749_ (.A1(_10839_),
    .A2(_10840_),
    .B(net20052),
    .ZN(_10841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19750_ (.A1(_10729_),
    .A2(net19407),
    .Z(_10842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19751_ (.A1(_10842_),
    .A2(net18934),
    .ZN(_10843_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19752_ (.A1(_10843_),
    .A2(net19848),
    .A3(_10599_),
    .ZN(_10844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19753_ (.A1(_10841_),
    .A2(_10844_),
    .B(net20643),
    .ZN(_10845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19754_ (.A1(_10838_),
    .A2(_10845_),
    .ZN(_10846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19755_ (.A1(_10746_),
    .A2(_10771_),
    .ZN(_10847_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19756_ (.A1(_10847_),
    .A2(net19840),
    .Z(_10848_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19757_ (.A1(_10717_),
    .A2(_10494_),
    .Z(_10849_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19758_ (.A1(net19413),
    .A2(net19869),
    .A3(_10849_),
    .Z(_10850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19759_ (.A1(_10848_),
    .A2(_10741_),
    .A3(_10850_),
    .ZN(_10851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19760_ (.A1(_10652_),
    .A2(net19413),
    .ZN(_10852_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19761_ (.A1(_10852_),
    .A2(net19864),
    .Z(_10853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19762_ (.A1(_10656_),
    .A2(net17970),
    .ZN(_10854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19763_ (.A1(_10854_),
    .A2(_10853_),
    .B(net20058),
    .ZN(_10855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19764_ (.A1(_10855_),
    .A2(_10851_),
    .ZN(_10856_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19765_ (.A1(_15703_[0]),
    .A2(net19412),
    .B(net19860),
    .ZN(_10857_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19766_ (.A1(_10857_),
    .A2(_10792_),
    .B(net19854),
    .ZN(_10858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19767_ (.A1(_10684_),
    .A2(net19416),
    .ZN(_10859_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19768_ (.A1(net19413),
    .A2(_15694_[0]),
    .Z(_10860_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19769_ (.A1(_10859_),
    .A2(net19860),
    .A3(_10860_),
    .ZN(_10861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19770_ (.A1(_10858_),
    .A2(_10861_),
    .ZN(_10862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19771_ (.A1(_10856_),
    .A2(_10862_),
    .A3(net20644),
    .ZN(_10863_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19772_ (.A1(_10846_),
    .A2(_10863_),
    .A3(_10643_),
    .ZN(_10864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19773_ (.A1(_10830_),
    .A2(_10864_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19774_ (.A1(_10669_),
    .A2(_10595_),
    .ZN(_10865_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19775_ (.A1(_10865_),
    .A2(_10532_),
    .Z(_10866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19776_ (.A1(net19400),
    .A2(net19868),
    .Z(_10867_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19777_ (.I(net18924),
    .ZN(_10868_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19778_ (.A1(_10866_),
    .A2(_10868_),
    .B(_10590_),
    .ZN(_10869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19779_ (.A1(_10648_),
    .A2(net17967),
    .ZN(_10870_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19780_ (.A1(_10779_),
    .A2(_10870_),
    .A3(net19842),
    .ZN(_10871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19781_ (.A1(_10869_),
    .A2(_10871_),
    .B(net19856),
    .ZN(_10872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19782_ (.A1(_10663_),
    .A2(_10669_),
    .ZN(_10873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19783_ (.A1(_10656_),
    .A2(net18928),
    .ZN(_10874_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19784_ (.A1(_10873_),
    .A2(net19865),
    .A3(_10874_),
    .ZN(_10875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19785_ (.A1(_10689_),
    .A2(net18928),
    .ZN(_10876_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19786_ (.I(_10650_),
    .ZN(_10877_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19787_ (.A1(_10876_),
    .A2(net19845),
    .A3(_10877_),
    .ZN(_10878_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19788_ (.A1(_10875_),
    .A2(_10878_),
    .A3(net20643),
    .ZN(_10879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19789_ (.A1(_10879_),
    .A2(_10872_),
    .B(net20642),
    .ZN(_10880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19790_ (.A1(_10497_),
    .A2(_10672_),
    .Z(_10881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19791_ (.A1(_10842_),
    .A2(_10881_),
    .ZN(_10882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19792_ (.A1(_10882_),
    .A2(net19865),
    .ZN(_10883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19793_ (.A1(_10775_),
    .A2(_10703_),
    .A3(_10688_),
    .Z(_10884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19794_ (.A1(_10883_),
    .A2(_10884_),
    .ZN(_10885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19795_ (.A1(_10676_),
    .A2(net17965),
    .ZN(_10886_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _19796_ (.A1(_10886_),
    .A2(net19847),
    .A3(_10670_),
    .Z(_10887_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19797_ (.A1(_10885_),
    .A2(_10887_),
    .B(_10631_),
    .ZN(_10888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19798_ (.A1(net17952),
    .A2(_10819_),
    .B(_10800_),
    .ZN(_10889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19799_ (.A1(_10889_),
    .A2(net19861),
    .ZN(_10890_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19800_ (.A1(_10881_),
    .A2(net19406),
    .Z(_10891_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19801_ (.A1(_10867_),
    .A2(net18351),
    .B(net19865),
    .ZN(_10892_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19802_ (.A1(_10746_),
    .A2(net18345),
    .Z(_10893_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19803_ (.I(_10893_),
    .ZN(_10894_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19804_ (.A1(_10891_),
    .A2(_10892_),
    .A3(_10894_),
    .ZN(_10895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19805_ (.A1(_10890_),
    .A2(_10895_),
    .A3(net20643),
    .ZN(_10896_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19806_ (.A1(_10888_),
    .A2(_10896_),
    .A3(net19854),
    .ZN(_10897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19807_ (.A1(_10880_),
    .A2(_10897_),
    .ZN(_10898_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19808_ (.A1(_10576_),
    .A2(_10446_),
    .Z(_10899_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19809_ (.A1(_10899_),
    .A2(_10893_),
    .B(net20054),
    .ZN(_10900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19810_ (.A1(_10767_),
    .A2(net19413),
    .Z(_10901_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _19811_ (.A1(_10901_),
    .A2(net19854),
    .B1(net19406),
    .B2(net18348),
    .ZN(_10902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19812_ (.A1(_10900_),
    .A2(_10902_),
    .ZN(_10903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19813_ (.A1(_10903_),
    .A2(net19840),
    .ZN(_10904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19814_ (.I(_10625_),
    .ZN(_10905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19815_ (.A1(_10905_),
    .A2(net19411),
    .ZN(_10906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19816_ (.A1(_10906_),
    .A2(_10556_),
    .Z(_10907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19817_ (.A1(_10907_),
    .A2(_10814_),
    .B(net19840),
    .ZN(_10908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19818_ (.A1(_10712_),
    .A2(net498),
    .ZN(_10909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _19819_ (.A1(net19867),
    .A2(_10849_),
    .ZN(_10910_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19820_ (.A1(net17953),
    .A2(_10910_),
    .A3(net19400),
    .ZN(_10911_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19821_ (.A1(_10909_),
    .A2(_10911_),
    .A3(net20055),
    .ZN(_10912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19822_ (.A1(_10908_),
    .A2(_10912_),
    .B(_10631_),
    .ZN(_10913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19823_ (.A1(_10904_),
    .A2(_10913_),
    .ZN(_10914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19824_ (.A1(_10562_),
    .A2(_10910_),
    .ZN(_10915_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19825_ (.A1(_10741_),
    .A2(_10915_),
    .A3(net19861),
    .ZN(_10916_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19826_ (.I(_10809_),
    .ZN(_10917_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19827_ (.A1(_10917_),
    .A2(net19840),
    .B(net19857),
    .ZN(_10918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19828_ (.A1(_10916_),
    .A2(_10918_),
    .B(net20644),
    .ZN(_10919_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19829_ (.A1(_10906_),
    .A2(net19840),
    .Z(_10920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19830_ (.A1(_10676_),
    .A2(net17953),
    .ZN(_10921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19831_ (.A1(net18926),
    .A2(net19425),
    .ZN(_10922_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19832_ (.A1(_10920_),
    .A2(_10921_),
    .A3(_10922_),
    .ZN(_10923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19833_ (.A1(_10750_),
    .A2(net19864),
    .A3(_10506_),
    .ZN(_10924_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19834_ (.A1(_10923_),
    .A2(_10924_),
    .A3(net19854),
    .ZN(_10925_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19835_ (.A1(_10919_),
    .A2(_10925_),
    .ZN(_10926_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19836_ (.A1(_10914_),
    .A2(_10926_),
    .A3(net20642),
    .ZN(_10927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19837_ (.A1(_10898_),
    .A2(_10927_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19838_ (.A1(net18932),
    .A2(net19413),
    .ZN(_10928_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _19839_ (.A1(net19840),
    .A2(_10730_),
    .A3(net17358),
    .A4(_10928_),
    .ZN(_10929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19840_ (.A1(_10663_),
    .A2(net17953),
    .ZN(_10930_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19841_ (.A1(net18927),
    .A2(net19845),
    .ZN(_10931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19842_ (.A1(_10930_),
    .A2(_10931_),
    .B(net19854),
    .ZN(_10932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19843_ (.A1(_10929_),
    .A2(_10932_),
    .ZN(_10933_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19844_ (.A1(_10752_),
    .A2(_10537_),
    .Z(_10934_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19845_ (.A1(_10616_),
    .A2(net19864),
    .A3(_10934_),
    .ZN(_10935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19846_ (.A1(_10718_),
    .A2(net19413),
    .ZN(_10936_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19847_ (.A1(_10936_),
    .A2(net19840),
    .Z(_10937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19848_ (.A1(net18935),
    .A2(net19403),
    .ZN(_10938_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19849_ (.A1(_10937_),
    .A2(_10938_),
    .B(net20059),
    .ZN(_10939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19850_ (.A1(_10935_),
    .A2(_10939_),
    .ZN(_10940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19851_ (.A1(_10933_),
    .A2(_10940_),
    .A3(_10631_),
    .ZN(_10941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19852_ (.A1(_10802_),
    .A2(net19413),
    .ZN(_10942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19853_ (.A1(_10942_),
    .A2(net19840),
    .Z(_10943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19854_ (.A1(_10562_),
    .A2(_10703_),
    .ZN(_10944_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19855_ (.A1(_10703_),
    .A2(net19409),
    .Z(_10945_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19856_ (.A1(_10943_),
    .A2(_10944_),
    .A3(_10945_),
    .ZN(_10946_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19857_ (.I(_15687_[0]),
    .ZN(_10947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19858_ (.A1(_10947_),
    .A2(net19414),
    .B(net19840),
    .ZN(_10948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19859_ (.A1(net18349),
    .A2(net19401),
    .ZN(_10949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19860_ (.A1(_10948_),
    .A2(_10949_),
    .B(net20057),
    .ZN(_10950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19861_ (.A1(_10946_),
    .A2(_10950_),
    .B(_10631_),
    .ZN(_10951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19862_ (.A1(_10729_),
    .A2(net19413),
    .ZN(_10952_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19863_ (.I(_10669_),
    .ZN(_10953_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19864_ (.A1(_10952_),
    .A2(_10953_),
    .ZN(_10954_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19865_ (.I(_10954_),
    .ZN(_10955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19866_ (.A1(net17596),
    .A2(net18940),
    .ZN(_10956_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19867_ (.A1(_10955_),
    .A2(_10956_),
    .A3(net19845),
    .ZN(_10957_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19868_ (.A1(_10609_),
    .A2(net19865),
    .A3(_10670_),
    .ZN(_10958_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19869_ (.A1(_10957_),
    .A2(_10958_),
    .A3(net20059),
    .ZN(_10959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19870_ (.A1(_10951_),
    .A2(_10959_),
    .ZN(_10960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19871_ (.A1(_10941_),
    .A2(net20642),
    .A3(_10960_),
    .ZN(_10961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19872_ (.A1(_10716_),
    .A2(net17955),
    .ZN(_10962_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19873_ (.A1(_10563_),
    .A2(net19864),
    .A3(_10962_),
    .ZN(_10963_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19874_ (.A1(_10536_),
    .A2(net19413),
    .ZN(_10964_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19875_ (.A1(_10964_),
    .A2(net17948),
    .ZN(_10965_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19876_ (.A1(_10763_),
    .A2(_10965_),
    .B(net20058),
    .ZN(_10966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19877_ (.A1(_10963_),
    .A2(_10966_),
    .B(_10631_),
    .ZN(_10967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19878_ (.A1(_10842_),
    .A2(_10448_),
    .ZN(_10968_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19879_ (.A1(_10968_),
    .A2(net19851),
    .A3(_10793_),
    .ZN(_10969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19880_ (.A1(net18937),
    .A2(_10499_),
    .ZN(_10970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19881_ (.A1(_10970_),
    .A2(net19402),
    .B(net19840),
    .ZN(_10971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19882_ (.A1(_10496_),
    .A2(_10971_),
    .ZN(_10972_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19883_ (.A1(_10969_),
    .A2(_10972_),
    .A3(net20058),
    .ZN(_10973_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19884_ (.A1(_10967_),
    .A2(_10973_),
    .B(net20642),
    .ZN(_10974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19885_ (.A1(_10835_),
    .A2(_10737_),
    .ZN(_10975_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19886_ (.A1(net18942),
    .A2(net19406),
    .A3(net17963),
    .Z(_10976_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19887_ (.A1(_10976_),
    .A2(_10954_),
    .B(net19846),
    .ZN(_10977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19888_ (.A1(_10975_),
    .A2(_10977_),
    .A3(net20059),
    .ZN(_10978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19889_ (.I(_10761_),
    .ZN(_10979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19890_ (.A1(_10979_),
    .A2(_10688_),
    .ZN(_10980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19891_ (.A1(_10689_),
    .A2(_10657_),
    .ZN(_10981_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19892_ (.A1(_10980_),
    .A2(net19865),
    .A3(_10981_),
    .ZN(_10982_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _19893_ (.A1(net17596),
    .A2(net19865),
    .A3(net18348),
    .Z(_10983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19894_ (.A1(_10982_),
    .A2(net19854),
    .A3(_10983_),
    .ZN(_10984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19895_ (.A1(_10978_),
    .A2(_10631_),
    .A3(_10984_),
    .ZN(_10985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19896_ (.A1(_10974_),
    .A2(_10985_),
    .ZN(_10986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19897_ (.A1(_10961_),
    .A2(_10986_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19898_ (.A1(_10613_),
    .A2(net18347),
    .ZN(_10987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19899_ (.A1(_10712_),
    .A2(_10771_),
    .ZN(_10988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19900_ (.A1(_10988_),
    .A2(net19843),
    .ZN(_10989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19901_ (.A1(_10987_),
    .A2(net19406),
    .B(_10989_),
    .ZN(_10990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19902_ (.A1(net19408),
    .A2(net19399),
    .ZN(_10991_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19903_ (.A1(_10955_),
    .A2(net19865),
    .A3(_10991_),
    .Z(_10992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19904_ (.A1(_10990_),
    .A2(_10992_),
    .B(net19855),
    .ZN(_10993_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19905_ (.A1(_10936_),
    .A2(net18352),
    .ZN(_10994_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19906_ (.A1(_10994_),
    .A2(_10964_),
    .B(net19849),
    .ZN(_10995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19907_ (.A1(_10808_),
    .A2(net19420),
    .ZN(_10996_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _19908_ (.A1(net17594),
    .A2(_10608_),
    .B(net19865),
    .C(_10996_),
    .ZN(_10997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19909_ (.A1(_10995_),
    .A2(_10997_),
    .ZN(_10998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19910_ (.A1(_10998_),
    .A2(net20060),
    .B(_10631_),
    .ZN(_10999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19911_ (.A1(_10993_),
    .A2(_10999_),
    .ZN(_11000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _19912_ (.A1(_10746_),
    .A2(net497),
    .B(net19840),
    .ZN(_11001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19913_ (.I(_10676_),
    .ZN(_11002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19914_ (.A1(_11001_),
    .A2(_11002_),
    .A3(net17591),
    .ZN(_11003_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19915_ (.A1(_10752_),
    .A2(net19840),
    .Z(_11004_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19916_ (.A1(_11004_),
    .A2(_10747_),
    .B(net19854),
    .ZN(_11005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19917_ (.A1(_11003_),
    .A2(_11005_),
    .B(net20643),
    .ZN(_11006_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19918_ (.A1(_10561_),
    .A2(net19412),
    .Z(_11007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19919_ (.A1(_10448_),
    .A2(_11007_),
    .ZN(_11008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19920_ (.A1(net19402),
    .A2(net18424),
    .ZN(_11009_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19921_ (.A1(_10574_),
    .A2(_11008_),
    .A3(_11009_),
    .ZN(_11010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19922_ (.A1(_10693_),
    .A2(net17964),
    .ZN(_11011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19923_ (.A1(_10701_),
    .A2(_11011_),
    .ZN(_11012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19924_ (.A1(_11010_),
    .A2(_11012_),
    .A3(net19859),
    .ZN(_11013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19925_ (.A1(_11006_),
    .A2(_11013_),
    .B(net20642),
    .ZN(_11014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19926_ (.A1(_11000_),
    .A2(_11014_),
    .ZN(_11015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19927_ (.I(_10613_),
    .ZN(_11016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19928_ (.A1(_10910_),
    .A2(net19410),
    .ZN(_11017_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _19929_ (.A1(_11016_),
    .A2(_10859_),
    .B(net19864),
    .C(_11017_),
    .ZN(_11018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19930_ (.I(_10693_),
    .ZN(_11019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19931_ (.A1(_10763_),
    .A2(_11019_),
    .B(net20058),
    .ZN(_11020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19932_ (.A1(_11018_),
    .A2(_11020_),
    .ZN(_11021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19933_ (.A1(_10656_),
    .A2(net18347),
    .ZN(_11022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19934_ (.A1(_10648_),
    .A2(net17953),
    .ZN(_11023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19935_ (.A1(_11022_),
    .A2(_11023_),
    .A3(net19844),
    .ZN(_11024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19936_ (.A1(net17961),
    .A2(net19419),
    .ZN(_11025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19937_ (.A1(net18346),
    .A2(net19406),
    .B(net19840),
    .ZN(_11026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19938_ (.A1(_11025_),
    .A2(_11026_),
    .ZN(_11027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19939_ (.A1(_11024_),
    .A2(_11027_),
    .A3(net20060),
    .ZN(_11028_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19940_ (.A1(_11021_),
    .A2(_11028_),
    .A3(net20643),
    .ZN(_11029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19941_ (.A1(net19428),
    .A2(net19406),
    .B(net19840),
    .ZN(_11030_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19942_ (.A1(_11030_),
    .A2(_10667_),
    .B(net20059),
    .ZN(_11031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19943_ (.A1(_10656_),
    .A2(_10684_),
    .ZN(_11032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19944_ (.A1(_11007_),
    .A2(_10703_),
    .ZN(_11033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19945_ (.A1(_11032_),
    .A2(_11033_),
    .A3(net19844),
    .ZN(_11034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19946_ (.A1(_11034_),
    .A2(_11031_),
    .B(net20643),
    .ZN(_11035_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19947_ (.A1(net17962),
    .A2(net19421),
    .A3(net17953),
    .ZN(_11036_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19948_ (.A1(_10653_),
    .A2(net19408),
    .B(net19865),
    .ZN(_11037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19949_ (.A1(_11036_),
    .A2(_11037_),
    .B(net19854),
    .ZN(_11038_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19950_ (.A1(_10616_),
    .A2(_10619_),
    .A3(net17947),
    .ZN(_11039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19951_ (.A1(_11038_),
    .A2(_11039_),
    .ZN(_11040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19952_ (.A1(_11035_),
    .A2(_11040_),
    .ZN(_11041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19953_ (.A1(_11029_),
    .A2(_11041_),
    .A3(net20642),
    .ZN(_11042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19954_ (.A1(_11015_),
    .A2(_11042_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19955_ (.A1(_11007_),
    .A2(_10706_),
    .ZN(_11043_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19956_ (.A1(_11043_),
    .A2(_10847_),
    .A3(_10569_),
    .ZN(_11044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19957_ (.A1(_11044_),
    .A2(net19860),
    .Z(_11045_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19958_ (.A1(_10626_),
    .A2(_10801_),
    .Z(_11046_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _19959_ (.A1(_10539_),
    .A2(_11046_),
    .A3(_10942_),
    .Z(_11047_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _19960_ (.A1(_11047_),
    .A2(_11045_),
    .B(net20056),
    .ZN(_11048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19961_ (.A1(_10508_),
    .A2(net19402),
    .ZN(_11049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _19962_ (.A1(_10852_),
    .A2(_11049_),
    .Z(_11050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19963_ (.A1(_11050_),
    .A2(_10920_),
    .B(net20059),
    .ZN(_11051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19964_ (.A1(_10842_),
    .A2(_10669_),
    .ZN(_11052_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _19965_ (.A1(_15692_[0]),
    .A2(_15701_[0]),
    .B(net19417),
    .ZN(_11053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19966_ (.A1(_11052_),
    .A2(net19865),
    .A3(_11053_),
    .ZN(_11054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19967_ (.A1(_11051_),
    .A2(_11054_),
    .B(net20643),
    .ZN(_11055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19968_ (.A1(_11055_),
    .A2(_11048_),
    .ZN(_11056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19969_ (.A1(_10979_),
    .A2(_10669_),
    .ZN(_11057_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19970_ (.A1(_10653_),
    .A2(net19413),
    .B(net19865),
    .ZN(_11058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19971_ (.A1(_11057_),
    .A2(_11058_),
    .B(net19854),
    .ZN(_11059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19972_ (.A1(_10775_),
    .A2(_10910_),
    .ZN(_11060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19973_ (.A1(_11001_),
    .A2(_10670_),
    .A3(_11060_),
    .ZN(_11061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19974_ (.A1(_11059_),
    .A2(_11061_),
    .B(_10631_),
    .ZN(_11062_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19975_ (.A1(_10684_),
    .A2(net19416),
    .A3(net17958),
    .ZN(_11063_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19976_ (.A1(_11063_),
    .A2(net19841),
    .A3(_10860_),
    .ZN(_11064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19977_ (.A1(_10684_),
    .A2(net19404),
    .A3(_10703_),
    .ZN(_11065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19978_ (.A1(net17949),
    .A2(net18343),
    .A3(net19416),
    .ZN(_11066_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19979_ (.A1(_11065_),
    .A2(_11066_),
    .A3(net19860),
    .ZN(_11067_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19980_ (.A1(_11064_),
    .A2(_11067_),
    .A3(net19857),
    .ZN(_11068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19981_ (.A1(_11062_),
    .A2(_11068_),
    .ZN(_11069_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19982_ (.A1(_11069_),
    .A2(_11056_),
    .A3(_10643_),
    .ZN(_11070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19983_ (.I(_10576_),
    .ZN(_11071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19984_ (.A1(_10944_),
    .A2(_11071_),
    .ZN(_11072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19985_ (.A1(_11072_),
    .A2(net19841),
    .ZN(_11073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19986_ (.A1(_10790_),
    .A2(net19860),
    .ZN(_11074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19987_ (.A1(_11073_),
    .A2(_11074_),
    .ZN(_11075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19988_ (.A1(_11075_),
    .A2(net20053),
    .ZN(_11076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19989_ (.A1(_10693_),
    .A2(net18343),
    .ZN(_11077_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19990_ (.A1(_11077_),
    .A2(net19851),
    .A3(_10724_),
    .ZN(_11078_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19991_ (.I(_15693_[0]),
    .ZN(_11079_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19992_ (.A1(_11079_),
    .A2(net19406),
    .B(net19840),
    .ZN(_11080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19993_ (.A1(_11080_),
    .A2(_11033_),
    .ZN(_11081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19994_ (.A1(_11078_),
    .A2(_11081_),
    .A3(net19856),
    .ZN(_11082_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19995_ (.A1(_11076_),
    .A2(_11082_),
    .A3(net20644),
    .ZN(_11083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19996_ (.A1(net18342),
    .A2(net19849),
    .A3(_10690_),
    .ZN(_11084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19997_ (.A1(_10811_),
    .A2(net17956),
    .ZN(_11085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _19998_ (.A1(_11001_),
    .A2(_11085_),
    .ZN(_11086_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _19999_ (.A1(_11084_),
    .A2(_11086_),
    .A3(net20053),
    .ZN(_11087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20000_ (.A1(net19412),
    .A2(net19399),
    .ZN(_11088_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20001_ (.A1(_10866_),
    .A2(net18923),
    .B(net20053),
    .ZN(_11089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20002_ (.A1(_10716_),
    .A2(net18941),
    .ZN(_11090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20003_ (.A1(_10865_),
    .A2(net19405),
    .ZN(_11091_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20004_ (.A1(_11090_),
    .A2(_11091_),
    .A3(net19840),
    .ZN(_11092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20005_ (.A1(_11089_),
    .A2(_11092_),
    .ZN(_11093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20006_ (.A1(_11087_),
    .A2(_11093_),
    .A3(_10631_),
    .ZN(_11094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20007_ (.A1(_11083_),
    .A2(_11094_),
    .A3(net20642),
    .ZN(_11095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20008_ (.A1(_11095_),
    .A2(_11070_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20009_ (.A1(_10532_),
    .A2(_10499_),
    .Z(_11096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20010_ (.A1(_11096_),
    .A2(_10510_),
    .Z(_11097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20011_ (.A1(net18932),
    .A2(net19402),
    .ZN(_11098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20012_ (.A1(_11097_),
    .A2(_11098_),
    .B(net19857),
    .ZN(_11099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20013_ (.A1(net19414),
    .A2(net18424),
    .ZN(_11100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20014_ (.A1(_11052_),
    .A2(net19853),
    .A3(_11100_),
    .ZN(_11101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20015_ (.A1(_11099_),
    .A2(_11101_),
    .B(net20643),
    .ZN(_11102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20016_ (.I(_10615_),
    .ZN(_11103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20017_ (.A1(net499),
    .A2(_10597_),
    .ZN(_11104_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20018_ (.A1(net18341),
    .A2(_10952_),
    .B1(_11104_),
    .B2(net19421),
    .ZN(_11105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20019_ (.A1(_11105_),
    .A2(_10853_),
    .ZN(_11106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20020_ (.A1(_11088_),
    .A2(_10572_),
    .Z(_11107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20021_ (.A1(_11103_),
    .A2(net19422),
    .ZN(_11108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20022_ (.A1(_11107_),
    .A2(_11108_),
    .Z(_11109_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20023_ (.A1(_11109_),
    .A2(_10915_),
    .B(net20059),
    .ZN(_11110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20024_ (.A1(_11106_),
    .A2(_11110_),
    .ZN(_11111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20025_ (.A1(_11102_),
    .A2(_11111_),
    .ZN(_11112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20026_ (.A1(_10712_),
    .A2(_10703_),
    .ZN(_11113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20027_ (.A1(_10650_),
    .A2(net18343),
    .ZN(_11114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20028_ (.A1(_11113_),
    .A2(_11114_),
    .A3(net19840),
    .ZN(_11115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20029_ (.A1(_10649_),
    .A2(_10625_),
    .Z(_11116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20030_ (.A1(net19406),
    .A2(_15701_[0]),
    .ZN(_11117_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20031_ (.A1(_11116_),
    .A2(net19400),
    .B(net19861),
    .C(_11117_),
    .ZN(_11118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20032_ (.A1(_11115_),
    .A2(_11118_),
    .A3(net20055),
    .ZN(_11119_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20033_ (.A1(net18421),
    .A2(net19414),
    .B(_10510_),
    .C(net19862),
    .ZN(_11120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20034_ (.A1(_10730_),
    .A2(net17947),
    .A3(_11107_),
    .ZN(_11121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20035_ (.A1(_11120_),
    .A2(_11121_),
    .A3(net19854),
    .ZN(_11122_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20036_ (.A1(_11119_),
    .A2(_11122_),
    .A3(net20643),
    .ZN(_11123_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20037_ (.A1(_11112_),
    .A2(_11123_),
    .A3(_10643_),
    .ZN(_11124_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20038_ (.A1(_10448_),
    .A2(net19406),
    .B(net19865),
    .ZN(_11125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20039_ (.A1(_10648_),
    .A2(net18935),
    .ZN(_11126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20040_ (.A1(_11125_),
    .A2(_11126_),
    .B(net19854),
    .ZN(_11127_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20041_ (.A1(_10867_),
    .A2(_10771_),
    .Z(_11128_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20042_ (.A1(_10901_),
    .A2(net19840),
    .A3(_11128_),
    .Z(_11129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20043_ (.A1(_11129_),
    .A2(_11127_),
    .B(_10631_),
    .ZN(_11130_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20044_ (.A1(net19428),
    .A2(net19406),
    .B(_10980_),
    .ZN(_11131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20045_ (.A1(_11131_),
    .A2(net19843),
    .ZN(_11132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20046_ (.A1(net18935),
    .A2(net19418),
    .A3(_10703_),
    .ZN(_11133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20047_ (.A1(_10835_),
    .A2(_11133_),
    .ZN(_11134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20048_ (.A1(_11132_),
    .A2(_11134_),
    .A3(net19855),
    .ZN(_11135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20049_ (.A1(_11135_),
    .A2(_11130_),
    .ZN(_11136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20050_ (.A1(_10448_),
    .A2(_10712_),
    .ZN(_11137_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20051_ (.A1(_10892_),
    .A2(_11137_),
    .A3(_10847_),
    .ZN(_11138_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20052_ (.A1(_10716_),
    .A2(net19840),
    .ZN(_11139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20053_ (.A1(_11139_),
    .A2(_10944_),
    .B(net20055),
    .ZN(_11140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20054_ (.A1(_11138_),
    .A2(_11140_),
    .B(net20643),
    .ZN(_11141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20055_ (.A1(_10843_),
    .A2(net19861),
    .A3(_11043_),
    .ZN(_11142_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20056_ (.A1(_10909_),
    .A2(_10758_),
    .A3(net19848),
    .ZN(_11143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20057_ (.A1(_11142_),
    .A2(_11143_),
    .A3(net20055),
    .ZN(_11144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20058_ (.A1(_11141_),
    .A2(_11144_),
    .B(_10643_),
    .ZN(_11145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20059_ (.A1(_11145_),
    .A2(_11136_),
    .ZN(_11146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20060_ (.A1(_11146_),
    .A2(_11124_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20061_ (.A1(\sa21_sr[1] ),
    .A2(\sa30_sub[1] ),
    .Z(_11147_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20062_ (.I(\sa01_sr[7] ),
    .ZN(_11148_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20063_ (.I(\sa01_sr[0] ),
    .ZN(_11149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20064_ (.A1(_11148_),
    .A2(_11149_),
    .ZN(_11150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20065_ (.A1(net21458),
    .A2(net21469),
    .ZN(_11151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20066_ (.A1(_11150_),
    .A2(_11151_),
    .ZN(_11152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20067_ (.A1(_11147_),
    .A2(_11152_),
    .ZN(_11153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20068_ (.A1(_11149_),
    .A2(net21458),
    .ZN(_11154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20069_ (.A1(_11148_),
    .A2(net21469),
    .ZN(_11155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20070_ (.A1(_11154_),
    .A2(_11155_),
    .ZN(_11156_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20071_ (.I(\sa21_sr[1] ),
    .ZN(_11157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20072_ (.I(\sa30_sub[1] ),
    .ZN(_11158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20073_ (.A1(_11158_),
    .A2(_11157_),
    .ZN(_11159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20074_ (.A1(\sa21_sr[1] ),
    .A2(\sa30_sub[1] ),
    .ZN(_11160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20075_ (.A1(_11159_),
    .A2(_11160_),
    .ZN(_11161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20076_ (.A1(_11156_),
    .A2(_11161_),
    .ZN(_11162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20077_ (.A1(_11153_),
    .A2(_11162_),
    .ZN(_11163_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20078_ (.I(_11163_),
    .ZN(_11164_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20079_ (.I(\sa11_sr[7] ),
    .ZN(_11165_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20080_ (.I(\sa11_sr[0] ),
    .ZN(_11166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20081_ (.A1(_11165_),
    .A2(_11166_),
    .ZN(_11167_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17538 (.I(_13710_),
    .Z(net17538));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20083_ (.A1(net21400),
    .A2(\sa11_sr[0] ),
    .ZN(_11169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20084_ (.A1(_11167_),
    .A2(_11169_),
    .ZN(_11170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20085_ (.A1(_11170_),
    .A2(net21409),
    .ZN(_11171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20086_ (.A1(_11166_),
    .A2(\sa11_sr[7] ),
    .ZN(_11172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20087_ (.A1(_11165_),
    .A2(\sa11_sr[0] ),
    .ZN(_11173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20088_ (.A1(_11172_),
    .A2(_11173_),
    .ZN(_11174_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20089_ (.I(\sa11_sr[1] ),
    .ZN(_11175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20090_ (.A1(_11174_),
    .A2(_11175_),
    .ZN(_11176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20091_ (.A1(_11171_),
    .A2(_11176_),
    .ZN(_11177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20092_ (.I(_11177_),
    .ZN(_11178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20093_ (.A1(_11164_),
    .A2(_11178_),
    .ZN(_11179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20094_ (.A1(_11163_),
    .A2(_11177_),
    .ZN(_11180_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20095_ (.A1(_11179_),
    .A2(_10378_),
    .A3(_11180_),
    .ZN(_11181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20096_ (.A1(net21493),
    .A2(\text_in_r[89] ),
    .ZN(_11182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20097_ (.A1(_11181_),
    .A2(_11182_),
    .ZN(_11183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20098_ (.A1(net19839),
    .A2(_07913_),
    .ZN(_11184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20099_ (.A1(_11181_),
    .A2(net21194),
    .A3(_11182_),
    .ZN(_11185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20100_ (.A1(_11184_),
    .A2(_11185_),
    .ZN(_11186_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17502 (.I(_00907_),
    .Z(net17502));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20102_ (.A1(_11148_),
    .A2(_11165_),
    .ZN(_11187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20103_ (.A1(net21458),
    .A2(net21401),
    .ZN(_11188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20104_ (.A1(_11187_),
    .A2(_11188_),
    .ZN(_11189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20105_ (.I(\sa30_sub[0] ),
    .ZN(_11190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20106_ (.A1(_11189_),
    .A2(net21042),
    .ZN(_11191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20107_ (.A1(net20954),
    .A2(net21297),
    .A3(_11188_),
    .ZN(_11192_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20108_ (.A1(net21043),
    .A2(net21360),
    .ZN(_11193_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20109_ (.I(\sa21_sr[0] ),
    .ZN(_11194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20110_ (.A1(net21041),
    .A2(net21411),
    .ZN(_11195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20111_ (.A1(_11193_),
    .A2(_11195_),
    .ZN(_11196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20112_ (.A1(_11191_),
    .A2(_11192_),
    .A3(_11196_),
    .ZN(_11197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20113_ (.A1(_11189_),
    .A2(net21297),
    .ZN(_11198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20114_ (.A1(net20954),
    .A2(net21042),
    .A3(_11188_),
    .ZN(_11199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20115_ (.I(_11196_),
    .ZN(_11200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20116_ (.A1(_11198_),
    .A2(_11199_),
    .A3(_11200_),
    .ZN(_11201_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17516 (.I(_15213_),
    .Z(net17516));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17526 (.I(_14468_),
    .Z(net17526));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20119_ (.A1(_11197_),
    .A2(_11201_),
    .B(net21493),
    .ZN(_11204_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20120_ (.I(\text_in_r[88] ),
    .ZN(_11205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20121_ (.A1(_11205_),
    .A2(net21493),
    .Z(_11206_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20122_ (.A1(net20445),
    .A2(net20953),
    .B(net21195),
    .ZN(_11207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20123_ (.A1(_11197_),
    .A2(_11201_),
    .ZN(_11208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20124_ (.A1(_11208_),
    .A2(net21073),
    .ZN(_11209_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20125_ (.I(_11206_),
    .ZN(_11210_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20126_ (.A1(net20279),
    .A2(_07908_),
    .A3(net20907),
    .ZN(_11211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20127_ (.A1(_11207_),
    .A2(_11211_),
    .ZN(_15714_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20128_ (.I(\sa01_sr[1] ),
    .ZN(_11212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20129_ (.A1(_11175_),
    .A2(_11212_),
    .ZN(_11213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20130_ (.A1(\sa11_sr[1] ),
    .A2(\sa01_sr[1] ),
    .ZN(_11214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20131_ (.A1(_11213_),
    .A2(_11214_),
    .ZN(_11215_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20132_ (.I(\sa21_sr[2] ),
    .ZN(_11216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20133_ (.A1(net20906),
    .A2(net21038),
    .ZN(_11217_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17493 (.I(_01094_),
    .Z(net17493));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20135_ (.A1(net20952),
    .A2(net21355),
    .A3(net21039),
    .ZN(_11219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20136_ (.A1(_11217_),
    .A2(_11219_),
    .ZN(_11220_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20137_ (.I(\sa30_sub[2] ),
    .ZN(_11221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20138_ (.A1(_11221_),
    .A2(\sa11_sr[2] ),
    .ZN(_11222_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20139_ (.I(\sa11_sr[2] ),
    .ZN(_11223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20140_ (.A1(_11223_),
    .A2(net21292),
    .ZN(_11224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20141_ (.A1(_11222_),
    .A2(_11224_),
    .ZN(_11225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20142_ (.I(_11225_),
    .ZN(_11226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20143_ (.A1(_11220_),
    .A2(_11226_),
    .ZN(_11227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20144_ (.A1(_11217_),
    .A2(_11219_),
    .A3(_11225_),
    .ZN(_11228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20145_ (.A1(_11227_),
    .A2(_11228_),
    .B(net21499),
    .ZN(_11229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20146_ (.I(\text_in_r[90] ),
    .ZN(_11230_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20147_ (.A1(_11230_),
    .A2(net21499),
    .Z(_11231_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20148_ (.A1(_11229_),
    .A2(_11231_),
    .B(_07917_),
    .ZN(_11232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20149_ (.A1(_11227_),
    .A2(_11228_),
    .ZN(_11233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20150_ (.A1(_11233_),
    .A2(net21073),
    .ZN(_11234_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20151_ (.I(_11231_),
    .ZN(_11235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20152_ (.A1(_11234_),
    .A2(net21193),
    .A3(_11235_),
    .ZN(_11236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20153_ (.A1(_11232_),
    .A2(_11236_),
    .ZN(_11237_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17485 (.I(_01348_),
    .Z(net17485));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17479 (.I(_01730_),
    .Z(net17479));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20156_ (.A1(_11204_),
    .A2(_11206_),
    .B(_07908_),
    .ZN(_11239_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20157_ (.A1(_11209_),
    .A2(net21195),
    .A3(_11210_),
    .ZN(_11240_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20158_ (.A1(_11239_),
    .A2(_11240_),
    .ZN(_15705_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20159_ (.A1(_11229_),
    .A2(_11231_),
    .B(net21193),
    .ZN(_11241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20160_ (.A1(_11234_),
    .A2(_07917_),
    .A3(_11235_),
    .ZN(_11242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20161_ (.A1(_11241_),
    .A2(_11242_),
    .ZN(_11243_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17496 (.I(_01062_),
    .Z(net17496));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20163_ (.I(_15715_[0]),
    .ZN(_11244_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20164_ (.A1(net19396),
    .A2(_11244_),
    .Z(_11245_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20165_ (.I(_15707_[0]),
    .ZN(_11246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20166_ (.A1(net20051),
    .A2(net19836),
    .A3(_11246_),
    .ZN(_11247_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20167_ (.I(_11247_),
    .ZN(_11248_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20168_ (.A1(\sa21_sr[3] ),
    .A2(\sa30_sub[3] ),
    .Z(_11249_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20169_ (.I(\sa01_sr[2] ),
    .ZN(_11250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20170_ (.A1(net21048),
    .A2(_11250_),
    .ZN(_11251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20171_ (.A1(net21459),
    .A2(net21464),
    .ZN(_11252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20172_ (.A1(_11251_),
    .A2(_11252_),
    .ZN(_11253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20173_ (.A1(_11249_),
    .A2(_11253_),
    .ZN(_11254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20174_ (.A1(net21035),
    .A2(net21459),
    .ZN(_11255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20175_ (.A1(net21048),
    .A2(net21464),
    .ZN(_11256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20176_ (.A1(_11255_),
    .A2(_11256_),
    .ZN(_11257_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20177_ (.I(\sa21_sr[3] ),
    .ZN(_11258_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20178_ (.I(\sa30_sub[3] ),
    .ZN(_11259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20179_ (.A1(_11258_),
    .A2(_11259_),
    .ZN(_11260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20180_ (.A1(net21353),
    .A2(\sa30_sub[3] ),
    .ZN(_11261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20181_ (.A1(_11260_),
    .A2(_11261_),
    .ZN(_11262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20182_ (.A1(_11257_),
    .A2(_11262_),
    .ZN(_11263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20183_ (.A1(_11254_),
    .A2(_11263_),
    .ZN(_11264_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20184_ (.I(_11264_),
    .ZN(_11265_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20185_ (.I(\sa11_sr[3] ),
    .ZN(_11266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20186_ (.A1(net21033),
    .A2(net21402),
    .ZN(_11267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20187_ (.A1(net21044),
    .A2(net21407),
    .ZN(_11268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20188_ (.A1(_11267_),
    .A2(_11268_),
    .ZN(_11269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20189_ (.A1(_11269_),
    .A2(net21408),
    .ZN(_11270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20190_ (.A1(net21044),
    .A2(_11266_),
    .ZN(_11271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20191_ (.A1(net21402),
    .A2(net21407),
    .ZN(_11272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20192_ (.A1(_11271_),
    .A2(_11272_),
    .ZN(_11273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20193_ (.A1(_11273_),
    .A2(net21037),
    .ZN(_11274_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20194_ (.A1(_11270_),
    .A2(_11274_),
    .ZN(_11275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20195_ (.A1(_11265_),
    .A2(_11275_),
    .ZN(_11276_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20196_ (.I(_11275_),
    .ZN(_11277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20197_ (.A1(_11277_),
    .A2(_11264_),
    .ZN(_11278_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17482 (.I(_01718_),
    .Z(net17482));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20199_ (.A1(_11276_),
    .A2(_11278_),
    .A3(net21070),
    .ZN(_11280_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20200_ (.A1(net21503),
    .A2(\text_in_r[91] ),
    .ZN(_11281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20201_ (.A1(_11280_),
    .A2(_07921_),
    .A3(_11281_),
    .ZN(_11282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20202_ (.A1(_11265_),
    .A2(_11277_),
    .ZN(_11283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20203_ (.A1(_11264_),
    .A2(_11275_),
    .ZN(_11284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20204_ (.A1(_11283_),
    .A2(net21070),
    .A3(_11284_),
    .ZN(_11285_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20205_ (.A1(net21070),
    .A2(\text_in_r[91] ),
    .Z(_11286_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20206_ (.A1(_11285_),
    .A2(net21192),
    .A3(_11286_),
    .ZN(_11287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20207_ (.A1(_11282_),
    .A2(_11287_),
    .ZN(_11288_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17512 (.I(_15227_),
    .Z(net17512));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17533 (.I(_13812_),
    .Z(net17533));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20210_ (.A1(_11245_),
    .A2(_11248_),
    .B(net19380),
    .ZN(_11291_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20211_ (.I(_15708_[0]),
    .ZN(_11292_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20212_ (.A1(net20051),
    .A2(net19836),
    .A3(_11292_),
    .ZN(_11293_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20213_ (.A1(_11280_),
    .A2(net21192),
    .A3(_11281_),
    .ZN(_11294_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20214_ (.A1(_11285_),
    .A2(_07921_),
    .A3(_11286_),
    .ZN(_11295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20215_ (.A1(_11294_),
    .A2(_11295_),
    .ZN(_11296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20216_ (.A1(net19363),
    .A2(_11293_),
    .ZN(_11297_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20217_ (.I(_11297_),
    .ZN(_11298_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20218_ (.A1(net20050),
    .A2(net19833),
    .A3(net18004),
    .ZN(_11299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20219_ (.A1(_11298_),
    .A2(_11299_),
    .ZN(_11300_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20220_ (.A1(net21459),
    .A2(net21462),
    .Z(_11301_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20221_ (.A1(\sa21_sr[4] ),
    .A2(\sa30_sub[4] ),
    .Z(_11302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20222_ (.A1(\sa21_sr[4] ),
    .A2(\sa30_sub[4] ),
    .ZN(_11303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20223_ (.A1(_11302_),
    .A2(_11303_),
    .ZN(_11304_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20224_ (.I(_11304_),
    .ZN(_11305_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20225_ (.A1(_11301_),
    .A2(_11305_),
    .Z(_11306_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20226_ (.A1(net21406),
    .A2(_11273_),
    .Z(_11307_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20227_ (.I(_11307_),
    .ZN(_11308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20228_ (.A1(_11306_),
    .A2(_11308_),
    .ZN(_11309_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20229_ (.A1(net20951),
    .A2(_11301_),
    .Z(_11310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20230_ (.A1(_11310_),
    .A2(_11307_),
    .ZN(_11311_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20231_ (.A1(_11309_),
    .A2(_11311_),
    .A3(net21069),
    .ZN(_11312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20232_ (.A1(net21505),
    .A2(\text_in_r[92] ),
    .ZN(_11313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20233_ (.A1(_11312_),
    .A2(_11313_),
    .ZN(_11314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20234_ (.A1(_11314_),
    .A2(net21191),
    .ZN(_11315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20235_ (.A1(_11312_),
    .A2(_07925_),
    .A3(_11313_),
    .ZN(_11316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20236_ (.A1(_11315_),
    .A2(_11316_),
    .ZN(_11317_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17475 (.I(_01750_),
    .Z(net17475));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17469 (.I(_01791_),
    .Z(net17469));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20239_ (.A1(_11291_),
    .A2(_11300_),
    .A3(net19360),
    .ZN(_11320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20240_ (.A1(_11183_),
    .A2(net21194),
    .ZN(_11321_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20241_ (.A1(_11181_),
    .A2(_07913_),
    .A3(_11182_),
    .ZN(_11322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20242_ (.A1(_11322_),
    .A2(_11321_),
    .ZN(_15706_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20243_ (.A1(net18918),
    .A2(net19374),
    .A3(net19395),
    .ZN(_11323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20244_ (.I(_11293_),
    .ZN(_11324_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17468 (.I(_01818_),
    .Z(net17468));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20246_ (.A1(_11324_),
    .A2(net19374),
    .ZN(_11326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20247_ (.A1(net19393),
    .A2(net17944),
    .ZN(_11327_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17465 (.I(_01864_),
    .Z(net17465));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20249_ (.A1(_11327_),
    .A2(net19363),
    .ZN(_11329_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20250_ (.A1(_11323_),
    .A2(_11326_),
    .A3(net17356),
    .ZN(_11330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20251_ (.A1(_11314_),
    .A2(_07925_),
    .ZN(_11331_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20252_ (.A1(_11312_),
    .A2(net21191),
    .A3(_11313_),
    .ZN(_11332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20253_ (.A1(_11331_),
    .A2(_11332_),
    .ZN(_11333_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17473 (.I(_01754_),
    .Z(net17473));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17464 (.I(_01877_),
    .Z(net17464));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20256_ (.A1(_11330_),
    .A2(net19351),
    .ZN(_11336_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20257_ (.A1(\sa21_sr[5] ),
    .A2(\sa30_sub[5] ),
    .Z(_11337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20258_ (.A1(\sa21_sr[5] ),
    .A2(\sa30_sub[5] ),
    .ZN(_11338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20259_ (.A1(_11337_),
    .A2(_11338_),
    .ZN(_11339_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20260_ (.A1(net21405),
    .A2(_11339_),
    .Z(_11340_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20261_ (.A1(\sa11_sr[4] ),
    .A2(\sa01_sr[4] ),
    .Z(_11341_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20262_ (.I(_11341_),
    .ZN(_11342_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20263_ (.A1(_11340_),
    .A2(net20949),
    .Z(_11343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20264_ (.A1(_11340_),
    .A2(net20949),
    .ZN(_11344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20265_ (.A1(_11343_),
    .A2(_11344_),
    .ZN(_11345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20266_ (.A1(net21495),
    .A2(\text_in_r[93] ),
    .ZN(_11346_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20267_ (.A1(_11345_),
    .A2(net21495),
    .B(_07929_),
    .C(_11346_),
    .ZN(_11347_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17463 (.I(_01907_),
    .Z(net17463));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20269_ (.A1(_11343_),
    .A2(net21067),
    .A3(_11344_),
    .ZN(_11349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20270_ (.A1(_11349_),
    .A2(_11346_),
    .ZN(_11350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20271_ (.A1(_11350_),
    .A2(net21190),
    .ZN(_11351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20272_ (.A1(_11347_),
    .A2(_11351_),
    .ZN(_11352_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17470 (.I(_01791_),
    .Z(net17470));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17457 (.I(_02427_),
    .Z(net17457));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20275_ (.A1(_11320_),
    .A2(_11336_),
    .A3(net20048),
    .ZN(_11355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20276_ (.A1(net19386),
    .A2(net19837),
    .ZN(_11356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20277_ (.A1(_11356_),
    .A2(net19374),
    .ZN(_11357_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20278_ (.I(_11357_),
    .ZN(_11358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20279_ (.A1(net18918),
    .A2(net19835),
    .ZN(_11359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20280_ (.A1(_11358_),
    .A2(net18338),
    .ZN(_11360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20281_ (.A1(net18922),
    .A2(net19835),
    .ZN(_11361_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17460 (.I(_01963_),
    .Z(net17460));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20283_ (.A1(_11237_),
    .A2(net19837),
    .ZN(_11363_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20284_ (.A1(_11361_),
    .A2(net19367),
    .A3(net18911),
    .ZN(_11364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20285_ (.A1(_11360_),
    .A2(_11364_),
    .A3(net19350),
    .ZN(_11365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20286_ (.A1(net18921),
    .A2(net19838),
    .A3(net19395),
    .ZN(_11366_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20287_ (.A1(net17587),
    .A2(net19374),
    .Z(_11367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20288_ (.A1(net18332),
    .A2(_11367_),
    .ZN(_11368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20289_ (.A1(net19393),
    .A2(net17945),
    .ZN(_11369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20290_ (.A1(net19386),
    .A2(_11244_),
    .ZN(_11370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20291_ (.A1(net17583),
    .A2(_11370_),
    .ZN(_11371_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17467 (.I(_01838_),
    .Z(net17467));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20293_ (.A1(_11371_),
    .A2(net19372),
    .ZN(_11373_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17459 (.I(_01974_),
    .Z(net17459));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20295_ (.A1(_11368_),
    .A2(_11373_),
    .A3(net19352),
    .ZN(_11375_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _20296_ (.I(_11352_),
    .ZN(_11376_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17518 (.I(_15210_),
    .Z(net17518));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20298_ (.A1(_11365_),
    .A2(_11375_),
    .A3(net19827),
    .ZN(_11378_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20299_ (.A1(\sa11_sr[5] ),
    .A2(\sa01_sr[5] ),
    .ZN(_11379_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20300_ (.A1(\sa21_sr[6] ),
    .A2(\sa30_sub[6] ),
    .Z(_11380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20301_ (.A1(\sa21_sr[6] ),
    .A2(\sa30_sub[6] ),
    .ZN(_11381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20302_ (.A1(_11380_),
    .A2(_11381_),
    .ZN(_11382_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20303_ (.A1(net21404),
    .A2(net20948),
    .Z(_11383_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20304_ (.A1(_11379_),
    .A2(_11383_),
    .Z(_11384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18536 (.I(net18532),
    .Z(net18536));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20306_ (.A1(net21505),
    .A2(\text_in_r[94] ),
    .Z(_11386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20307_ (.A1(_11384_),
    .A2(net21069),
    .B(_11386_),
    .ZN(_11387_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20308_ (.A1(_07729_),
    .A2(_11387_),
    .Z(_11388_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _20309_ (.I(net20444),
    .ZN(_11389_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17453 (.I(_02586_),
    .Z(net17453));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20311_ (.A1(_11355_),
    .A2(_11378_),
    .A3(_11389_),
    .ZN(_11391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20312_ (.A1(_11237_),
    .A2(net19835),
    .ZN(_11392_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20313_ (.I(_11392_),
    .ZN(_11393_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20314_ (.I(_15721_[0]),
    .ZN(_11394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20315_ (.A1(net19387),
    .A2(_11394_),
    .ZN(_11395_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20316_ (.I(_11395_),
    .ZN(_11396_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17451 (.I(_02608_),
    .Z(net17451));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20318_ (.A1(net18331),
    .A2(_11396_),
    .A3(net19385),
    .Z(_11398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20319_ (.A1(_11393_),
    .A2(net18921),
    .ZN(_11399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20320_ (.A1(net18918),
    .A2(net19386),
    .ZN(_11400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20321_ (.A1(net17943),
    .A2(net19385),
    .A3(net18329),
    .ZN(_11401_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20322_ (.A1(_11398_),
    .A2(_11401_),
    .A3(net19347),
    .ZN(_11402_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20323_ (.A1(net20051),
    .A2(net19836),
    .A3(net18000),
    .ZN(_11403_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17445 (.I(_02756_),
    .Z(net17445));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20325_ (.A1(net19363),
    .A2(_11403_),
    .ZN(_11405_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20326_ (.I(_11405_),
    .ZN(_11406_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20327_ (.A1(_11406_),
    .A2(_11323_),
    .Z(_11407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20328_ (.A1(net19363),
    .A2(net19390),
    .ZN(_11408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20329_ (.A1(net19363),
    .A2(net19838),
    .ZN(_11409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20330_ (.A1(_11408_),
    .A2(_11409_),
    .ZN(_11410_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20331_ (.I(_11356_),
    .ZN(_11411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20332_ (.A1(_11411_),
    .A2(net18921),
    .ZN(_11412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20333_ (.A1(_11410_),
    .A2(_11412_),
    .ZN(_11413_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20334_ (.A1(_11407_),
    .A2(_11413_),
    .A3(net19356),
    .ZN(_11414_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20335_ (.A1(_11402_),
    .A2(net20048),
    .A3(_11414_),
    .ZN(_11415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20336_ (.A1(_11392_),
    .A2(net19374),
    .ZN(_11416_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18278 (.I(_13181_),
    .Z(net18278));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20338_ (.A1(_11416_),
    .A2(net19359),
    .Z(_11418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20339_ (.A1(net20050),
    .A2(net19833),
    .B(net17998),
    .ZN(_11419_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _20340_ (.A1(_11419_),
    .A2(net19374),
    .ZN(_11420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20341_ (.A1(_11399_),
    .A2(_11420_),
    .ZN(_11421_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18252 (.I(_13916_),
    .Z(net18252));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20343_ (.A1(_11418_),
    .A2(_11421_),
    .B(net20047),
    .ZN(_11423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20344_ (.A1(net19392),
    .A2(net18003),
    .ZN(_11424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20345_ (.A1(net19397),
    .A2(net17994),
    .ZN(_11425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20346_ (.A1(_11424_),
    .A2(_11425_),
    .ZN(_11426_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18388 (.I(net18387),
    .Z(net18388));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20348_ (.A1(_11426_),
    .A2(net19372),
    .B(net19352),
    .ZN(_11428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20349_ (.A1(net19386),
    .A2(net19835),
    .ZN(_11429_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20350_ (.A1(net18905),
    .A2(net19374),
    .Z(_11430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20351_ (.A1(_11430_),
    .A2(_11361_),
    .ZN(_11431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20352_ (.A1(_11428_),
    .A2(_11431_),
    .ZN(_11432_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18378 (.I(_16055_[0]),
    .Z(net18378));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20354_ (.A1(_11423_),
    .A2(_11432_),
    .B(_11389_),
    .ZN(_11434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20355_ (.A1(_11415_),
    .A2(_11434_),
    .ZN(_11435_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18729 (.I(_15150_),
    .Z(net18729));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20357_ (.A1(\sa11_sr[6] ),
    .A2(\sa01_sr[6] ),
    .Z(_11437_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20358_ (.A1(net21403),
    .A2(_11437_),
    .Z(_11438_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _20359_ (.A1(net689),
    .A2(net21285),
    .A3(_11438_),
    .Z(_11439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20360_ (.I0(_11439_),
    .I1(\text_in_r[95] ),
    .S(net21505),
    .Z(_11440_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20361_ (.A1(_07936_),
    .A2(_11440_),
    .Z(_11441_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17449 (.I(_02695_),
    .Z(net17449));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20363_ (.A1(_11391_),
    .A2(_11435_),
    .A3(net20641),
    .ZN(_11443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20364_ (.A1(net18002),
    .A2(net19833),
    .A3(net20050),
    .ZN(_11444_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20365_ (.A1(net19363),
    .A2(net17941),
    .B(net19341),
    .ZN(_11445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20366_ (.A1(net19363),
    .A2(_15728_[0]),
    .Z(_11446_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20367_ (.A1(_11445_),
    .A2(_11446_),
    .Z(_11447_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20368_ (.A1(_11447_),
    .A2(net20047),
    .Z(_11448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20369_ (.A1(_11363_),
    .A2(net17589),
    .ZN(_11449_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18633 (.I(net18623),
    .Z(net18633));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17443 (.I(_02771_),
    .Z(net17443));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20372_ (.A1(_11449_),
    .A2(net19367),
    .B(net19341),
    .ZN(_11452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20373_ (.A1(net18919),
    .A2(net19386),
    .ZN(_11453_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20374_ (.I(_15712_[0]),
    .ZN(_11454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20375_ (.A1(net19395),
    .A2(net17939),
    .ZN(_11455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20376_ (.A1(net18324),
    .A2(net19380),
    .A3(_11455_),
    .ZN(_11456_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20377_ (.I(_15709_[0]),
    .ZN(_11457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20378_ (.A1(net19395),
    .A2(_11457_),
    .ZN(_11458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20379_ (.A1(net18325),
    .A2(net17578),
    .ZN(_11459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20380_ (.A1(_11452_),
    .A2(net17353),
    .A3(_11459_),
    .ZN(_11460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20381_ (.A1(_11448_),
    .A2(_11460_),
    .ZN(_11461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20382_ (.I(_11403_),
    .ZN(_11462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20383_ (.A1(_11462_),
    .A2(net19371),
    .ZN(_11463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20384_ (.A1(_11463_),
    .A2(net19351),
    .Z(_11464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20385_ (.I(_11429_),
    .ZN(_11465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20386_ (.A1(_11465_),
    .A2(net18921),
    .ZN(_11466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20387_ (.A1(net19395),
    .A2(net17996),
    .ZN(_11467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20388_ (.A1(_11467_),
    .A2(net19374),
    .ZN(_11468_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20389_ (.I(_11468_),
    .ZN(_11469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20390_ (.A1(_11466_),
    .A2(net17352),
    .ZN(_11470_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20391_ (.A1(_11464_),
    .A2(_11470_),
    .B(net20049),
    .ZN(_11471_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20392_ (.I(_15717_[0]),
    .ZN(_11472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20393_ (.A1(_11237_),
    .A2(_11472_),
    .ZN(_11473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20394_ (.A1(_11473_),
    .A2(net19363),
    .ZN(_11474_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20395_ (.I(_11474_),
    .ZN(_11475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20396_ (.A1(_11466_),
    .A2(_11475_),
    .ZN(_11476_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20397_ (.A1(_11476_),
    .A2(net19356),
    .A3(net17354),
    .ZN(_11477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20398_ (.A1(_11471_),
    .A2(_11477_),
    .ZN(_11478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20399_ (.A1(_11461_),
    .A2(_11478_),
    .A3(_11389_),
    .ZN(_11479_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20400_ (.A1(_11453_),
    .A2(net19374),
    .Z(_11480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20401_ (.A1(_11480_),
    .A2(net17940),
    .ZN(_11481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20402_ (.A1(net17938),
    .A2(net19363),
    .Z(_11482_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20403_ (.A1(_11482_),
    .A2(net18906),
    .ZN(_11483_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20404_ (.A1(net17574),
    .A2(net19352),
    .A3(_11483_),
    .ZN(_11484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20405_ (.I(_11369_),
    .ZN(_11485_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20406_ (.A1(_11485_),
    .A2(_11462_),
    .B(net19375),
    .ZN(_11486_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20407_ (.A1(net17580),
    .A2(net19356),
    .ZN(_11487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20408_ (.A1(_11486_),
    .A2(_11487_),
    .B(net20047),
    .ZN(_11488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20409_ (.A1(_11484_),
    .A2(_11488_),
    .B(_11389_),
    .ZN(_11489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20410_ (.A1(net19394),
    .A2(net17997),
    .ZN(_11490_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20411_ (.A1(_11490_),
    .A2(net19363),
    .Z(_11491_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20412_ (.A1(_11491_),
    .A2(net19341),
    .Z(_11492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20413_ (.A1(net19391),
    .A2(net17995),
    .ZN(_11493_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20414_ (.A1(_11493_),
    .A2(net19363),
    .ZN(_11494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20415_ (.I(_11494_),
    .ZN(_11495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20416_ (.A1(_11492_),
    .A2(net17357),
    .A3(_11495_),
    .ZN(_11496_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20417_ (.A1(_11413_),
    .A2(net17573),
    .A3(net19356),
    .ZN(_11497_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20418_ (.A1(_11496_),
    .A2(net20047),
    .A3(_11497_),
    .ZN(_11498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20419_ (.A1(_11489_),
    .A2(_11498_),
    .ZN(_11499_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _20420_ (.I(_11441_),
    .ZN(_11500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20421_ (.A1(_11479_),
    .A2(_11499_),
    .A3(_11500_),
    .ZN(_11501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20422_ (.A1(_11443_),
    .A2(_11501_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20423_ (.A1(net20050),
    .A2(net19833),
    .A3(_11394_),
    .ZN(_11502_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20424_ (.A1(_11502_),
    .A2(net19363),
    .Z(_11503_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20425_ (.A1(_11503_),
    .A2(_11400_),
    .B(net19352),
    .ZN(_11504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20426_ (.A1(_11400_),
    .A2(net18905),
    .ZN(_11505_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18615 (.I(net449),
    .Z(net18615));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20428_ (.A1(_11505_),
    .A2(net19385),
    .ZN(_11507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20429_ (.A1(_11504_),
    .A2(_11507_),
    .ZN(_11508_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20430_ (.A1(_11366_),
    .A2(net19373),
    .A3(_11424_),
    .ZN(_11509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20431_ (.A1(net19389),
    .A2(net17997),
    .Z(_11510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20432_ (.A1(_11510_),
    .A2(net19379),
    .B(net19341),
    .ZN(_11511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20433_ (.A1(_11509_),
    .A2(_11511_),
    .ZN(_11512_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20434_ (.A1(_11508_),
    .A2(_11512_),
    .ZN(_11513_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17456 (.I(_02442_),
    .Z(net17456));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20436_ (.A1(_11513_),
    .A2(net19828),
    .ZN(_11515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20437_ (.A1(_11444_),
    .A2(net19374),
    .ZN(_11516_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20438_ (.A1(_11516_),
    .A2(_11465_),
    .B(net19352),
    .ZN(_11517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20439_ (.A1(net18921),
    .A2(net19838),
    .ZN(_11518_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20440_ (.A1(_11518_),
    .A2(net18905),
    .B(net19382),
    .ZN(_11519_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20441_ (.A1(_11517_),
    .A2(_11519_),
    .ZN(_11520_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20442_ (.A1(net18909),
    .A2(net17589),
    .A3(net19382),
    .ZN(_11521_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20443_ (.A1(net17936),
    .A2(net17586),
    .A3(net19369),
    .ZN(_11522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20444_ (.A1(_11521_),
    .A2(_11522_),
    .B(net19352),
    .ZN(_11523_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17450 (.I(_02641_),
    .Z(net17450));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20446_ (.A1(_11520_),
    .A2(_11523_),
    .B(net20047),
    .ZN(_11525_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17441 (.I(_02886_),
    .Z(net17441));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20448_ (.A1(_11515_),
    .A2(_11525_),
    .A3(net20444),
    .ZN(_11527_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20449_ (.A1(net19363),
    .A2(net19396),
    .Z(_11528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20450_ (.A1(_11528_),
    .A2(_11361_),
    .B(net19341),
    .ZN(_11529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20451_ (.A1(net18324),
    .A2(_11359_),
    .A3(net19380),
    .ZN(_11530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20452_ (.A1(_11529_),
    .A2(_11530_),
    .ZN(_11531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20453_ (.A1(net19388),
    .A2(_11454_),
    .ZN(_11532_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20454_ (.A1(net18909),
    .A2(net17569),
    .A3(net19381),
    .ZN(_11533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20455_ (.A1(net18908),
    .A2(net17586),
    .A3(net19369),
    .ZN(_11534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20456_ (.A1(_11533_),
    .A2(_11534_),
    .A3(net19341),
    .ZN(_11535_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20457_ (.A1(_11531_),
    .A2(_11535_),
    .A3(_11376_),
    .ZN(_11536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20458_ (.A1(net18921),
    .A2(net19395),
    .ZN(_11537_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20459_ (.A1(_11537_),
    .A2(net19363),
    .B(net19352),
    .ZN(_11538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20460_ (.A1(_11538_),
    .A2(_11456_),
    .B(_11376_),
    .ZN(_11539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20461_ (.A1(net18913),
    .A2(_11490_),
    .ZN(_11540_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20462_ (.I(_11400_),
    .ZN(_11541_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20463_ (.A1(_11540_),
    .A2(_11541_),
    .B(net19376),
    .ZN(_11542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20464_ (.A1(net19388),
    .A2(net17994),
    .ZN(_11543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20465_ (.A1(_11444_),
    .A2(_11543_),
    .ZN(_11544_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20466_ (.A1(_11544_),
    .A2(net19372),
    .B(net19341),
    .ZN(_11545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20467_ (.A1(_11542_),
    .A2(_11545_),
    .ZN(_11546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20468_ (.A1(_11539_),
    .A2(_11546_),
    .ZN(_11547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20469_ (.A1(_11536_),
    .A2(_11547_),
    .ZN(_11548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20470_ (.A1(_11548_),
    .A2(_11389_),
    .ZN(_11549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20471_ (.A1(_11527_),
    .A2(_11549_),
    .ZN(_11550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20472_ (.A1(_11550_),
    .A2(_11500_),
    .ZN(_11551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20473_ (.I(_11363_),
    .ZN(_11552_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20474_ (.A1(_11552_),
    .A2(net19383),
    .B(net19352),
    .ZN(_11553_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20475_ (.A1(_11247_),
    .A2(net19374),
    .ZN(_11554_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20476_ (.A1(_11405_),
    .A2(_11554_),
    .ZN(_11555_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20477_ (.I(_11444_),
    .ZN(_11556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20478_ (.A1(_11556_),
    .A2(net19370),
    .ZN(_11557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20479_ (.A1(_11553_),
    .A2(_11555_),
    .A3(_11557_),
    .ZN(_11558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20480_ (.A1(net18917),
    .A2(net19394),
    .ZN(_11559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20481_ (.A1(_11420_),
    .A2(net18322),
    .ZN(_11560_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20482_ (.A1(net18912),
    .A2(_11299_),
    .A3(net19376),
    .ZN(_11561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20483_ (.A1(_11560_),
    .A2(net19357),
    .A3(_11561_),
    .ZN(_11562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20484_ (.A1(_11558_),
    .A2(_11562_),
    .A3(_11376_),
    .ZN(_11563_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20485_ (.I(_11416_),
    .ZN(_11564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20486_ (.A1(_11564_),
    .A2(_11412_),
    .ZN(_11565_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20487_ (.A1(_11297_),
    .A2(net19352),
    .Z(_11566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20488_ (.A1(_11565_),
    .A2(_11566_),
    .B(_11376_),
    .ZN(_11567_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20489_ (.A1(_11395_),
    .A2(net19383),
    .Z(_11568_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20490_ (.A1(_11568_),
    .A2(net17578),
    .B(net19361),
    .ZN(_11569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20491_ (.A1(_11569_),
    .A2(_11509_),
    .ZN(_11570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20492_ (.A1(_11567_),
    .A2(_11570_),
    .ZN(_11571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20493_ (.A1(_11571_),
    .A2(_11563_),
    .B(_11389_),
    .ZN(_11572_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20494_ (.A1(net18905),
    .A2(net18910),
    .A3(net18921),
    .ZN(_11573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20495_ (.A1(_11573_),
    .A2(net19366),
    .ZN(_11574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20496_ (.A1(_11430_),
    .A2(_11299_),
    .ZN(_11575_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20497_ (.A1(_11574_),
    .A2(_11376_),
    .A3(_11575_),
    .ZN(_11576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20498_ (.A1(_11358_),
    .A2(net18323),
    .ZN(_11577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20499_ (.A1(_11577_),
    .A2(net20047),
    .A3(_11560_),
    .ZN(_11578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20500_ (.A1(_11576_),
    .A2(_11578_),
    .ZN(_11579_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20501_ (.I(_15731_[0]),
    .ZN(_11580_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20502_ (.A1(net19368),
    .A2(_11580_),
    .Z(_11581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20503_ (.A1(_11581_),
    .A2(net20045),
    .B(net19341),
    .ZN(_11582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20504_ (.A1(_11469_),
    .A2(_11412_),
    .ZN(_11583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20505_ (.A1(_11582_),
    .A2(_11583_),
    .ZN(_11584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20506_ (.A1(_11584_),
    .A2(_11389_),
    .ZN(_11585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20507_ (.A1(_11579_),
    .A2(net19345),
    .B(_11585_),
    .ZN(_11586_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20508_ (.A1(_11572_),
    .A2(_11586_),
    .B(net20641),
    .ZN(_11587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20509_ (.A1(_11551_),
    .A2(_11587_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20510_ (.A1(_11559_),
    .A2(net19363),
    .Z(_11588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20511_ (.A1(_11588_),
    .A2(net18906),
    .ZN(_11589_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20512_ (.A1(net17574),
    .A2(_11589_),
    .B(net20047),
    .ZN(_11590_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20513_ (.A1(net17940),
    .A2(net19363),
    .Z(_11591_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20514_ (.A1(_11591_),
    .A2(net17582),
    .B(_11376_),
    .ZN(_11592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20515_ (.A1(net17937),
    .A2(net17583),
    .ZN(_11593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20516_ (.A1(_11592_),
    .A2(_11593_),
    .Z(_11594_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20517_ (.A1(_11590_),
    .A2(_11594_),
    .B(net19341),
    .ZN(_11595_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20518_ (.I(_11329_),
    .ZN(_11596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20519_ (.A1(_11466_),
    .A2(_11596_),
    .ZN(_11597_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17446 (.I(_02756_),
    .Z(net17446));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20521_ (.A1(net17993),
    .A2(net19378),
    .B(net20045),
    .ZN(_11599_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18614 (.I(net18605),
    .Z(net18614));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20523_ (.A1(_11597_),
    .A2(_11599_),
    .B(net19346),
    .ZN(_11601_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20524_ (.A1(net18324),
    .A2(net18337),
    .A3(net19367),
    .ZN(_11602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20525_ (.A1(net19377),
    .A2(net17931),
    .ZN(_11603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20526_ (.A1(_11602_),
    .A2(net20045),
    .A3(_11603_),
    .ZN(_11604_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20527_ (.A1(_11601_),
    .A2(_11604_),
    .B(_11389_),
    .ZN(_11605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20528_ (.A1(_11595_),
    .A2(_11605_),
    .ZN(_11606_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20529_ (.A1(_11457_),
    .A2(_11454_),
    .Z(_11607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20530_ (.I(_11607_),
    .ZN(_11608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20531_ (.A1(net19390),
    .A2(_11608_),
    .ZN(_11609_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20532_ (.A1(net18322),
    .A2(net18908),
    .A3(_11609_),
    .ZN(_11610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20533_ (.A1(_11610_),
    .A2(net19364),
    .ZN(_11611_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20534_ (.A1(_11611_),
    .A2(net19343),
    .A3(_11583_),
    .ZN(_11612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20535_ (.A1(_11248_),
    .A2(net19380),
    .ZN(_11613_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20536_ (.A1(_11613_),
    .A2(net19355),
    .Z(_11614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20537_ (.A1(_11298_),
    .A2(net17579),
    .ZN(_11615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20538_ (.A1(_11614_),
    .A2(_11615_),
    .B(net20046),
    .ZN(_11616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20539_ (.A1(_11616_),
    .A2(_11612_),
    .ZN(_11617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20540_ (.A1(net18324),
    .A2(_11361_),
    .A3(net19368),
    .ZN(_11618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20541_ (.A1(_15735_[0]),
    .A2(net19377),
    .B(net19353),
    .ZN(_11619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20542_ (.A1(_11618_),
    .A2(_11619_),
    .B(net19832),
    .ZN(_11620_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20543_ (.A1(net19374),
    .A2(_15726_[0]),
    .Z(_11621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20544_ (.A1(net18918),
    .A2(net19374),
    .ZN(_11622_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20545_ (.A1(net18326),
    .A2(_11621_),
    .A3(_11622_),
    .ZN(_11623_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20546_ (.A1(_11623_),
    .A2(net19341),
    .Z(_11624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20547_ (.A1(_11620_),
    .A2(_11624_),
    .ZN(_11625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20548_ (.A1(_11617_),
    .A2(_11625_),
    .A3(_11389_),
    .ZN(_11626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20549_ (.A1(_11626_),
    .A2(_11606_),
    .A3(_11500_),
    .ZN(_11627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20550_ (.A1(_11366_),
    .A2(net19372),
    .ZN(_11628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20551_ (.A1(net17943),
    .A2(net19385),
    .ZN(_11629_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20552_ (.A1(net17355),
    .A2(_11628_),
    .B(_11629_),
    .C(net19356),
    .ZN(_11630_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20553_ (.A1(_11424_),
    .A2(net19374),
    .Z(_11631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20554_ (.A1(_11631_),
    .A2(net18322),
    .ZN(_11632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20555_ (.A1(net19394),
    .A2(net18001),
    .ZN(_11633_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20556_ (.A1(net18912),
    .A2(net17928),
    .A3(net19372),
    .ZN(_11634_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20557_ (.A1(_11632_),
    .A2(_11634_),
    .ZN(_11635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20558_ (.A1(_11635_),
    .A2(net19347),
    .B(net20048),
    .ZN(_11636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20559_ (.A1(_11630_),
    .A2(_11636_),
    .B(net20444),
    .ZN(_11637_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20560_ (.A1(net18914),
    .A2(_11490_),
    .A3(net19363),
    .ZN(_11638_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20561_ (.A1(_11638_),
    .A2(_11541_),
    .B(net19352),
    .ZN(_11639_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20562_ (.I(_11481_),
    .ZN(_11640_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20563_ (.A1(_11639_),
    .A2(_11640_),
    .Z(_11641_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20564_ (.I(_11618_),
    .ZN(_11642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20565_ (.A1(_11532_),
    .A2(net19374),
    .ZN(_11643_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20566_ (.I(_11502_),
    .ZN(_11644_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20567_ (.A1(_11643_),
    .A2(_11644_),
    .ZN(_11645_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17448 (.I(_02700_),
    .Z(net17448));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20569_ (.A1(_11642_),
    .A2(_11645_),
    .B(net19341),
    .ZN(_11647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20570_ (.A1(_11641_),
    .A2(_11647_),
    .ZN(_11648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20571_ (.A1(_11648_),
    .A2(net20047),
    .ZN(_11649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20572_ (.A1(_11637_),
    .A2(_11649_),
    .ZN(_11650_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20573_ (.A1(_11473_),
    .A2(net19374),
    .Z(_11651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20574_ (.A1(_11651_),
    .A2(net18906),
    .ZN(_11652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20575_ (.A1(_11591_),
    .A2(net17585),
    .ZN(_11653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20576_ (.A1(_11652_),
    .A2(_11653_),
    .B(net19341),
    .ZN(_11654_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20577_ (.I(_11425_),
    .ZN(_11655_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20578_ (.A1(net18339),
    .A2(_11655_),
    .B(net19341),
    .ZN(_11656_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20579_ (.A1(net18322),
    .A2(net19363),
    .A3(net17934),
    .Z(_11657_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20580_ (.A1(_11656_),
    .A2(_11657_),
    .ZN(_11658_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20581_ (.A1(_11654_),
    .A2(_11658_),
    .B(_11376_),
    .ZN(_11659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20582_ (.A1(net19352),
    .A2(net17935),
    .ZN(_11660_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20583_ (.A1(net17572),
    .A2(_11660_),
    .ZN(_11661_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20584_ (.A1(net18920),
    .A2(net19368),
    .Z(_11662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20585_ (.A1(_11662_),
    .A2(net19389),
    .ZN(_11663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20586_ (.A1(_11661_),
    .A2(_11663_),
    .B(_11376_),
    .ZN(_11664_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20587_ (.A1(_11495_),
    .A2(net19341),
    .Z(_11665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20588_ (.A1(_11425_),
    .A2(net19375),
    .ZN(_11666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20589_ (.A1(net17567),
    .A2(_11666_),
    .ZN(_11667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20590_ (.A1(_11665_),
    .A2(_11667_),
    .ZN(_11668_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20591_ (.A1(_11664_),
    .A2(_11668_),
    .B(_11389_),
    .ZN(_11669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20592_ (.A1(_11659_),
    .A2(_11669_),
    .B(_11500_),
    .ZN(_11670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20593_ (.A1(_11650_),
    .A2(_11670_),
    .ZN(_11671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20594_ (.A1(_11627_),
    .A2(_11671_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20595_ (.A1(_11363_),
    .A2(_11370_),
    .Z(_11672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20596_ (.A1(_11588_),
    .A2(_11672_),
    .ZN(_11673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20597_ (.A1(_11518_),
    .A2(net19390),
    .ZN(_11674_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20598_ (.I(_11516_),
    .ZN(_11675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20599_ (.A1(_11674_),
    .A2(_11675_),
    .ZN(_11676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20600_ (.A1(_11673_),
    .A2(_11676_),
    .A3(net19354),
    .ZN(_11677_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20601_ (.I(_11245_),
    .ZN(_11678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20602_ (.A1(_11367_),
    .A2(_11678_),
    .ZN(_11679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20603_ (.A1(_11364_),
    .A2(_11679_),
    .A3(net19341),
    .ZN(_11680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20604_ (.A1(_11677_),
    .A2(_11680_),
    .ZN(_11681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20605_ (.A1(_11681_),
    .A2(net19827),
    .ZN(_11682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20606_ (.A1(net19352),
    .A2(_11363_),
    .ZN(_11683_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20607_ (.I(_11359_),
    .ZN(_11684_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20608_ (.A1(_11683_),
    .A2(_11684_),
    .ZN(_11685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20609_ (.A1(_11685_),
    .A2(net18907),
    .B(_11376_),
    .ZN(_11686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20610_ (.A1(_11651_),
    .A2(net17942),
    .ZN(_11687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20611_ (.A1(_11504_),
    .A2(_11687_),
    .ZN(_11688_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20612_ (.A1(_11686_),
    .A2(_11688_),
    .B(_11389_),
    .ZN(_11689_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20613_ (.A1(_11682_),
    .A2(_11689_),
    .B(net20641),
    .ZN(_11690_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20614_ (.A1(_11672_),
    .A2(net19369),
    .ZN(_11691_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20615_ (.A1(net17584),
    .A2(net17589),
    .B(net19382),
    .ZN(_11692_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _20616_ (.A1(_11691_),
    .A2(net19354),
    .A3(_11692_),
    .Z(_11693_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18613 (.I(net18612),
    .Z(net18613));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20618_ (.A1(net17579),
    .A2(net17581),
    .A3(net19373),
    .ZN(_11695_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20619_ (.A1(_11632_),
    .A2(net19362),
    .A3(_11695_),
    .ZN(_11696_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20620_ (.A1(_11693_),
    .A2(net19828),
    .A3(_11696_),
    .ZN(_11697_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20621_ (.A1(_11358_),
    .A2(_11537_),
    .Z(_11698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20622_ (.I(_11327_),
    .ZN(_11699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20623_ (.A1(_11699_),
    .A2(net19370),
    .Z(_11700_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20624_ (.A1(_11698_),
    .A2(_11700_),
    .B(net19347),
    .ZN(_11701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20625_ (.A1(_11358_),
    .A2(net18334),
    .ZN(_11702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20626_ (.A1(_11298_),
    .A2(net18322),
    .ZN(_11703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20627_ (.A1(_11702_),
    .A2(_11703_),
    .A3(net19362),
    .ZN(_11704_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20628_ (.A1(_11701_),
    .A2(_11704_),
    .A3(net20048),
    .ZN(_11705_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20629_ (.A1(_11697_),
    .A2(_11705_),
    .A3(_11389_),
    .ZN(_11706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20630_ (.A1(_11690_),
    .A2(_11706_),
    .ZN(_11707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20631_ (.I(_11493_),
    .ZN(_11708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20632_ (.A1(net17566),
    .A2(net19371),
    .B(net20049),
    .ZN(_11709_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20633_ (.A1(_11652_),
    .A2(_11709_),
    .B(net19351),
    .ZN(_11710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20634_ (.A1(net19390),
    .A2(_11607_),
    .ZN(_11711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20635_ (.A1(_11711_),
    .A2(net19364),
    .ZN(_11712_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20636_ (.A1(_11712_),
    .A2(_11644_),
    .Z(_11713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20637_ (.A1(_11564_),
    .A2(net17586),
    .ZN(_11714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20638_ (.A1(_11713_),
    .A2(_11714_),
    .A3(net20047),
    .ZN(_11715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20639_ (.A1(_11710_),
    .A2(_11715_),
    .B(net20444),
    .ZN(_11716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20640_ (.I(_11326_),
    .ZN(_11717_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20641_ (.A1(_11717_),
    .A2(_11376_),
    .B1(net19371),
    .B2(net17577),
    .ZN(_11718_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20642_ (.I(net18324),
    .ZN(_11719_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20643_ (.A1(net17576),
    .A2(_11719_),
    .ZN(_11720_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20644_ (.A1(_11720_),
    .A2(_11700_),
    .B(net20048),
    .ZN(_11721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20645_ (.A1(_11718_),
    .A2(_11721_),
    .ZN(_11722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20646_ (.A1(_11722_),
    .A2(net19351),
    .ZN(_11723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20647_ (.A1(_11716_),
    .A2(_11723_),
    .B(_11500_),
    .ZN(_11724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20648_ (.A1(_11475_),
    .A2(net17344),
    .ZN(_11725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20649_ (.A1(_11583_),
    .A2(_11725_),
    .B(net19343),
    .ZN(_11726_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20650_ (.I(_11656_),
    .ZN(_11727_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20651_ (.A1(_11726_),
    .A2(_11727_),
    .B(net20047),
    .ZN(_11728_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20652_ (.A1(net18331),
    .A2(_11708_),
    .B(net19370),
    .ZN(_11729_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18728 (.I(net18727),
    .Z(net18728));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20654_ (.A1(_11426_),
    .A2(net19384),
    .ZN(_11731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20655_ (.A1(_11729_),
    .A2(net19347),
    .A3(_11731_),
    .ZN(_11732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20656_ (.A1(_11452_),
    .A2(_11530_),
    .ZN(_11733_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20657_ (.A1(_11732_),
    .A2(_11733_),
    .A3(net19827),
    .ZN(_11734_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20658_ (.A1(_11728_),
    .A2(net20444),
    .A3(_11734_),
    .ZN(_11735_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20659_ (.A1(_11724_),
    .A2(_11735_),
    .ZN(_11736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20660_ (.A1(_11707_),
    .A2(_11736_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20661_ (.I(net18322),
    .ZN(_11737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20662_ (.A1(_11466_),
    .A2(net19372),
    .ZN(_11738_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20663_ (.A1(_11645_),
    .A2(net19357),
    .ZN(_11739_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20664_ (.A1(_11737_),
    .A2(_11738_),
    .B(_11739_),
    .ZN(_11740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20665_ (.I(_11554_),
    .ZN(_11741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20666_ (.A1(_11741_),
    .A2(net19352),
    .Z(_11742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20667_ (.A1(_11662_),
    .A2(net19395),
    .ZN(_11743_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20668_ (.A1(net17348),
    .A2(_11742_),
    .A3(_11743_),
    .ZN(_11744_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20669_ (.A1(_11740_),
    .A2(_11744_),
    .A3(net20047),
    .ZN(_11745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20670_ (.A1(_11557_),
    .A2(_11493_),
    .Z(_11746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20671_ (.A1(_11492_),
    .A2(_11746_),
    .B(net20048),
    .ZN(_11747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20672_ (.A1(net17568),
    .A2(net19375),
    .ZN(_11748_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20673_ (.A1(_11476_),
    .A2(_11748_),
    .A3(net19356),
    .ZN(_11749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20674_ (.A1(_11747_),
    .A2(_11749_),
    .B(net20444),
    .ZN(_11750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20675_ (.A1(_11745_),
    .A2(_11750_),
    .ZN(_11751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20676_ (.A1(net18322),
    .A2(net18912),
    .ZN(_11752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20677_ (.A1(_11752_),
    .A2(net19366),
    .ZN(_11753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20678_ (.A1(_11753_),
    .A2(_11575_),
    .A3(net19360),
    .ZN(_11754_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20679_ (.A1(net19351),
    .A2(_11403_),
    .Z(_11755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20680_ (.A1(_11755_),
    .A2(net17351),
    .B(net20048),
    .ZN(_11756_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20681_ (.A1(_11754_),
    .A2(_11756_),
    .B(_11389_),
    .ZN(_11757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20682_ (.A1(_11602_),
    .A2(_11577_),
    .A3(net19360),
    .ZN(_11758_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20683_ (.A1(net18328),
    .A2(_11518_),
    .A3(net19380),
    .ZN(_11759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20684_ (.A1(net18328),
    .A2(net19366),
    .A3(_11299_),
    .ZN(_11760_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20685_ (.A1(_11759_),
    .A2(_11760_),
    .A3(net19350),
    .ZN(_11761_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20686_ (.A1(_11758_),
    .A2(_11761_),
    .A3(net20047),
    .ZN(_11762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20687_ (.A1(_11757_),
    .A2(_11762_),
    .ZN(_11763_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20688_ (.A1(_11751_),
    .A2(_11763_),
    .A3(_11500_),
    .ZN(_11764_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20689_ (.A1(net18333),
    .A2(net18322),
    .A3(net19385),
    .ZN(_11765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20690_ (.A1(_11475_),
    .A2(net18912),
    .ZN(_11766_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20691_ (.A1(_11765_),
    .A2(_11766_),
    .A3(net19349),
    .ZN(_11767_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20692_ (.A1(_11486_),
    .A2(_11364_),
    .A3(net19356),
    .ZN(_11768_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20693_ (.A1(_11767_),
    .A2(_11768_),
    .A3(net20048),
    .ZN(_11769_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20694_ (.A1(net19381),
    .A2(net19390),
    .Z(_11770_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20695_ (.A1(_11770_),
    .A2(_11361_),
    .B(net19358),
    .ZN(_11771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20696_ (.A1(_11475_),
    .A2(net18330),
    .ZN(_11772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20697_ (.A1(_11771_),
    .A2(_11772_),
    .ZN(_11773_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20698_ (.I(_15719_[0]),
    .ZN(_11774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20699_ (.A1(net19374),
    .A2(_11774_),
    .Z(_11775_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20700_ (.A1(_11591_),
    .A2(net19341),
    .A3(_11775_),
    .Z(_11776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20701_ (.A1(_11773_),
    .A2(_11776_),
    .A3(_11376_),
    .ZN(_11777_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20702_ (.A1(_11769_),
    .A2(_11389_),
    .A3(_11777_),
    .ZN(_11778_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20703_ (.A1(net19348),
    .A2(_11560_),
    .A3(net17232),
    .A4(net18340),
    .ZN(_11779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20704_ (.A1(_11358_),
    .A2(net17571),
    .ZN(_11780_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20705_ (.A1(net18904),
    .A2(net19349),
    .ZN(_11781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20706_ (.A1(_11780_),
    .A2(_11781_),
    .B(_11376_),
    .ZN(_11782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20707_ (.A1(_11779_),
    .A2(_11782_),
    .ZN(_11783_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20708_ (.A1(_11643_),
    .A2(_11556_),
    .Z(_11784_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20709_ (.A1(_11413_),
    .A2(_11784_),
    .A3(net19356),
    .ZN(_11785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20710_ (.A1(_11458_),
    .A2(net19383),
    .ZN(_11786_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20711_ (.A1(_11786_),
    .A2(net19341),
    .Z(_11787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20712_ (.A1(_11787_),
    .A2(_11628_),
    .B(net20048),
    .ZN(_11788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20713_ (.A1(_11785_),
    .A2(_11788_),
    .ZN(_11789_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20714_ (.A1(_11783_),
    .A2(_11789_),
    .A3(net20444),
    .ZN(_11790_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20715_ (.A1(_11778_),
    .A2(_11790_),
    .A3(net20641),
    .ZN(_11791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20716_ (.A1(_11764_),
    .A2(_11791_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20717_ (.A1(_11674_),
    .A2(net19365),
    .A3(_11678_),
    .Z(_11792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20718_ (.A1(_11564_),
    .A2(_11518_),
    .Z(_11793_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20719_ (.A1(_11792_),
    .A2(_11793_),
    .B(net19341),
    .ZN(_11794_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20720_ (.A1(_11662_),
    .A2(net19345),
    .ZN(_11795_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20721_ (.A1(_11759_),
    .A2(_11795_),
    .B(net20047),
    .ZN(_11796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20722_ (.A1(_11794_),
    .A2(_11796_),
    .ZN(_11797_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20723_ (.A1(_11786_),
    .A2(_11719_),
    .ZN(_11798_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20724_ (.I(_11557_),
    .ZN(_11799_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20725_ (.A1(_11798_),
    .A2(_11799_),
    .B(net19347),
    .ZN(_11800_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20726_ (.A1(net17357),
    .A2(net17350),
    .B(_11666_),
    .C(net19356),
    .ZN(_11801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20727_ (.A1(_11800_),
    .A2(_11801_),
    .ZN(_11802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20728_ (.A1(_11802_),
    .A2(net20048),
    .ZN(_11803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20729_ (.A1(_11797_),
    .A2(_11389_),
    .A3(_11803_),
    .ZN(_11804_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20730_ (.A1(_11367_),
    .A2(net19351),
    .ZN(_11805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20731_ (.A1(_11729_),
    .A2(_11805_),
    .B(_11376_),
    .ZN(_11806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20732_ (.A1(net18904),
    .A2(_11361_),
    .ZN(_11807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20733_ (.A1(_11807_),
    .A2(net19351),
    .A3(net17347),
    .ZN(_11808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20734_ (.A1(_11806_),
    .A2(_11808_),
    .B(_11389_),
    .ZN(_11809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20735_ (.A1(_11651_),
    .A2(_11466_),
    .ZN(_11810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20736_ (.A1(net19371),
    .A2(net17999),
    .ZN(_11811_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20737_ (.A1(_11464_),
    .A2(_11810_),
    .A3(_11811_),
    .ZN(_11812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20738_ (.A1(net17349),
    .A2(net17570),
    .ZN(_11813_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20739_ (.A1(_11407_),
    .A2(_11813_),
    .A3(net19356),
    .ZN(_11814_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20740_ (.A1(_11812_),
    .A2(_11814_),
    .A3(_11376_),
    .ZN(_11815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20741_ (.A1(_11809_),
    .A2(_11815_),
    .B(net20641),
    .ZN(_11816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20742_ (.A1(_11804_),
    .A2(_11816_),
    .ZN(_11817_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20743_ (.I(_11503_),
    .ZN(_11818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20744_ (.A1(_11492_),
    .A2(_11818_),
    .B(net20048),
    .ZN(_11819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20745_ (.A1(_11573_),
    .A2(net19380),
    .ZN(_11820_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20746_ (.A1(_11820_),
    .A2(net19352),
    .A3(net17231),
    .ZN(_11821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20747_ (.A1(_11819_),
    .A2(_11821_),
    .ZN(_11822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20748_ (.A1(_11412_),
    .A2(net19381),
    .ZN(_11823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20749_ (.A1(net17946),
    .A2(net19364),
    .B(net19341),
    .ZN(_11824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20750_ (.A1(_11823_),
    .A2(_11824_),
    .B(_11376_),
    .ZN(_11825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20751_ (.A1(_11631_),
    .A2(net17571),
    .ZN(_11826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20752_ (.A1(_11298_),
    .A2(net17938),
    .ZN(_11827_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20753_ (.A1(_11826_),
    .A2(_11827_),
    .A3(net19348),
    .ZN(_11828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20754_ (.A1(_11825_),
    .A2(_11828_),
    .ZN(_11829_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20755_ (.A1(_11822_),
    .A2(_11829_),
    .A3(_11389_),
    .ZN(_11830_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20756_ (.A1(_11409_),
    .A2(net19359),
    .Z(_11831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20757_ (.A1(_11360_),
    .A2(_11831_),
    .B(net20047),
    .ZN(_11832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20758_ (.A1(_11651_),
    .A2(net18330),
    .ZN(_11833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20759_ (.A1(_11399_),
    .A2(_11298_),
    .ZN(_11834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20760_ (.A1(_11833_),
    .A2(_11834_),
    .A3(net19348),
    .ZN(_11835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20761_ (.A1(_11832_),
    .A2(_11835_),
    .B(_11389_),
    .ZN(_11836_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20762_ (.A1(_11245_),
    .A2(net19365),
    .B(net19358),
    .ZN(_11837_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20763_ (.A1(_11823_),
    .A2(net17346),
    .B(_11837_),
    .ZN(_11838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20764_ (.A1(_11540_),
    .A2(net19376),
    .ZN(_11839_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20765_ (.A1(_11413_),
    .A2(net19357),
    .A3(_11839_),
    .ZN(_11840_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20766_ (.A1(_11838_),
    .A2(_11840_),
    .A3(net20047),
    .ZN(_11841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20767_ (.A1(_11836_),
    .A2(_11841_),
    .ZN(_11842_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20768_ (.A1(_11830_),
    .A2(_11842_),
    .A3(net20641),
    .ZN(_11843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20769_ (.A1(_11817_),
    .A2(_11843_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20770_ (.A1(_15724_[0]),
    .A2(_15733_[0]),
    .Z(_11844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20771_ (.A1(net19377),
    .A2(_11844_),
    .ZN(_11845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20772_ (.A1(_11845_),
    .A2(net19353),
    .ZN(_11846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20773_ (.A1(net17930),
    .A2(net18335),
    .B(_11846_),
    .ZN(_11847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20774_ (.A1(_11613_),
    .A2(net19346),
    .ZN(_11848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20775_ (.A1(net17929),
    .A2(net17934),
    .B(net19379),
    .ZN(_11849_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20776_ (.A1(_11848_),
    .A2(_11849_),
    .ZN(_11850_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20777_ (.A1(_11847_),
    .A2(_11850_),
    .B(net20444),
    .ZN(_11851_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20778_ (.I(_11399_),
    .ZN(_11852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20779_ (.A1(net18329),
    .A2(net19372),
    .ZN(_11853_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20780_ (.A1(_11852_),
    .A2(_11853_),
    .B(_11786_),
    .ZN(_11854_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20781_ (.I(_11424_),
    .ZN(_11855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20782_ (.A1(_11855_),
    .A2(net19385),
    .B(net19341),
    .ZN(_11856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20783_ (.A1(_11854_),
    .A2(_11856_),
    .ZN(_11857_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20784_ (.A1(_11326_),
    .A2(net19341),
    .Z(_11858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20785_ (.A1(_11623_),
    .A2(_11858_),
    .B(net20444),
    .ZN(_11859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20786_ (.A1(_11857_),
    .A2(_11859_),
    .ZN(_11860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20787_ (.A1(_11851_),
    .A2(_11860_),
    .ZN(_11861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20788_ (.A1(_11861_),
    .A2(net19830),
    .ZN(_11862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20789_ (.A1(net17575),
    .A2(_11395_),
    .A3(net19374),
    .ZN(_11863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20790_ (.A1(_11528_),
    .A2(_11518_),
    .ZN(_11864_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20791_ (.A1(_11863_),
    .A2(_11864_),
    .A3(_11463_),
    .ZN(_11865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20792_ (.A1(_11865_),
    .A2(net19352),
    .ZN(_11866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20793_ (.A1(_11411_),
    .A2(net19377),
    .Z(_11867_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20794_ (.A1(_11445_),
    .A2(_11867_),
    .ZN(_11868_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20795_ (.A1(net19363),
    .A2(net17935),
    .A3(net17929),
    .A4(net17934),
    .ZN(_11869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20796_ (.A1(_11868_),
    .A2(_11869_),
    .ZN(_11870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20797_ (.A1(_11866_),
    .A2(_11870_),
    .ZN(_11871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20798_ (.A1(_11871_),
    .A2(net20444),
    .ZN(_11872_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20799_ (.A1(net17590),
    .A2(net19377),
    .B(net19353),
    .ZN(_11873_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20800_ (.A1(net18327),
    .A2(net18918),
    .B(net19369),
    .ZN(_11874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20801_ (.A1(_11873_),
    .A2(_11874_),
    .B(net20444),
    .ZN(_11875_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20802_ (.A1(_11466_),
    .A2(net19369),
    .A3(_11363_),
    .ZN(_11876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20803_ (.A1(_11675_),
    .A2(net17345),
    .B(net19341),
    .ZN(_11877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20804_ (.A1(_11876_),
    .A2(_11877_),
    .ZN(_11878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20805_ (.A1(_11875_),
    .A2(_11878_),
    .B(net19831),
    .ZN(_11879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20806_ (.A1(_11872_),
    .A2(_11879_),
    .ZN(_11880_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20807_ (.A1(_11862_),
    .A2(_11880_),
    .A3(_11500_),
    .ZN(_11881_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20808_ (.A1(net17565),
    .A2(_11818_),
    .B(_11553_),
    .ZN(_11882_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20809_ (.I(_15725_[0]),
    .ZN(_11883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20810_ (.A1(_11883_),
    .A2(net19369),
    .B(net19341),
    .ZN(_11884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20811_ (.A1(_11833_),
    .A2(_11884_),
    .ZN(_11885_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20812_ (.A1(_11882_),
    .A2(_11376_),
    .A3(_11885_),
    .ZN(_11886_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20813_ (.A1(net17351),
    .A2(_11541_),
    .B(net17576),
    .ZN(_11887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20814_ (.A1(_11887_),
    .A2(net19341),
    .ZN(_11888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20815_ (.A1(_11888_),
    .A2(_11639_),
    .ZN(_11889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20816_ (.A1(_11889_),
    .A2(net20047),
    .ZN(_11890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20817_ (.A1(_11886_),
    .A2(_11890_),
    .A3(_11389_),
    .ZN(_11891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20818_ (.A1(net17933),
    .A2(_11431_),
    .ZN(_11892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20819_ (.A1(_11729_),
    .A2(_11856_),
    .ZN(_11893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20820_ (.A1(_11892_),
    .A2(_11893_),
    .A3(net20047),
    .ZN(_11894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20821_ (.A1(_11685_),
    .A2(net18321),
    .B(net20045),
    .ZN(_11895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20822_ (.A1(net18336),
    .A2(net19369),
    .A3(_11363_),
    .ZN(_11896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20823_ (.A1(net18908),
    .A2(net17932),
    .ZN(_11897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20824_ (.A1(_11897_),
    .A2(net19377),
    .ZN(_11898_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20825_ (.A1(_11896_),
    .A2(_11898_),
    .A3(net19344),
    .ZN(_11899_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20826_ (.A1(_11895_),
    .A2(_11899_),
    .ZN(_11900_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20827_ (.A1(_11894_),
    .A2(_11900_),
    .A3(net20444),
    .ZN(_11901_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20828_ (.A1(_11891_),
    .A2(_11901_),
    .A3(net20641),
    .ZN(_11902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20829_ (.A1(_11881_),
    .A2(_11902_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20830_ (.A1(_11589_),
    .A2(net19356),
    .A3(_11863_),
    .ZN(_11903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20831_ (.A1(net17568),
    .A2(net19372),
    .ZN(_11904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20832_ (.A1(_11714_),
    .A2(_11904_),
    .A3(net19341),
    .ZN(_11905_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20833_ (.A1(_11903_),
    .A2(net20047),
    .A3(_11905_),
    .ZN(_11906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20834_ (.A1(_11552_),
    .A2(net19380),
    .ZN(_11907_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20835_ (.A1(_11864_),
    .A2(_11907_),
    .A3(_11741_),
    .Z(_11908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20836_ (.A1(_11908_),
    .A2(_11771_),
    .ZN(_11909_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20837_ (.A1(_11568_),
    .A2(net19341),
    .ZN(_11910_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20838_ (.A1(_11910_),
    .A2(_11772_),
    .B(net20047),
    .ZN(_11911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20839_ (.A1(_11909_),
    .A2(_11911_),
    .ZN(_11912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20840_ (.A1(_11906_),
    .A2(_11912_),
    .A3(net20444),
    .ZN(_11913_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20841_ (.A1(net19361),
    .A2(_11326_),
    .Z(_11914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20842_ (.A1(_11505_),
    .A2(net19373),
    .ZN(_11915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20843_ (.A1(_11914_),
    .A2(_11915_),
    .B(_11376_),
    .ZN(_11916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20844_ (.A1(_11631_),
    .A2(_11366_),
    .ZN(_11917_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20845_ (.A1(_11917_),
    .A2(_11738_),
    .A3(net19349),
    .ZN(_11918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20846_ (.A1(_11918_),
    .A2(_11916_),
    .B(net20444),
    .ZN(_11919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20847_ (.A1(_11719_),
    .A2(net19380),
    .B(net19341),
    .ZN(_11920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20848_ (.A1(_11920_),
    .A2(_11602_),
    .A3(_11759_),
    .ZN(_11921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20849_ (.A1(net19380),
    .A2(net19838),
    .ZN(_11922_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20850_ (.A1(_11752_),
    .A2(net19380),
    .B(net19350),
    .C(_11922_),
    .ZN(_11923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20851_ (.A1(_11921_),
    .A2(_11923_),
    .A3(net19829),
    .ZN(_11924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20852_ (.A1(_11924_),
    .A2(_11919_),
    .ZN(_11925_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20853_ (.A1(_11925_),
    .A2(net20641),
    .A3(_11913_),
    .ZN(_11926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20854_ (.A1(net17927),
    .A2(net19363),
    .B(net19341),
    .ZN(_11927_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20855_ (.A1(_11633_),
    .A2(net19363),
    .Z(_11928_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20856_ (.A1(_11927_),
    .A2(_11928_),
    .B(net20047),
    .ZN(_11929_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20857_ (.I(_11867_),
    .ZN(_11930_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20858_ (.A1(_11622_),
    .A2(net19341),
    .Z(_11931_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20859_ (.A1(_11930_),
    .A2(_11560_),
    .A3(_11931_),
    .ZN(_11932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20860_ (.A1(_11929_),
    .A2(_11932_),
    .B(net20444),
    .ZN(_11933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20861_ (.A1(_11564_),
    .A2(net18328),
    .ZN(_11934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20862_ (.A1(_11596_),
    .A2(net17942),
    .ZN(_11935_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20863_ (.A1(_11934_),
    .A2(_11935_),
    .A3(net19345),
    .ZN(_11936_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20864_ (.A1(net19369),
    .A2(_15733_[0]),
    .Z(_11937_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20865_ (.A1(_11937_),
    .A2(net19342),
    .ZN(_11938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20866_ (.A1(_11699_),
    .A2(net19375),
    .ZN(_11939_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20867_ (.A1(_11938_),
    .A2(_11495_),
    .A3(_11939_),
    .ZN(_11940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20868_ (.A1(_11936_),
    .A2(_11940_),
    .A3(net20047),
    .ZN(_11941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20869_ (.A1(_11933_),
    .A2(_11941_),
    .B(net20641),
    .ZN(_11942_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20870_ (.A1(_11518_),
    .A2(net19395),
    .A3(net19376),
    .Z(_11943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20871_ (.A1(_11482_),
    .A2(net17942),
    .ZN(_11944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20872_ (.A1(_11614_),
    .A2(_11944_),
    .ZN(_11945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20873_ (.A1(net18331),
    .A2(net19374),
    .ZN(_11946_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20874_ (.A1(_11725_),
    .A2(_11931_),
    .A3(_11946_),
    .ZN(_11947_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20875_ (.A1(_11943_),
    .A2(_11945_),
    .B(_11947_),
    .C(net19832),
    .ZN(_11948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20876_ (.A1(net19352),
    .A2(net17588),
    .Z(_11949_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20877_ (.A1(_11949_),
    .A2(_11928_),
    .Z(_11950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20878_ (.A1(net18904),
    .A2(net18918),
    .ZN(_11951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20879_ (.A1(_11950_),
    .A2(_11951_),
    .B(_11376_),
    .ZN(_11952_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20880_ (.A1(_11588_),
    .A2(net18335),
    .ZN(_11953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20881_ (.A1(net19379),
    .A2(net17997),
    .ZN(_11954_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20882_ (.A1(_11953_),
    .A2(_11954_),
    .A3(net19346),
    .ZN(_11955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20883_ (.A1(_11952_),
    .A2(_11955_),
    .B(_11389_),
    .ZN(_11956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20884_ (.A1(_11948_),
    .A2(_11956_),
    .ZN(_11957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20885_ (.A1(_11942_),
    .A2(_11957_),
    .ZN(_11958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20886_ (.A1(_11926_),
    .A2(_11958_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20887_ (.I(\sa20_sub[1] ),
    .ZN(_11959_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20888_ (.I(\sa31_sub[1] ),
    .ZN(_11960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20889_ (.A1(_11959_),
    .A2(_11960_),
    .ZN(_11961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20890_ (.A1(\sa20_sub[1] ),
    .A2(\sa31_sub[1] ),
    .ZN(_11962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20891_ (.A1(_11961_),
    .A2(_11962_),
    .ZN(_11963_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20892_ (.I(_11963_),
    .ZN(_11964_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20893_ (.I(\sa02_sr[7] ),
    .ZN(_11965_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20894_ (.I(\sa02_sr[0] ),
    .ZN(_11966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20895_ (.A1(_11965_),
    .A2(_11966_),
    .ZN(_11967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20896_ (.A1(net21444),
    .A2(net21454),
    .ZN(_11968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20897_ (.A1(_11968_),
    .A2(_11967_),
    .ZN(_11969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20898_ (.A1(_11969_),
    .A2(_11964_),
    .ZN(_11970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20899_ (.A1(_11966_),
    .A2(net21444),
    .ZN(_11971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20900_ (.A1(_11965_),
    .A2(net21454),
    .ZN(_11972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20901_ (.A1(_11972_),
    .A2(_11971_),
    .ZN(_11973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20902_ (.A1(_11973_),
    .A2(net20903),
    .ZN(_11974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20903_ (.A1(_11970_),
    .A2(_11974_),
    .ZN(_11975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20904_ (.I(_11975_),
    .ZN(_11976_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20905_ (.A1(\sa12_sr[7] ),
    .A2(\sa12_sr[0] ),
    .Z(_11977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20906_ (.I(\sa12_sr[1] ),
    .ZN(_11978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20907_ (.A1(_11977_),
    .A2(net21027),
    .ZN(_11979_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20908_ (.I(\sa12_sr[7] ),
    .ZN(_11980_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20909_ (.I(\sa12_sr[0] ),
    .ZN(_11981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20910_ (.A1(_11980_),
    .A2(_11981_),
    .ZN(_11982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20911_ (.A1(net21386),
    .A2(\sa12_sr[0] ),
    .ZN(_11983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20912_ (.A1(_11982_),
    .A2(_11983_),
    .ZN(_11984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20913_ (.A1(_11984_),
    .A2(net21397),
    .ZN(_11985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20914_ (.A1(_11979_),
    .A2(_11985_),
    .ZN(_11986_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20915_ (.I(_11986_),
    .ZN(_11987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20916_ (.A1(_11976_),
    .A2(_11987_),
    .ZN(_11988_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17434 (.I(net17433),
    .Z(net17434));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20918_ (.A1(_11975_),
    .A2(_11986_),
    .ZN(_11990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20919_ (.A1(_11988_),
    .A2(_10378_),
    .A3(_11990_),
    .ZN(_11991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20920_ (.A1(net21501),
    .A2(\text_in_r[57] ),
    .ZN(_11992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20921_ (.A1(_11992_),
    .A2(_11991_),
    .ZN(_11993_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20922_ (.I(net21168),
    .ZN(_11994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20923_ (.A1(_11994_),
    .A2(net398),
    .ZN(_11995_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20924_ (.A1(net21023),
    .A2(net21168),
    .A3(net19826),
    .ZN(_11996_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20925_ (.A1(_11995_),
    .A2(_11996_),
    .ZN(_11997_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17431 (.I(_03230_),
    .Z(net17431));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20927_ (.A1(net21029),
    .A2(_11980_),
    .ZN(_11998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20928_ (.A1(net21444),
    .A2(net21384),
    .ZN(_11999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20929_ (.A1(_11998_),
    .A2(_11999_),
    .ZN(_12000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20930_ (.A1(_12000_),
    .A2(net21284),
    .ZN(_12001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20931_ (.I(\sa31_sub[0] ),
    .ZN(_12002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20932_ (.A1(_11998_),
    .A2(net21022),
    .A3(_11999_),
    .ZN(_12003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20933_ (.A1(_12001_),
    .A2(_12003_),
    .ZN(_12004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20934_ (.A1(net21024),
    .A2(net21345),
    .ZN(_12005_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20935_ (.I(\sa20_sub[0] ),
    .ZN(_12006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20936_ (.A1(net21020),
    .A2(net21398),
    .ZN(_12007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20937_ (.A1(_12005_),
    .A2(_12007_),
    .ZN(_12008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20938_ (.A1(_12004_),
    .A2(_12008_),
    .ZN(_12009_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20939_ (.I(_12008_),
    .ZN(_12010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20940_ (.A1(_12001_),
    .A2(_12003_),
    .A3(_12010_),
    .ZN(_12011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20941_ (.A1(_12009_),
    .A2(_12011_),
    .B(net21501),
    .ZN(_12012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20942_ (.I(\text_in_r[56] ),
    .ZN(_12013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20943_ (.A1(_12013_),
    .A2(net21501),
    .Z(_12014_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20944_ (.A1(net20278),
    .A2(_12014_),
    .B(net21169),
    .ZN(_12015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20945_ (.A1(_12009_),
    .A2(_12011_),
    .ZN(_12016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20946_ (.A1(_12016_),
    .A2(net21082),
    .ZN(_12017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20947_ (.I(net21169),
    .ZN(_12018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20948_ (.I(_12014_),
    .ZN(_12019_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20949_ (.A1(_12017_),
    .A2(_12018_),
    .A3(_12019_),
    .ZN(_12020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20950_ (.A1(_12020_),
    .A2(_12015_),
    .ZN(_15746_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20951_ (.I(\sa02_sr[1] ),
    .ZN(_12021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20952_ (.A1(_11978_),
    .A2(_12021_),
    .ZN(_12022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20953_ (.A1(\sa12_sr[1] ),
    .A2(\sa02_sr[1] ),
    .ZN(_12023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20954_ (.A1(_12022_),
    .A2(_12023_),
    .ZN(_12024_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20955_ (.I(\sa20_sub[2] ),
    .ZN(_12025_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20956_ (.A1(net20899),
    .A2(net21017),
    .ZN(_12026_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17430 (.I(_03233_),
    .Z(net17430));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20958_ (.A1(net20947),
    .A2(net21341),
    .A3(net21018),
    .ZN(_12028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20959_ (.A1(_12026_),
    .A2(_12028_),
    .ZN(_12029_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20960_ (.I(\sa31_sub[2] ),
    .ZN(_12030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20961_ (.A1(_12030_),
    .A2(net21395),
    .ZN(_12031_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20962_ (.I(\sa12_sr[2] ),
    .ZN(_12032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20963_ (.A1(_12032_),
    .A2(\sa31_sub[2] ),
    .ZN(_12033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20964_ (.A1(_12031_),
    .A2(_12033_),
    .ZN(_12034_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20965_ (.I(_12034_),
    .ZN(_12035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20966_ (.A1(_12029_),
    .A2(_12035_),
    .ZN(_12036_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20967_ (.A1(_12026_),
    .A2(_12028_),
    .A3(_12034_),
    .ZN(_12037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20968_ (.A1(_12036_),
    .A2(_12037_),
    .B(net21509),
    .ZN(_12038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20969_ (.I(\text_in_r[58] ),
    .ZN(_12039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20970_ (.A1(_12039_),
    .A2(net21509),
    .Z(_12040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20971_ (.I(net21167),
    .ZN(_12041_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20972_ (.A1(_12038_),
    .A2(_12040_),
    .B(_12041_),
    .ZN(_12042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20973_ (.A1(_12036_),
    .A2(_12037_),
    .ZN(_12043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20974_ (.A1(_12043_),
    .A2(net21082),
    .ZN(_12044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20975_ (.I(_12040_),
    .ZN(_12045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20976_ (.A1(_12044_),
    .A2(net21167),
    .A3(_12045_),
    .ZN(_12046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20977_ (.A1(_12042_),
    .A2(_12046_),
    .ZN(_12047_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place17428 (.I(_03239_),
    .Z(net17428));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20979_ (.A1(_12012_),
    .A2(_12014_),
    .B(_12018_),
    .ZN(_12048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20980_ (.A1(_12017_),
    .A2(net21169),
    .A3(_12019_),
    .ZN(_12049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20981_ (.A1(_12049_),
    .A2(_12048_),
    .ZN(_15737_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20982_ (.A1(_12038_),
    .A2(_12040_),
    .B(net21167),
    .ZN(_12050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20983_ (.A1(_12044_),
    .A2(_12041_),
    .A3(_12045_),
    .ZN(_12051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20984_ (.A1(_12050_),
    .A2(_12051_),
    .ZN(_12052_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18612 (.I(net18605),
    .Z(net18612));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20986_ (.A1(_12047_),
    .A2(net19333),
    .ZN(_12053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _20987_ (.I(_15753_[0]),
    .ZN(_12054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20988_ (.A1(net17564),
    .A2(net19329),
    .ZN(_12055_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20989_ (.A1(\sa20_sub[3] ),
    .A2(\sa31_sub[3] ),
    .Z(_12056_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20990_ (.I(\sa02_sr[2] ),
    .ZN(_12057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20991_ (.A1(net21030),
    .A2(_12057_),
    .ZN(_12058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20992_ (.A1(net21446),
    .A2(net21451),
    .ZN(_12059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20993_ (.A1(_12058_),
    .A2(_12059_),
    .ZN(_12060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20994_ (.A1(_12056_),
    .A2(_12060_),
    .ZN(_12061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20995_ (.A1(_12057_),
    .A2(net21446),
    .ZN(_12062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20996_ (.A1(net21030),
    .A2(net21451),
    .ZN(_12063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20997_ (.A1(_12062_),
    .A2(_12063_),
    .ZN(_12064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20998_ (.I(\sa20_sub[3] ),
    .ZN(_12065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20999_ (.I(\sa31_sub[3] ),
    .ZN(_12066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21000_ (.A1(_12065_),
    .A2(_12066_),
    .ZN(_12067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21001_ (.A1(\sa20_sub[3] ),
    .A2(\sa31_sub[3] ),
    .ZN(_12068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21002_ (.A1(_12067_),
    .A2(_12068_),
    .ZN(_12069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21003_ (.A1(_12064_),
    .A2(_12069_),
    .ZN(_12070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21004_ (.A1(_12061_),
    .A2(_12070_),
    .ZN(_12071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21005_ (.I(_12071_),
    .ZN(_12072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21006_ (.I(\sa12_sr[3] ),
    .ZN(_12073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21007_ (.A1(_12073_),
    .A2(net21385),
    .ZN(_12074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21008_ (.A1(net21025),
    .A2(\sa12_sr[3] ),
    .ZN(_12075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21009_ (.A1(_12074_),
    .A2(_12075_),
    .ZN(_12076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21010_ (.A1(_12076_),
    .A2(net21394),
    .ZN(_12077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21011_ (.A1(net21025),
    .A2(_12073_),
    .ZN(_12078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21012_ (.A1(net21385),
    .A2(net21391),
    .ZN(_12079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21013_ (.A1(_12078_),
    .A2(_12079_),
    .ZN(_12080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21014_ (.A1(_12080_),
    .A2(net21016),
    .ZN(_12081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21015_ (.A1(_12077_),
    .A2(_12081_),
    .ZN(_12082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21016_ (.A1(_12072_),
    .A2(net20639),
    .ZN(_12083_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21017_ (.I(_12082_),
    .ZN(_12084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21018_ (.A1(_12084_),
    .A2(net20640),
    .ZN(_12085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21019_ (.A1(_12083_),
    .A2(_12085_),
    .A3(net21082),
    .ZN(_12086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21020_ (.A1(net21513),
    .A2(\text_in_r[59] ),
    .ZN(_12087_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21021_ (.A1(_12086_),
    .A2(net21166),
    .A3(_12087_),
    .ZN(_12088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21022_ (.A1(_12072_),
    .A2(_12084_),
    .ZN(_12089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21023_ (.A1(_12071_),
    .A2(_12082_),
    .ZN(_12090_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21024_ (.A1(_12089_),
    .A2(_12090_),
    .A3(net21082),
    .ZN(_12091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21025_ (.I(net21166),
    .ZN(_12092_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21026_ (.A1(net21082),
    .A2(\text_in_r[59] ),
    .Z(_12093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21027_ (.A1(_12091_),
    .A2(_12092_),
    .A3(_12093_),
    .ZN(_12094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21028_ (.A1(_12088_),
    .A2(_12094_),
    .ZN(_12095_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place17436 (.I(_03156_),
    .Z(net17436));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17424 (.I(_03252_),
    .Z(net17424));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21031_ (.A1(net18902),
    .A2(_12055_),
    .A3(net19319),
    .Z(_12098_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21032_ (.A1(\sa12_sr[4] ),
    .A2(\sa31_sub[4] ),
    .Z(_12099_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21033_ (.A1(_12099_),
    .A2(_12076_),
    .Z(_12100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21034_ (.A1(_12099_),
    .A2(_12076_),
    .ZN(_12101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21035_ (.A1(_12100_),
    .A2(_12101_),
    .ZN(_12102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21036_ (.I(_12102_),
    .ZN(_12103_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21037_ (.A1(net21446),
    .A2(\sa02_sr[3] ),
    .Z(_12104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21038_ (.I(\sa20_sub[4] ),
    .ZN(_12105_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21039_ (.A1(_12104_),
    .A2(_12105_),
    .ZN(_12106_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21040_ (.I(_12106_),
    .ZN(_12107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21041_ (.A1(_12104_),
    .A2(_12105_),
    .ZN(_12108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21042_ (.A1(_12107_),
    .A2(_12108_),
    .ZN(_12109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21043_ (.A1(_12103_),
    .A2(_12109_),
    .ZN(_12110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21044_ (.I(_12108_),
    .ZN(_12111_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21045_ (.A1(_12111_),
    .A2(_12106_),
    .ZN(_12112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21046_ (.A1(_12112_),
    .A2(_12102_),
    .ZN(_12113_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21047_ (.A1(_12110_),
    .A2(_12113_),
    .A3(net21081),
    .ZN(_12114_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18611 (.I(net449),
    .Z(net18611));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21049_ (.A1(net21510),
    .A2(\text_in_r[60] ),
    .ZN(_12116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21050_ (.A1(_12116_),
    .A2(_12114_),
    .ZN(_12117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21051_ (.A1(_12117_),
    .A2(net21165),
    .ZN(_12118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21052_ (.I(net21165),
    .ZN(_12119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21053_ (.A1(_12114_),
    .A2(_12119_),
    .A3(_12116_),
    .ZN(_12120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21054_ (.A1(_12118_),
    .A2(_12120_),
    .ZN(_12121_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18588 (.I(net18587),
    .Z(net18588));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21056_ (.A1(_12098_),
    .A2(net18894),
    .ZN(_12123_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21057_ (.I(_12053_),
    .ZN(_12124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21058_ (.A1(_12124_),
    .A2(net18319),
    .ZN(_12125_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21059_ (.A1(_12086_),
    .A2(_12092_),
    .A3(_12087_),
    .ZN(_12126_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21060_ (.A1(_12091_),
    .A2(net21166),
    .A3(_12093_),
    .ZN(_12127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21061_ (.A1(_12127_),
    .A2(_12126_),
    .ZN(_12128_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17417 (.I(_03291_),
    .Z(net17417));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17415 (.I(_03366_),
    .Z(net17415));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21064_ (.A1(_11993_),
    .A2(net21168),
    .ZN(_12131_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21065_ (.A1(_11994_),
    .A2(_11991_),
    .A3(_11992_),
    .ZN(_12132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21066_ (.A1(_12132_),
    .A2(_12131_),
    .ZN(_15738_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21067_ (.A1(net19331),
    .A2(net18316),
    .ZN(_12133_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17418 (.I(_03288_),
    .Z(net17418));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21069_ (.A1(_12125_),
    .A2(net19308),
    .A3(net17925),
    .ZN(_12135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21070_ (.A1(_12123_),
    .A2(_12135_),
    .ZN(_12136_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21071_ (.I(_15741_[0]),
    .ZN(_12137_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _21072_ (.A1(_12047_),
    .A2(_12137_),
    .ZN(_12138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21073_ (.A1(net19303),
    .A2(_12138_),
    .ZN(_12139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21074_ (.A1(net18887),
    .A2(_12139_),
    .ZN(_12140_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18610 (.I(net449),
    .Z(net18610));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21076_ (.A1(net18316),
    .A2(net19303),
    .A3(net19338),
    .ZN(_12142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21077_ (.I(_12142_),
    .ZN(_12143_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21078_ (.A1(net681),
    .A2(_12143_),
    .ZN(_12144_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21079_ (.A1(net641),
    .A2(net19340),
    .A3(net19330),
    .ZN(_12145_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21080_ (.A1(_12145_),
    .A2(net19322),
    .A3(net18900),
    .ZN(_12146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21081_ (.A1(_12144_),
    .A2(_12146_),
    .ZN(_12147_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21082_ (.A1(\sa12_sr[4] ),
    .A2(\sa02_sr[4] ),
    .Z(_12148_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21083_ (.A1(\sa20_sub[5] ),
    .A2(\sa31_sub[5] ),
    .Z(_12149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21084_ (.A1(\sa20_sub[5] ),
    .A2(\sa31_sub[5] ),
    .ZN(_12150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21085_ (.A1(_12149_),
    .A2(_12150_),
    .ZN(_12151_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21086_ (.A1(\sa12_sr[5] ),
    .A2(net20946),
    .Z(_12152_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21087_ (.A1(net21013),
    .A2(_12152_),
    .Z(_12153_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21088_ (.I(net21164),
    .ZN(_12154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21089_ (.A1(net21510),
    .A2(\text_in_r[61] ),
    .ZN(_12155_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21090_ (.A1(_12153_),
    .A2(net21510),
    .B(_12154_),
    .C(_12155_),
    .ZN(_12156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21091_ (.A1(_12153_),
    .A2(net21083),
    .ZN(_12157_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21092_ (.A1(net21083),
    .A2(\text_in_r[61] ),
    .Z(_12158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21093_ (.A1(_12157_),
    .A2(net21164),
    .A3(_12158_),
    .ZN(_12159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21094_ (.A1(_12156_),
    .A2(_12159_),
    .ZN(_12160_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17413 (.I(_03416_),
    .Z(net17413));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21096_ (.A1(_12136_),
    .A2(_12147_),
    .A3(net20276),
    .ZN(_12162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21097_ (.I(_15744_[0]),
    .ZN(_12163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21098_ (.A1(_12052_),
    .A2(_12163_),
    .ZN(_12164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21099_ (.A1(_12164_),
    .A2(net19317),
    .ZN(_12165_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21100_ (.I(_12165_),
    .ZN(_12166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21101_ (.A1(_12125_),
    .A2(_12166_),
    .ZN(_12167_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17411 (.I(_03483_),
    .Z(net17411));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18695 (.I(net18694),
    .Z(net18695));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21104_ (.A1(net18901),
    .A2(net19303),
    .Z(_12170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21105_ (.I(_12170_),
    .ZN(_12171_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21106_ (.A1(_12167_),
    .A2(net18894),
    .A3(_12171_),
    .ZN(_12172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17421 (.I(_03274_),
    .Z(net17421));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21108_ (.A1(net19334),
    .A2(net19330),
    .ZN(_12174_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17416 (.I(_03366_),
    .Z(net17416));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21110_ (.A1(_12125_),
    .A2(net19316),
    .A3(net18886),
    .ZN(_12176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21111_ (.A1(net17609),
    .A2(net19331),
    .ZN(_12177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21112_ (.A1(net20043),
    .A2(net19824),
    .A3(net17606),
    .ZN(_12178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21113_ (.A1(_12177_),
    .A2(_12178_),
    .ZN(_12179_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17412 (.I(_03441_),
    .Z(net17412));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17405 (.I(_04085_),
    .Z(net17405));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21116_ (.A1(_12179_),
    .A2(net19319),
    .B(net18887),
    .ZN(_12182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21117_ (.A1(_12176_),
    .A2(_12182_),
    .ZN(_12183_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21118_ (.I(_12160_),
    .ZN(_12184_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17402 (.I(_04147_),
    .Z(net17402));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21120_ (.A1(_12172_),
    .A2(_12183_),
    .A3(net20040),
    .ZN(_12186_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21121_ (.A1(\sa12_sr[5] ),
    .A2(\sa02_sr[5] ),
    .ZN(_12187_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21122_ (.A1(\sa20_sub[6] ),
    .A2(\sa31_sub[6] ),
    .Z(_12188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21123_ (.A1(\sa20_sub[6] ),
    .A2(\sa31_sub[6] ),
    .ZN(_12189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21124_ (.A1(_12188_),
    .A2(_12189_),
    .ZN(_12190_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21125_ (.A1(net21388),
    .A2(_12190_),
    .Z(_12191_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21126_ (.A1(_12187_),
    .A2(_12191_),
    .Z(_12192_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17400 (.I(_04199_),
    .Z(net17400));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21128_ (.A1(net21507),
    .A2(\text_in_r[62] ),
    .Z(_12194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21129_ (.A1(_12192_),
    .A2(net21081),
    .B(_12194_),
    .ZN(_12195_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21130_ (.A1(net21162),
    .A2(_12195_),
    .Z(_12196_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17404 (.I(_04129_),
    .Z(net17404));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _21132_ (.I(_12196_),
    .ZN(_12198_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17454 (.I(_02586_),
    .Z(net17454));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21134_ (.A1(_12162_),
    .A2(_12186_),
    .A3(net20273),
    .ZN(_12200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21135_ (.A1(net19330),
    .A2(net19340),
    .ZN(_12201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21136_ (.A1(_12201_),
    .A2(net19303),
    .Z(_12202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21137_ (.A1(net645),
    .A2(net19334),
    .ZN(_12203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21138_ (.A1(_12202_),
    .A2(_12203_),
    .ZN(_12204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21139_ (.A1(net19334),
    .A2(net18319),
    .ZN(_12205_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17395 (.I(_04286_),
    .Z(net17395));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17406 (.I(_03972_),
    .Z(net17406));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21142_ (.A1(net19338),
    .A2(net19340),
    .ZN(_12208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21143_ (.A1(_12205_),
    .A2(net19319),
    .A3(_12208_),
    .ZN(_12209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21144_ (.A1(_12117_),
    .A2(_12119_),
    .ZN(_12210_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21145_ (.A1(net20042),
    .A2(net21165),
    .A3(_12116_),
    .ZN(_12211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21146_ (.A1(_12211_),
    .A2(_12210_),
    .ZN(_12212_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17422 (.I(_03274_),
    .Z(net17422));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17392 (.I(_04836_),
    .Z(net17392));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21149_ (.A1(_12204_),
    .A2(_12209_),
    .A3(net648),
    .ZN(_12215_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21150_ (.I(_15739_[0]),
    .ZN(_12216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21151_ (.A1(net19338),
    .A2(_12216_),
    .ZN(_12217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21152_ (.I(_15747_[0]),
    .ZN(_12218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21153_ (.A1(net19331),
    .A2(_12218_),
    .ZN(_12219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21154_ (.A1(_12217_),
    .A2(_12219_),
    .ZN(_12220_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17399 (.I(_04250_),
    .Z(net17399));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17389 (.I(_05433_),
    .Z(net17389));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21157_ (.A1(_12220_),
    .A2(net19319),
    .B(net648),
    .ZN(_12223_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21158_ (.A1(net19338),
    .A2(net19340),
    .Z(_12224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21159_ (.A1(net18319),
    .A2(_12224_),
    .ZN(_12225_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21160_ (.I(_15740_[0]),
    .ZN(_12226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21161_ (.A1(_12226_),
    .A2(net19331),
    .ZN(_12227_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21162_ (.A1(net17337),
    .A2(net647),
    .Z(_12228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21163_ (.A1(_12225_),
    .A2(_12228_),
    .ZN(_12229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21164_ (.A1(_12223_),
    .A2(_12229_),
    .ZN(_12230_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21165_ (.A1(_12215_),
    .A2(_12230_),
    .A3(net20040),
    .ZN(_12231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21166_ (.A1(net647),
    .A2(net17559),
    .A3(net19331),
    .ZN(_12232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21167_ (.A1(net654),
    .A2(net19337),
    .ZN(_12233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21168_ (.A1(net19317),
    .A2(_12233_),
    .ZN(_12234_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21169_ (.A1(net17921),
    .A2(_12232_),
    .A3(_12234_),
    .ZN(_12235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21170_ (.A1(_12235_),
    .A2(net648),
    .ZN(_12236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21171_ (.A1(net19331),
    .A2(_12216_),
    .ZN(_12237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21172_ (.A1(_12218_),
    .A2(net19338),
    .ZN(_12238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21173_ (.A1(net17334),
    .A2(_12238_),
    .ZN(_12239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21174_ (.A1(_12239_),
    .A2(net19314),
    .ZN(_12240_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21175_ (.A1(_12047_),
    .A2(net17610),
    .ZN(_12241_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17397 (.I(_04266_),
    .Z(net17397));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21177_ (.A1(net17337),
    .A2(_12241_),
    .A3(net19319),
    .ZN(_12243_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17391 (.I(_05088_),
    .Z(net17391));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21179_ (.A1(_12240_),
    .A2(_12243_),
    .A3(net18892),
    .ZN(_12245_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17386 (.I(_05505_),
    .Z(net17386));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21181_ (.A1(_12236_),
    .A2(_12245_),
    .A3(net20276),
    .ZN(_12247_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17387 (.I(_05499_),
    .Z(net17387));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21183_ (.A1(_12231_),
    .A2(_12247_),
    .A3(net20442),
    .ZN(_12249_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17382 (.I(_05726_),
    .Z(net17382));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17380 (.I(_06082_),
    .Z(net17380));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21186_ (.A1(net21387),
    .A2(net21447),
    .Z(_12252_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21187_ (.A1(net21385),
    .A2(_12252_),
    .Z(_12253_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _21188_ (.A1(net21332),
    .A2(net21274),
    .A3(_12253_),
    .Z(_12254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21189_ (.I0(_12254_),
    .I1(\text_in_r[63] ),
    .S(net21507),
    .Z(_12255_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21190_ (.A1(net21161),
    .A2(_12255_),
    .ZN(_12256_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17379 (.I(_06172_),
    .Z(net17379));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21192_ (.A1(_12200_),
    .A2(_12249_),
    .A3(net20637),
    .ZN(_12258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21193_ (.A1(net19335),
    .A2(net17607),
    .ZN(_12259_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _21194_ (.I(_12259_),
    .ZN(_12260_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17383 (.I(_05680_),
    .Z(net17383));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21196_ (.A1(_12260_),
    .A2(net19304),
    .B(net18875),
    .ZN(_12262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21197_ (.A1(_12146_),
    .A2(_12262_),
    .ZN(_12263_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21198_ (.A1(net20044),
    .A2(net19825),
    .A3(_15749_[0]),
    .ZN(_12264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21199_ (.A1(_12259_),
    .A2(net17558),
    .B(net19325),
    .ZN(_12265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21200_ (.A1(net487),
    .A2(net19317),
    .ZN(_12266_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21201_ (.I(_12266_),
    .ZN(_12267_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21202_ (.A1(_12265_),
    .A2(net524),
    .ZN(_12268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21203_ (.A1(_12268_),
    .A2(net648),
    .ZN(_12269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21204_ (.A1(_12263_),
    .A2(_12269_),
    .A3(_12198_),
    .ZN(_12270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21205_ (.A1(_12208_),
    .A2(_12237_),
    .ZN(_12271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21206_ (.A1(_12271_),
    .A2(net19328),
    .B(net18875),
    .ZN(_12272_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21207_ (.A1(net19334),
    .A2(net435),
    .A3(net19330),
    .ZN(_12273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21208_ (.A1(net20043),
    .A2(net19824),
    .A3(_12163_),
    .ZN(_12274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21209_ (.A1(_12273_),
    .A2(net19301),
    .A3(_12274_),
    .ZN(_12275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21210_ (.A1(net19335),
    .A2(net17608),
    .Z(_12276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21211_ (.A1(net647),
    .A2(_12276_),
    .ZN(_12277_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21212_ (.A1(_12272_),
    .A2(_12275_),
    .A3(_12277_),
    .ZN(_12278_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21213_ (.A1(net20043),
    .A2(_15740_[0]),
    .A3(net19823),
    .ZN(_12279_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21214_ (.I(_12279_),
    .ZN(_12280_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17375 (.I(_06225_),
    .Z(net17375));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21216_ (.A1(net19301),
    .A2(_12280_),
    .B(net18887),
    .ZN(_12282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21217_ (.A1(net19318),
    .A2(_15760_[0]),
    .ZN(_12283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21218_ (.A1(_12282_),
    .A2(_12283_),
    .B(_12198_),
    .ZN(_12284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21219_ (.A1(_12278_),
    .A2(_12284_),
    .ZN(_12285_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21220_ (.A1(_12270_),
    .A2(_12285_),
    .A3(net20274),
    .ZN(_12286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21221_ (.A1(net17340),
    .A2(net19320),
    .ZN(_12287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21222_ (.A1(_12287_),
    .A2(net648),
    .Z(_12288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21223_ (.A1(net19336),
    .A2(_15747_[0]),
    .ZN(_12289_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21224_ (.A1(_12289_),
    .A2(net19303),
    .Z(_12290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21225_ (.A1(net17328),
    .A2(net643),
    .ZN(_12291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21226_ (.A1(_12288_),
    .A2(_12291_),
    .B(_12198_),
    .ZN(_12292_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21227_ (.I(_12140_),
    .ZN(_12293_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21228_ (.I(_15749_[0]),
    .ZN(_12294_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21229_ (.A1(_12294_),
    .A2(net19823),
    .A3(net20043),
    .ZN(_12295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21230_ (.A1(net19317),
    .A2(_12295_),
    .Z(_12296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21231_ (.A1(_12273_),
    .A2(_12296_),
    .ZN(_12297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21232_ (.A1(net682),
    .A2(_12297_),
    .ZN(_12298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21233_ (.A1(_12292_),
    .A2(_12298_),
    .B(net20274),
    .ZN(_12299_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21234_ (.A1(_12139_),
    .A2(_12165_),
    .Z(_12300_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21235_ (.I(_12217_),
    .ZN(_12301_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17396 (.I(_04275_),
    .Z(net17396));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21237_ (.A1(_12301_),
    .A2(net19305),
    .ZN(_12303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21238_ (.A1(_12300_),
    .A2(_12303_),
    .B(net18887),
    .ZN(_12304_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _21239_ (.I(_12201_),
    .ZN(_12305_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21240_ (.I(_12238_),
    .ZN(_12306_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21241_ (.A1(_12305_),
    .A2(_12306_),
    .B(net19319),
    .ZN(_12307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21242_ (.A1(net19330),
    .A2(net18319),
    .ZN(_12308_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21243_ (.A1(_12308_),
    .A2(net19316),
    .A3(net17554),
    .ZN(_12309_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17388 (.I(_05485_),
    .Z(net17388));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21245_ (.A1(_12307_),
    .A2(_12309_),
    .B(net648),
    .ZN(_12311_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21246_ (.A1(_12304_),
    .A2(_12311_),
    .B(_12198_),
    .ZN(_12312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21247_ (.A1(_12299_),
    .A2(_12312_),
    .ZN(_12313_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21248_ (.I(_12256_),
    .ZN(_12314_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21249_ (.A1(_12286_),
    .A2(_12313_),
    .A3(_12314_),
    .ZN(_12315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21250_ (.A1(_12258_),
    .A2(_12315_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21251_ (.A1(net18316),
    .A2(net19338),
    .ZN(_12316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21252_ (.A1(_12166_),
    .A2(_12316_),
    .ZN(_12317_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21253_ (.A1(net18883),
    .A2(_12241_),
    .A3(net19308),
    .ZN(_12318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21254_ (.A1(_12317_),
    .A2(net18898),
    .A3(_12318_),
    .ZN(_12319_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17370 (.I(_06338_),
    .Z(net17370));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21256_ (.A1(net17342),
    .A2(net19308),
    .B(net18894),
    .ZN(_12321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21257_ (.A1(net17333),
    .A2(net17554),
    .ZN(_12322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21258_ (.A1(_12322_),
    .A2(net19324),
    .ZN(_12323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21259_ (.A1(net18874),
    .A2(net19309),
    .ZN(_12324_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21260_ (.A1(_12321_),
    .A2(_12323_),
    .A3(_12324_),
    .ZN(_12325_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17398 (.I(_04261_),
    .Z(net17398));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21262_ (.A1(_12319_),
    .A2(_12325_),
    .A3(net20040),
    .ZN(_12327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21263_ (.A1(_12170_),
    .A2(net17920),
    .ZN(_12328_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21264_ (.A1(net18887),
    .A2(_12266_),
    .Z(_12329_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21265_ (.A1(_12328_),
    .A2(_12329_),
    .B(net20040),
    .ZN(_12330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21266_ (.A1(net19307),
    .A2(_12055_),
    .Z(_12331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21267_ (.A1(net19336),
    .A2(_12137_),
    .ZN(_12332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21268_ (.A1(_12331_),
    .A2(net17326),
    .B(net18887),
    .ZN(_12333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21269_ (.A1(_12225_),
    .A2(net19319),
    .A3(net17562),
    .ZN(_12334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21270_ (.A1(_12333_),
    .A2(_12334_),
    .ZN(_12335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21271_ (.A1(_12330_),
    .A2(_12335_),
    .ZN(_12336_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21272_ (.A1(_12336_),
    .A2(_12327_),
    .B(net20442),
    .ZN(_12337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21273_ (.A1(net18319),
    .A2(net19338),
    .ZN(_12338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21274_ (.A1(_12202_),
    .A2(_12338_),
    .ZN(_12339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21275_ (.A1(_12339_),
    .A2(_12317_),
    .ZN(_12340_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21276_ (.A1(_12340_),
    .A2(net20275),
    .B(net18896),
    .ZN(_12341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21277_ (.A1(_12305_),
    .A2(net641),
    .B(net19313),
    .ZN(_12342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21278_ (.A1(_12342_),
    .A2(_12125_),
    .ZN(_12343_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21279_ (.A1(_12174_),
    .A2(_12241_),
    .A3(net19313),
    .ZN(_12344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21280_ (.A1(_12343_),
    .A2(_12344_),
    .ZN(_12345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21281_ (.A1(_12345_),
    .A2(net20040),
    .ZN(_12346_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21282_ (.A1(net20638),
    .A2(net20443),
    .B(_15763_[0]),
    .ZN(_12347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21283_ (.A1(_12347_),
    .A2(net19321),
    .ZN(_12348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21284_ (.A1(_12290_),
    .A2(_12145_),
    .ZN(_12349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21285_ (.A1(_12348_),
    .A2(_12349_),
    .A3(net18895),
    .ZN(_12350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21286_ (.A1(_12350_),
    .A2(net20442),
    .ZN(_12351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21287_ (.A1(_12341_),
    .A2(_12346_),
    .B(_12351_),
    .ZN(_12352_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21288_ (.A1(_12352_),
    .A2(_12337_),
    .B(net20637),
    .ZN(_12353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21289_ (.A1(net19336),
    .A2(_12054_),
    .ZN(_12354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21290_ (.A1(_12354_),
    .A2(net19322),
    .ZN(_12355_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21291_ (.I(_12355_),
    .ZN(_12356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21292_ (.A1(_12356_),
    .A2(net642),
    .B(net18888),
    .ZN(_12357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21293_ (.A1(net17923),
    .A2(net18885),
    .ZN(_12358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21294_ (.A1(_12358_),
    .A2(net19302),
    .ZN(_12359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21295_ (.A1(_12357_),
    .A2(_12359_),
    .ZN(_12360_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21296_ (.A1(net19331),
    .A2(net17607),
    .Z(_12361_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21297_ (.A1(_12361_),
    .A2(net647),
    .B(net18875),
    .ZN(_12362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21298_ (.A1(_12334_),
    .A2(_12362_),
    .ZN(_12363_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21299_ (.A1(_12360_),
    .A2(_12363_),
    .A3(net20040),
    .ZN(_12364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21300_ (.A1(net19340),
    .A2(net18319),
    .ZN(_12365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21301_ (.A1(_12365_),
    .A2(net655),
    .ZN(_12366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21302_ (.A1(_12366_),
    .A2(net19328),
    .ZN(_12367_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21303_ (.A1(net17554),
    .A2(net19301),
    .Z(_12368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21304_ (.A1(_12368_),
    .A2(net18886),
    .ZN(_12369_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21305_ (.A1(_12367_),
    .A2(net18893),
    .A3(_12369_),
    .ZN(_12370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21306_ (.A1(_12259_),
    .A2(net17336),
    .ZN(_12371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21307_ (.A1(_12371_),
    .A2(net19325),
    .ZN(_12372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21308_ (.A1(_12271_),
    .A2(net19301),
    .ZN(_12373_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21309_ (.A1(_12372_),
    .A2(_12373_),
    .A3(net648),
    .ZN(_12374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21310_ (.A1(_12370_),
    .A2(_12374_),
    .A3(net20277),
    .ZN(_12375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21311_ (.A1(_12364_),
    .A2(_12375_),
    .A3(net20273),
    .ZN(_12376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21312_ (.A1(_12338_),
    .A2(net19319),
    .ZN(_12377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21313_ (.A1(_12377_),
    .A2(net642),
    .Z(_12378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21314_ (.A1(_12260_),
    .A2(net19305),
    .B(net18887),
    .ZN(_12379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21315_ (.A1(_12378_),
    .A2(_12379_),
    .B(net20040),
    .ZN(_12380_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _21316_ (.I(_12234_),
    .ZN(_12381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21317_ (.A1(net17343),
    .A2(_12381_),
    .ZN(_12382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21318_ (.A1(_12275_),
    .A2(net18887),
    .A3(_12382_),
    .ZN(_12383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21319_ (.A1(_12380_),
    .A2(_12383_),
    .ZN(_12384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21320_ (.A1(_12164_),
    .A2(net19303),
    .Z(_12385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21321_ (.A1(net17227),
    .A2(net18882),
    .ZN(_12386_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18700 (.I(net18699),
    .Z(net18700));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17378 (.I(_06201_),
    .Z(net17378));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21324_ (.A1(net18903),
    .A2(net17338),
    .A3(net19319),
    .ZN(_12389_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21325_ (.A1(_12389_),
    .A2(net648),
    .A3(_12386_),
    .ZN(_12390_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21326_ (.A1(net19317),
    .A2(net19336),
    .Z(_12391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21327_ (.A1(net18873),
    .A2(_12205_),
    .B(net18875),
    .ZN(_12392_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21328_ (.A1(_12308_),
    .A2(_12203_),
    .A3(net19309),
    .ZN(_12393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21329_ (.A1(_12392_),
    .A2(_12393_),
    .ZN(_12394_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21330_ (.A1(_12390_),
    .A2(net20040),
    .A3(_12394_),
    .ZN(_12395_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21331_ (.A1(_12384_),
    .A2(_12395_),
    .A3(net20442),
    .ZN(_12396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21332_ (.A1(_12376_),
    .A2(_12396_),
    .A3(_12314_),
    .ZN(_12397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21333_ (.A1(_12353_),
    .A2(_12397_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21334_ (.A1(net18320),
    .A2(net19335),
    .ZN(_12398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21335_ (.A1(_12274_),
    .A2(net19317),
    .ZN(_12399_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21336_ (.A1(_12398_),
    .A2(_12399_),
    .ZN(_12400_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21337_ (.A1(_12400_),
    .A2(_12265_),
    .B(net18891),
    .ZN(_12401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21338_ (.A1(net17558),
    .A2(_12178_),
    .ZN(_12402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21339_ (.A1(_12402_),
    .A2(net19301),
    .ZN(_12403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21340_ (.A1(_12174_),
    .A2(net19326),
    .A3(_12274_),
    .ZN(_12404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21341_ (.A1(_12403_),
    .A2(_12404_),
    .ZN(_12405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21342_ (.A1(_12405_),
    .A2(net648),
    .ZN(_12406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21343_ (.A1(_12401_),
    .A2(_12406_),
    .A3(net20274),
    .ZN(_12407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21344_ (.A1(net17914),
    .A2(net19326),
    .A3(net17558),
    .ZN(_12408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21345_ (.A1(net18884),
    .A2(net19301),
    .A3(_12178_),
    .ZN(_12409_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21346_ (.A1(_12408_),
    .A2(net18876),
    .A3(_12409_),
    .ZN(_12410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21347_ (.A1(_12174_),
    .A2(net19301),
    .A3(net17327),
    .ZN(_12411_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21348_ (.A1(net17336),
    .A2(net17553),
    .A3(net19325),
    .ZN(_12412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21349_ (.A1(_12411_),
    .A2(_12412_),
    .ZN(_12413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21350_ (.A1(_12413_),
    .A2(net18889),
    .ZN(_12414_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21351_ (.A1(_12410_),
    .A2(_12414_),
    .A3(net20040),
    .ZN(_12415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21352_ (.A1(_12407_),
    .A2(_12415_),
    .ZN(_12416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21353_ (.A1(_12416_),
    .A2(_12198_),
    .B(_12314_),
    .ZN(_12417_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21354_ (.A1(_12308_),
    .A2(_12205_),
    .A3(net19319),
    .ZN(_12418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21355_ (.A1(_12385_),
    .A2(net17325),
    .ZN(_12419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21356_ (.A1(_12418_),
    .A2(_12419_),
    .ZN(_12420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21357_ (.A1(_12420_),
    .A2(net18879),
    .ZN(_12421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21358_ (.A1(_12174_),
    .A2(_12274_),
    .ZN(_12422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21359_ (.A1(_12422_),
    .A2(net19319),
    .A3(_12133_),
    .ZN(_12423_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21360_ (.A1(_12423_),
    .A2(net18893),
    .A3(_12309_),
    .ZN(_12424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21361_ (.A1(_12421_),
    .A2(_12424_),
    .ZN(_12425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21362_ (.A1(_12425_),
    .A2(net20277),
    .ZN(_12426_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21363_ (.A1(net17916),
    .A2(net19328),
    .A3(net17343),
    .ZN(_12427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21364_ (.A1(_12125_),
    .A2(net19315),
    .ZN(_12428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21365_ (.A1(_12427_),
    .A2(net18892),
    .A3(_12428_),
    .ZN(_12429_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21366_ (.A1(_12305_),
    .A2(net17556),
    .B(net19319),
    .ZN(_12430_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21367_ (.A1(_12338_),
    .A2(net19314),
    .A3(net488),
    .ZN(_12431_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21368_ (.A1(_12430_),
    .A2(_12431_),
    .A3(net18879),
    .ZN(_12432_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21369_ (.A1(_12429_),
    .A2(net20040),
    .A3(_12432_),
    .ZN(_12433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21370_ (.A1(_12426_),
    .A2(_12433_),
    .A3(net20442),
    .ZN(_12434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21371_ (.A1(_12417_),
    .A2(_12434_),
    .ZN(_12435_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21372_ (.A1(_12308_),
    .A2(net19307),
    .A3(_12217_),
    .Z(_12436_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21373_ (.A1(_12219_),
    .A2(net19317),
    .A3(net17554),
    .Z(_12437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21374_ (.A1(_12436_),
    .A2(_12437_),
    .B(net18877),
    .ZN(_12438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21375_ (.A1(_12308_),
    .A2(_12203_),
    .A3(net19322),
    .ZN(_12439_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21376_ (.A1(net19321),
    .A2(_15763_[0]),
    .Z(_12440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21377_ (.A1(_12439_),
    .A2(net18896),
    .A3(_12440_),
    .ZN(_12441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21378_ (.A1(_12438_),
    .A2(net20274),
    .A3(_12441_),
    .ZN(_12442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21379_ (.A1(_12381_),
    .A2(net644),
    .ZN(_12443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21380_ (.A1(_15760_[0]),
    .A2(net19301),
    .B(net18875),
    .ZN(_12444_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17371 (.I(_06330_),
    .Z(net17371));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21382_ (.A1(_12443_),
    .A2(_12444_),
    .B(net20274),
    .ZN(_12446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21383_ (.A1(net645),
    .A2(net19338),
    .B(net647),
    .ZN(_12447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21384_ (.A1(_12447_),
    .A2(net18885),
    .ZN(_12448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21385_ (.A1(_12448_),
    .A2(_12309_),
    .A3(net18878),
    .ZN(_12449_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21386_ (.A1(_12446_),
    .A2(_12449_),
    .B(net20442),
    .ZN(_12450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21387_ (.A1(_12442_),
    .A2(_12450_),
    .ZN(_12451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21388_ (.A1(_12391_),
    .A2(_12365_),
    .ZN(_12452_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21389_ (.A1(_12452_),
    .A2(net18875),
    .Z(_12453_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21390_ (.A1(_12137_),
    .A2(_12163_),
    .Z(_12454_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21391_ (.A1(net647),
    .A2(net19336),
    .A3(_12454_),
    .Z(_12455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21392_ (.A1(_12453_),
    .A2(_12349_),
    .A3(_12455_),
    .ZN(_12456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21393_ (.A1(net17329),
    .A2(_12267_),
    .ZN(_12457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21394_ (.I(_12237_),
    .ZN(_12458_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21395_ (.A1(_12458_),
    .A2(net19308),
    .B(net18875),
    .ZN(_12459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21396_ (.A1(_12459_),
    .A2(_12457_),
    .B(net20274),
    .ZN(_12460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21397_ (.A1(_12456_),
    .A2(_12460_),
    .ZN(_12461_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21398_ (.A1(_15767_[0]),
    .A2(net19315),
    .B(net18899),
    .ZN(_12462_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21399_ (.A1(_12418_),
    .A2(_12462_),
    .B(net20040),
    .ZN(_12463_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21400_ (.A1(net19310),
    .A2(_15758_[0]),
    .Z(_12464_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21401_ (.A1(_12428_),
    .A2(net18899),
    .A3(_12464_),
    .ZN(_12465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21402_ (.A1(_12463_),
    .A2(_12465_),
    .ZN(_12466_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21403_ (.A1(net20442),
    .A2(_12466_),
    .A3(_12461_),
    .ZN(_12467_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21404_ (.A1(_12467_),
    .A2(_12451_),
    .A3(_12314_),
    .ZN(_12468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21405_ (.A1(_12468_),
    .A2(_12435_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21406_ (.A1(_12208_),
    .A2(_12219_),
    .Z(_12469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21407_ (.A1(_12447_),
    .A2(_12469_),
    .ZN(_12470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21408_ (.A1(_12365_),
    .A2(net19332),
    .ZN(_12471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21409_ (.A1(_12471_),
    .A2(_12368_),
    .ZN(_12472_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21410_ (.A1(_12470_),
    .A2(_12472_),
    .A3(net18892),
    .Z(_12473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21411_ (.A1(_12228_),
    .A2(net17332),
    .ZN(_12474_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21412_ (.A1(_12474_),
    .A2(_12209_),
    .A3(net648),
    .Z(_12475_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21413_ (.A1(_12475_),
    .A2(_12473_),
    .B(net20041),
    .ZN(_12476_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _21414_ (.A1(_12203_),
    .A2(net18899),
    .A3(_12208_),
    .Z(_12477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21415_ (.A1(net19317),
    .A2(net19332),
    .ZN(_12478_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21416_ (.A1(_12477_),
    .A2(net18872),
    .B(net20040),
    .ZN(_12479_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21417_ (.A1(_12295_),
    .A2(net19301),
    .Z(_12480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21418_ (.A1(_12480_),
    .A2(net17562),
    .ZN(_12481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21419_ (.A1(_12357_),
    .A2(_12481_),
    .ZN(_12482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21420_ (.A1(_12479_),
    .A2(_12482_),
    .B(net20442),
    .ZN(_12483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21421_ (.A1(_12476_),
    .A2(_12483_),
    .ZN(_12484_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21422_ (.A1(_12234_),
    .A2(net648),
    .Z(_12485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21423_ (.A1(net17914),
    .A2(net19302),
    .A3(net18885),
    .ZN(_12486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21424_ (.A1(_12485_),
    .A2(_12486_),
    .B(net20040),
    .ZN(_12487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21425_ (.A1(_12202_),
    .A2(net17917),
    .ZN(_12488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21426_ (.A1(_12267_),
    .A2(net17914),
    .ZN(_12489_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21427_ (.A1(_12489_),
    .A2(_12488_),
    .A3(net18889),
    .ZN(_12490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21428_ (.A1(_12490_),
    .A2(_12487_),
    .B(_12198_),
    .ZN(_12491_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21429_ (.A1(_12469_),
    .A2(net19327),
    .Z(_12492_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21430_ (.I(_12478_),
    .ZN(_12493_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21431_ (.A1(_12493_),
    .A2(net17561),
    .B(net18887),
    .ZN(_12494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21432_ (.I(_12233_),
    .ZN(_12495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21433_ (.A1(_12495_),
    .A2(net19326),
    .Z(_12496_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21434_ (.I(_12496_),
    .ZN(_12497_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21435_ (.A1(_12492_),
    .A2(_12494_),
    .A3(_12497_),
    .ZN(_12498_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21436_ (.A1(net17914),
    .A2(net19301),
    .A3(net17563),
    .ZN(_12499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21437_ (.A1(net17343),
    .A2(net17330),
    .A3(net19327),
    .ZN(_12500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21438_ (.A1(_12499_),
    .A2(net18890),
    .A3(_12500_),
    .ZN(_12501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21439_ (.A1(_12498_),
    .A2(net20040),
    .A3(_12501_),
    .ZN(_12502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21440_ (.A1(_12502_),
    .A2(_12491_),
    .ZN(_12503_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21441_ (.A1(_12503_),
    .A2(_12314_),
    .A3(_12484_),
    .ZN(_12504_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21442_ (.I(_12264_),
    .ZN(_12505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21443_ (.A1(net19326),
    .A2(net17322),
    .B(net20274),
    .ZN(_12506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21444_ (.A1(_12506_),
    .A2(_12411_),
    .B(net648),
    .ZN(_12507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21445_ (.A1(_12170_),
    .A2(net17336),
    .ZN(_12508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21446_ (.A1(_12454_),
    .A2(net19330),
    .ZN(_12509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21447_ (.A1(_12509_),
    .A2(net19322),
    .ZN(_12510_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21448_ (.I(_12354_),
    .ZN(_12511_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21449_ (.A1(_12510_),
    .A2(_12511_),
    .Z(_12512_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21450_ (.A1(_12508_),
    .A2(_12512_),
    .A3(net20274),
    .ZN(_12513_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21451_ (.A1(_12507_),
    .A2(_12513_),
    .B(_12198_),
    .ZN(_12514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21452_ (.A1(net17923),
    .A2(net17331),
    .B(net19326),
    .ZN(_12515_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21453_ (.A1(_12515_),
    .A2(_12496_),
    .B(net20274),
    .ZN(_12516_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21454_ (.I(_12232_),
    .ZN(_12517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21455_ (.A1(_12517_),
    .A2(net20040),
    .B1(net19326),
    .B2(net17341),
    .ZN(_12518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21456_ (.A1(_12516_),
    .A2(_12518_),
    .ZN(_12519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21457_ (.A1(_12519_),
    .A2(net18876),
    .ZN(_12520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21458_ (.A1(_12514_),
    .A2(_12520_),
    .B(_12314_),
    .ZN(_12521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21459_ (.A1(_12296_),
    .A2(net17224),
    .ZN(_12522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21460_ (.A1(_12522_),
    .A2(_12349_),
    .B(net648),
    .ZN(_12523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21461_ (.A1(_12409_),
    .A2(net18876),
    .ZN(_12524_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21462_ (.I(_12524_),
    .ZN(_12525_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21463_ (.A1(_12523_),
    .A2(_12525_),
    .B(net20274),
    .ZN(_12526_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21464_ (.A1(net18317),
    .A2(_12505_),
    .B(net19319),
    .ZN(_12527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21465_ (.A1(_12179_),
    .A2(net19314),
    .ZN(_12528_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21466_ (.A1(_12527_),
    .A2(net18879),
    .A3(_12528_),
    .ZN(_12529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21467_ (.A1(_12272_),
    .A2(_12393_),
    .ZN(_12530_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21468_ (.A1(_12529_),
    .A2(_12530_),
    .A3(net20041),
    .ZN(_12531_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21469_ (.A1(_12526_),
    .A2(_12531_),
    .A3(_12198_),
    .ZN(_12532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21470_ (.A1(_12521_),
    .A2(_12532_),
    .ZN(_12533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21471_ (.A1(_12504_),
    .A2(_12533_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21472_ (.A1(_12332_),
    .A2(net19303),
    .Z(_12534_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21473_ (.A1(_12534_),
    .A2(net18897),
    .ZN(_12535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21474_ (.A1(_12225_),
    .A2(net19322),
    .ZN(_12536_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21475_ (.A1(_12535_),
    .A2(_12536_),
    .B(net20275),
    .ZN(_12537_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21476_ (.A1(_12385_),
    .A2(net17555),
    .B(net18875),
    .ZN(_12538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21477_ (.A1(_12538_),
    .A2(_12146_),
    .ZN(_12539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21478_ (.A1(_12537_),
    .A2(_12539_),
    .ZN(_12540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21479_ (.A1(_12202_),
    .A2(net17324),
    .ZN(_12541_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21480_ (.A1(_12391_),
    .A2(net18875),
    .ZN(_12542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21481_ (.A1(_12541_),
    .A2(_12542_),
    .B(net20040),
    .ZN(_12543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21482_ (.A1(_12458_),
    .A2(net647),
    .B(net18894),
    .ZN(_12544_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21483_ (.A1(_12317_),
    .A2(_12544_),
    .A3(net17921),
    .ZN(_12545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21484_ (.A1(_12543_),
    .A2(_12545_),
    .ZN(_12546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21485_ (.A1(_12540_),
    .A2(_12546_),
    .ZN(_12547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21486_ (.A1(_12547_),
    .A2(_12198_),
    .ZN(_12548_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21487_ (.A1(net436),
    .A2(net18884),
    .B(net19317),
    .ZN(_12549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21488_ (.A1(_12296_),
    .A2(_12133_),
    .ZN(_12550_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21489_ (.I(_12550_),
    .ZN(_12551_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21490_ (.A1(_12549_),
    .A2(_12551_),
    .B(net18877),
    .ZN(_12552_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21491_ (.A1(_15751_[0]),
    .A2(net19306),
    .B(net648),
    .ZN(_12553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21492_ (.A1(_12280_),
    .A2(net19318),
    .ZN(_12554_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21493_ (.A1(_12553_),
    .A2(_12554_),
    .B(net20274),
    .ZN(_12555_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21494_ (.A1(_12552_),
    .A2(_12555_),
    .B(_12198_),
    .ZN(_12556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21495_ (.A1(_12303_),
    .A2(_12209_),
    .A3(_12293_),
    .ZN(_12557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21496_ (.A1(_12205_),
    .A2(_12316_),
    .A3(net19313),
    .ZN(_12558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21497_ (.A1(_12296_),
    .A2(net18884),
    .ZN(_12559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21498_ (.A1(_12558_),
    .A2(_12559_),
    .A3(net648),
    .ZN(_12560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21499_ (.A1(_12560_),
    .A2(_12557_),
    .ZN(_12561_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21500_ (.A1(net20274),
    .A2(_12561_),
    .ZN(_12562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21501_ (.A1(_12556_),
    .A2(_12562_),
    .ZN(_12563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21502_ (.A1(_12563_),
    .A2(_12548_),
    .ZN(_12564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21503_ (.A1(_12564_),
    .A2(net20637),
    .ZN(_12565_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21504_ (.A1(_12377_),
    .A2(net17226),
    .B(net18887),
    .ZN(_12566_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21505_ (.A1(_12422_),
    .A2(net19307),
    .A3(_12133_),
    .Z(_12567_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21506_ (.A1(_12566_),
    .A2(_12567_),
    .ZN(_12568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21507_ (.A1(_12447_),
    .A2(_12273_),
    .ZN(_12569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21508_ (.A1(_12569_),
    .A2(_12419_),
    .B(net18893),
    .ZN(_12570_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21509_ (.A1(_12568_),
    .A2(_12570_),
    .B(net20277),
    .ZN(_12571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21510_ (.A1(_12554_),
    .A2(net17557),
    .Z(_12572_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21511_ (.A1(_12572_),
    .A2(_12379_),
    .B(net20274),
    .ZN(_12573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21512_ (.A1(_12331_),
    .A2(net17335),
    .ZN(_12574_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21513_ (.A1(_12574_),
    .A2(_12297_),
    .A3(net18888),
    .ZN(_12575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21514_ (.A1(_12573_),
    .A2(_12575_),
    .B(_12198_),
    .ZN(_12576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21515_ (.A1(_12576_),
    .A2(_12571_),
    .ZN(_12577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21516_ (.A1(_12439_),
    .A2(_12339_),
    .A3(net18896),
    .ZN(_12578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21517_ (.A1(net17913),
    .A2(net17924),
    .A3(net19311),
    .ZN(_12579_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21518_ (.A1(net17924),
    .A2(net19323),
    .A3(_12241_),
    .ZN(_12580_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21519_ (.A1(_12579_),
    .A2(_12580_),
    .A3(net18881),
    .ZN(_12581_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21520_ (.A1(_12578_),
    .A2(_12581_),
    .A3(net20275),
    .ZN(_12582_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21521_ (.A1(_12338_),
    .A2(net19322),
    .A3(_12174_),
    .ZN(_12583_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21522_ (.A1(_12583_),
    .A2(net18896),
    .A3(_12344_),
    .ZN(_12584_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21523_ (.I(net17229),
    .ZN(_12585_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21524_ (.A1(net17342),
    .A2(net18896),
    .ZN(_12586_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21525_ (.A1(_12585_),
    .A2(_12586_),
    .B(net20275),
    .ZN(_12587_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21526_ (.A1(_12584_),
    .A2(_12587_),
    .B(net20442),
    .ZN(_12588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21527_ (.A1(_12582_),
    .A2(_12588_),
    .ZN(_12589_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21528_ (.A1(_12577_),
    .A2(net20440),
    .A3(_12589_),
    .ZN(_12590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21529_ (.A1(_12565_),
    .A2(_12590_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21530_ (.A1(_12471_),
    .A2(net19328),
    .A3(_12238_),
    .ZN(_12591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21531_ (.A1(_12170_),
    .A2(_12365_),
    .ZN(_12592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21532_ (.A1(_12592_),
    .A2(_12591_),
    .ZN(_12593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21533_ (.A1(net20040),
    .A2(_12593_),
    .ZN(_12594_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21534_ (.A1(_12554_),
    .A2(net20274),
    .Z(_12595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21535_ (.A1(_12534_),
    .A2(net17915),
    .ZN(_12596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21536_ (.A1(_12595_),
    .A2(_12596_),
    .B(net18896),
    .ZN(_12597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21537_ (.A1(_12594_),
    .A2(_12597_),
    .ZN(_12598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21538_ (.A1(_12178_),
    .A2(net19305),
    .ZN(_12599_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21539_ (.A1(_12301_),
    .A2(net17230),
    .B(net20274),
    .C(_12599_),
    .ZN(_12600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21540_ (.A1(net18315),
    .A2(net19321),
    .B(_12160_),
    .ZN(_12601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21541_ (.A1(_12601_),
    .A2(_12558_),
    .ZN(_12602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21542_ (.A1(_12602_),
    .A2(_12600_),
    .ZN(_12603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21543_ (.A1(_12603_),
    .A2(net18895),
    .ZN(_12604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21544_ (.A1(_12604_),
    .A2(net20442),
    .A3(_12598_),
    .ZN(_12605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21545_ (.A1(_12356_),
    .A2(net17339),
    .ZN(_12606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21546_ (.A1(_12144_),
    .A2(_12606_),
    .ZN(_12607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21547_ (.A1(net644),
    .A2(_12480_),
    .ZN(_12608_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21548_ (.A1(net17607),
    .A2(net19317),
    .B(net18887),
    .ZN(_12609_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21549_ (.A1(_12608_),
    .A2(_12609_),
    .A3(_12287_),
    .ZN(_12610_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21550_ (.A1(_12607_),
    .A2(_12610_),
    .A3(net20040),
    .ZN(_12611_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21551_ (.A1(_12228_),
    .A2(net18875),
    .ZN(_12612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21552_ (.A1(_12612_),
    .A2(_12527_),
    .ZN(_12613_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21553_ (.A1(net17227),
    .A2(net18899),
    .ZN(_12614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21554_ (.A1(net18873),
    .A2(_12205_),
    .ZN(_12615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21555_ (.A1(_12614_),
    .A2(_12615_),
    .ZN(_12616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21556_ (.A1(_12613_),
    .A2(_12616_),
    .A3(net20275),
    .ZN(_12617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21557_ (.A1(_12617_),
    .A2(_12198_),
    .A3(_12611_),
    .ZN(_12618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21558_ (.A1(_12605_),
    .A2(_12618_),
    .A3(net20440),
    .ZN(_12619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21559_ (.A1(net17919),
    .A2(net19312),
    .ZN(_12620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21560_ (.A1(_12306_),
    .A2(net19322),
    .ZN(_12621_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21561_ (.A1(_12620_),
    .A2(net17223),
    .B(net18880),
    .C(_12621_),
    .ZN(_12622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21562_ (.A1(_12305_),
    .A2(net19304),
    .ZN(_12623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21563_ (.A1(_12146_),
    .A2(_12262_),
    .A3(_12623_),
    .ZN(_12624_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21564_ (.A1(_12622_),
    .A2(_12624_),
    .A3(net20274),
    .ZN(_12625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21565_ (.A1(net19340),
    .A2(net19322),
    .B(net18875),
    .ZN(_12626_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21566_ (.A1(_12204_),
    .A2(_12626_),
    .B(net20275),
    .ZN(_12627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21567_ (.A1(_12267_),
    .A2(net17926),
    .ZN(_12628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21568_ (.A1(_12480_),
    .A2(net642),
    .ZN(_12629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21569_ (.A1(_12628_),
    .A2(net648),
    .A3(_12629_),
    .ZN(_12630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21570_ (.A1(_12630_),
    .A2(_12627_),
    .B(net20442),
    .ZN(_12631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21571_ (.A1(_12631_),
    .A2(_12625_),
    .ZN(_12632_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21572_ (.I(_12177_),
    .ZN(_12633_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21573_ (.A1(_12633_),
    .A2(_12511_),
    .A3(net19322),
    .Z(_12634_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21574_ (.A1(_12267_),
    .A2(net17552),
    .ZN(_12635_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21575_ (.A1(_12635_),
    .A2(net18880),
    .A3(_12634_),
    .ZN(_12636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21576_ (.A1(net17560),
    .A2(net19322),
    .B(net18875),
    .ZN(_12637_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21577_ (.A1(_12620_),
    .A2(_12637_),
    .B(net20040),
    .ZN(_12638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21578_ (.A1(_12636_),
    .A2(_12638_),
    .ZN(_12639_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21579_ (.I(net17919),
    .ZN(_12640_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21580_ (.A1(_12510_),
    .A2(net18896),
    .Z(_12641_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21581_ (.A1(_12428_),
    .A2(_12640_),
    .B(_12641_),
    .ZN(_12642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21582_ (.A1(_12379_),
    .A2(net17228),
    .B(net20275),
    .ZN(_12643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21583_ (.A1(_12642_),
    .A2(_12643_),
    .ZN(_12644_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21584_ (.A1(net20442),
    .A2(_12644_),
    .A3(_12639_),
    .ZN(_12645_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21585_ (.A1(_12645_),
    .A2(_12632_),
    .A3(net20637),
    .ZN(_12646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21586_ (.A1(_12646_),
    .A2(_12619_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21587_ (.A1(_12125_),
    .A2(net19315),
    .A3(net17338),
    .ZN(_12647_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21588_ (.A1(_12647_),
    .A2(net648),
    .A3(_12464_),
    .ZN(_12648_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21589_ (.A1(net17926),
    .A2(net19324),
    .A3(net17924),
    .ZN(_12649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21590_ (.A1(net17222),
    .A2(net17563),
    .ZN(_12650_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21591_ (.A1(_12649_),
    .A2(net18894),
    .A3(_12650_),
    .ZN(_12651_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21592_ (.A1(_12648_),
    .A2(_12651_),
    .A3(net20040),
    .ZN(_12652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21593_ (.A1(_12306_),
    .A2(net19308),
    .B(net18898),
    .ZN(_12653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21594_ (.A1(net18883),
    .A2(net641),
    .ZN(_12654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21595_ (.A1(_12654_),
    .A2(net19322),
    .ZN(_12655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21596_ (.A1(_12653_),
    .A2(_12655_),
    .B(net20040),
    .ZN(_12656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21597_ (.A1(_12368_),
    .A2(net17225),
    .B(net18875),
    .ZN(_12657_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21598_ (.A1(_12273_),
    .A2(net19324),
    .A3(net18882),
    .ZN(_12658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21599_ (.A1(_12658_),
    .A2(_12657_),
    .ZN(_12659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21600_ (.A1(_12656_),
    .A2(_12659_),
    .B(_12198_),
    .ZN(_12660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21601_ (.A1(_12660_),
    .A2(_12652_),
    .ZN(_12661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21602_ (.A1(net19335),
    .A2(net17608),
    .ZN(_12662_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _21603_ (.A1(net19318),
    .A2(_12259_),
    .A3(_12662_),
    .A4(net17557),
    .ZN(_12663_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21604_ (.A1(_12663_),
    .A2(_12282_),
    .A3(_12623_),
    .ZN(_12664_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21605_ (.A1(_12055_),
    .A2(net17327),
    .A3(net19301),
    .ZN(_12665_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21606_ (.A1(_12452_),
    .A2(_12287_),
    .A3(_12665_),
    .ZN(_12666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21607_ (.A1(_12666_),
    .A2(net18891),
    .ZN(_12667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21608_ (.A1(_12664_),
    .A2(_12667_),
    .ZN(_12668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21609_ (.A1(_12668_),
    .A2(net20274),
    .ZN(_12669_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21610_ (.A1(net17556),
    .A2(net17323),
    .B(net19319),
    .ZN(_12670_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21611_ (.A1(_12544_),
    .A2(_12670_),
    .B(net20275),
    .ZN(_12671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21612_ (.A1(_12447_),
    .A2(net17917),
    .ZN(_12672_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21613_ (.A1(_15756_[0]),
    .A2(_15765_[0]),
    .B(net647),
    .ZN(_12673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21614_ (.A1(_12672_),
    .A2(net18897),
    .A3(_12673_),
    .ZN(_12674_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21615_ (.A1(_12674_),
    .A2(_12671_),
    .B(net20442),
    .ZN(_12675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21616_ (.A1(_12669_),
    .A2(_12675_),
    .ZN(_12676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21617_ (.A1(_12676_),
    .A2(_12661_),
    .A3(net20441),
    .ZN(_12677_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21618_ (.A1(net19329),
    .A2(net17606),
    .Z(_12678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21619_ (.A1(net18317),
    .A2(_12678_),
    .B(net19308),
    .ZN(_12679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21620_ (.A1(net17918),
    .A2(net19324),
    .A3(net18882),
    .ZN(_12680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21621_ (.A1(_12679_),
    .A2(_12680_),
    .A3(net648),
    .ZN(_12681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21622_ (.A1(net645),
    .A2(net19309),
    .ZN(_12682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21623_ (.A1(_12477_),
    .A2(net17911),
    .ZN(_12683_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21624_ (.A1(_12681_),
    .A2(_12683_),
    .A3(net20040),
    .ZN(_12684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21625_ (.A1(net17321),
    .A2(net19308),
    .B(net18875),
    .ZN(_12685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21626_ (.A1(_12527_),
    .A2(_12685_),
    .B(net20040),
    .ZN(_12686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21627_ (.A1(_12377_),
    .A2(net18875),
    .Z(_12687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21628_ (.A1(_12176_),
    .A2(_12687_),
    .ZN(_12688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21629_ (.A1(_12686_),
    .A2(_12688_),
    .ZN(_12689_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21630_ (.A1(_12684_),
    .A2(_12198_),
    .A3(_12689_),
    .ZN(_12690_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21631_ (.A1(_12551_),
    .A2(net17328),
    .B(net18877),
    .ZN(_12691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21632_ (.A1(_12423_),
    .A2(net18887),
    .ZN(_12692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21633_ (.A1(_12691_),
    .A2(_12692_),
    .ZN(_12693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21634_ (.A1(_12693_),
    .A2(net20276),
    .ZN(_12694_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21635_ (.A1(net17321),
    .A2(net17228),
    .B(_12324_),
    .C(net648),
    .ZN(_12695_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21636_ (.I(_15757_[0]),
    .ZN(_12696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21637_ (.A1(_12696_),
    .A2(net19323),
    .B(net18875),
    .ZN(_12697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21638_ (.A1(_12697_),
    .A2(_12629_),
    .B(net20275),
    .ZN(_12698_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21639_ (.A1(_12695_),
    .A2(_12698_),
    .B(_12198_),
    .ZN(_12699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21640_ (.A1(_12694_),
    .A2(_12699_),
    .ZN(_12700_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21641_ (.A1(_12690_),
    .A2(_12700_),
    .A3(net20637),
    .ZN(_12701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21642_ (.A1(_12701_),
    .A2(_12677_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21643_ (.A1(net18894),
    .A2(_12237_),
    .Z(_12702_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21644_ (.A1(_12277_),
    .A2(_12702_),
    .Z(_12703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21645_ (.A1(net18873),
    .A2(net645),
    .ZN(_12704_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21646_ (.A1(_12704_),
    .A2(_12703_),
    .B(net20040),
    .ZN(_12705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21647_ (.A1(net19312),
    .A2(net17607),
    .ZN(_12706_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21648_ (.A1(_12672_),
    .A2(_12706_),
    .A3(net648),
    .ZN(_12707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21649_ (.A1(_12707_),
    .A2(_12705_),
    .B(net20442),
    .ZN(_12708_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21650_ (.A1(net19303),
    .A2(net19334),
    .Z(_12709_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21651_ (.A1(_12709_),
    .A2(net19338),
    .Z(_12710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21652_ (.A1(_12682_),
    .A2(net648),
    .ZN(_12711_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21653_ (.A1(_12710_),
    .A2(_12711_),
    .ZN(_12712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21654_ (.A1(_12522_),
    .A2(_12712_),
    .B(net20275),
    .ZN(_12713_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21655_ (.A1(_12710_),
    .A2(_12143_),
    .ZN(_12714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21656_ (.A1(net17552),
    .A2(net17563),
    .A3(net19322),
    .ZN(_12715_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21657_ (.A1(_12714_),
    .A2(_12459_),
    .A3(_12715_),
    .ZN(_12716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21658_ (.A1(_12713_),
    .A2(_12716_),
    .ZN(_12717_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21659_ (.A1(_12717_),
    .A2(_12708_),
    .ZN(_12718_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21660_ (.A1(_12505_),
    .A2(net19301),
    .Z(_12719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21661_ (.A1(net19327),
    .A2(_15765_[0]),
    .ZN(_12720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21662_ (.A1(_12720_),
    .A2(net18890),
    .ZN(_12721_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21663_ (.A1(_12719_),
    .A2(_12721_),
    .ZN(_12722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21664_ (.A1(_12495_),
    .A2(net19301),
    .ZN(_12723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21665_ (.A1(_12722_),
    .A2(_12723_),
    .B(net20040),
    .ZN(_12724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21666_ (.A1(_12170_),
    .A2(net17922),
    .ZN(_12725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21667_ (.A1(_12381_),
    .A2(net17563),
    .ZN(_12726_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21668_ (.A1(_12725_),
    .A2(_12726_),
    .A3(net648),
    .ZN(_12727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21669_ (.A1(_12724_),
    .A2(_12727_),
    .ZN(_12728_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21670_ (.I(_15751_[0]),
    .ZN(_12729_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21671_ (.A1(_12729_),
    .A2(net19320),
    .B(net18875),
    .ZN(_12730_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21672_ (.A1(_12730_),
    .A2(_12277_),
    .B(net20275),
    .ZN(_12731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21673_ (.A1(_12654_),
    .A2(net19308),
    .ZN(_12732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21674_ (.A1(_12317_),
    .A2(net648),
    .A3(_12732_),
    .ZN(_12733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21675_ (.A1(_12731_),
    .A2(_12733_),
    .ZN(_12734_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21676_ (.A1(_12728_),
    .A2(net20442),
    .A3(_12734_),
    .ZN(_12735_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21677_ (.A1(_12735_),
    .A2(net20441),
    .A3(_12718_),
    .ZN(_12736_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _21678_ (.A1(_12331_),
    .A2(net18877),
    .ZN(_12737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21679_ (.A1(net17202),
    .A2(_12737_),
    .B(net20442),
    .ZN(_12738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21680_ (.A1(_12170_),
    .A2(_12273_),
    .ZN(_12739_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21681_ (.A1(_12494_),
    .A2(_12739_),
    .A3(net17551),
    .ZN(_12740_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21682_ (.A1(_12740_),
    .A2(_12738_),
    .B(net20276),
    .ZN(_12741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21683_ (.A1(_12225_),
    .A2(net19311),
    .A3(net17924),
    .ZN(_12742_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21684_ (.A1(_12742_),
    .A2(net18894),
    .A3(_12439_),
    .ZN(_12743_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21685_ (.I(_12709_),
    .ZN(_12744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21686_ (.A1(_12583_),
    .A2(_12744_),
    .ZN(_12745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21687_ (.A1(_12745_),
    .A2(net18881),
    .ZN(_12746_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21688_ (.A1(_12743_),
    .A2(_12746_),
    .A3(net20442),
    .ZN(_12747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21689_ (.A1(_12747_),
    .A2(_12741_),
    .ZN(_12748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21690_ (.A1(_12232_),
    .A2(net18889),
    .Z(_12749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21691_ (.A1(net18313),
    .A2(net17912),
    .ZN(_12750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21692_ (.A1(_12749_),
    .A2(_12750_),
    .B(_12198_),
    .ZN(_12751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21693_ (.A1(net644),
    .A2(net19327),
    .B(net18889),
    .ZN(_12752_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21694_ (.A1(net17916),
    .A2(net19301),
    .A3(net17563),
    .ZN(_12753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21695_ (.A1(_12752_),
    .A2(_12753_),
    .ZN(_12754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21696_ (.A1(_12751_),
    .A2(_12754_),
    .B(net20040),
    .ZN(_12755_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21697_ (.A1(_12508_),
    .A2(_12382_),
    .A3(net18878),
    .ZN(_12756_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21698_ (.A1(_12448_),
    .A2(net18889),
    .A3(net17221),
    .ZN(_12757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21699_ (.A1(_12198_),
    .A2(_12757_),
    .A3(_12756_),
    .ZN(_12758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21700_ (.A1(_12755_),
    .A2(_12758_),
    .ZN(_12759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21701_ (.A1(_12748_),
    .A2(_12759_),
    .A3(net20637),
    .ZN(_12760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21702_ (.A1(_12760_),
    .A2(_12736_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21703_ (.I(\sa03_sr[7] ),
    .ZN(_12761_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21704_ (.I(\sa03_sr[0] ),
    .ZN(_12762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21705_ (.A1(_12762_),
    .A2(_12761_),
    .ZN(_12763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21706_ (.A1(net21433),
    .A2(\sa03_sr[0] ),
    .ZN(_12764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21707_ (.A1(_12764_),
    .A2(_12763_),
    .ZN(_12765_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21708_ (.I(\sa32_sub[1] ),
    .ZN(_12766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21709_ (.A1(_12766_),
    .A2(net21327),
    .ZN(_12767_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21710_ (.I(\sa21_sub[1] ),
    .ZN(_12768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21711_ (.A1(_12768_),
    .A2(net21269),
    .ZN(_12769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21712_ (.A1(_12769_),
    .A2(_12767_),
    .ZN(_12770_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21713_ (.A1(_12770_),
    .A2(_12765_),
    .ZN(_12771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21714_ (.A1(net21433),
    .A2(_12762_),
    .ZN(_12772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21715_ (.A1(_12761_),
    .A2(\sa03_sr[0] ),
    .ZN(_12773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21716_ (.A1(_12773_),
    .A2(_12772_),
    .ZN(_12774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21717_ (.A1(_12768_),
    .A2(_12766_),
    .ZN(_12775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21718_ (.A1(net21326),
    .A2(net21269),
    .ZN(_12776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21719_ (.A1(_12776_),
    .A2(_12775_),
    .ZN(_12777_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21720_ (.A1(_12777_),
    .A2(_12774_),
    .ZN(_12778_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21721_ (.A1(_12778_),
    .A2(_12771_),
    .ZN(_12779_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _21722_ (.I(\sa10_sub[0] ),
    .ZN(_12780_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17542 (.I(_13196_),
    .Z(net17542));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21724_ (.A1(net21006),
    .A2(net21374),
    .ZN(_12782_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21725_ (.I(\sa10_sub[7] ),
    .ZN(_12783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21726_ (.A1(_12783_),
    .A2(net21383),
    .ZN(_12784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21727_ (.A1(_12782_),
    .A2(_12784_),
    .ZN(_12785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21728_ (.A1(_12785_),
    .A2(net21382),
    .ZN(_12786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21729_ (.A1(_12783_),
    .A2(net21006),
    .ZN(_12787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21730_ (.A1(net21374),
    .A2(net21383),
    .ZN(_12788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21731_ (.A1(_12787_),
    .A2(_12788_),
    .ZN(_12789_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21732_ (.I(\sa10_sub[1] ),
    .ZN(_12790_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21733_ (.A1(_12789_),
    .A2(net21003),
    .ZN(_12791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21734_ (.A1(_12786_),
    .A2(_12791_),
    .ZN(_12792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21735_ (.A1(_12792_),
    .A2(_12779_),
    .ZN(_12793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21736_ (.A1(_12774_),
    .A2(_12777_),
    .ZN(_12794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21737_ (.A1(_12765_),
    .A2(_12770_),
    .ZN(_12795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21738_ (.A1(_12794_),
    .A2(_12795_),
    .ZN(_12796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21739_ (.A1(_12789_),
    .A2(net21382),
    .ZN(_12797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21740_ (.A1(_12785_),
    .A2(net21003),
    .ZN(_12798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21741_ (.A1(_12797_),
    .A2(_12798_),
    .ZN(_12799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21742_ (.A1(_12796_),
    .A2(_12799_),
    .ZN(_12800_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21743_ (.A1(_12800_),
    .A2(_12793_),
    .A3(_10378_),
    .ZN(_12801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21744_ (.A1(net21486),
    .A2(\text_in_r[25] ),
    .ZN(_12802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21745_ (.A1(_12802_),
    .A2(_12801_),
    .ZN(_12803_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21746_ (.I(net21144),
    .ZN(_12804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21747_ (.A1(net20039),
    .A2(_12804_),
    .ZN(_12805_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21748_ (.A1(net20272),
    .A2(net21144),
    .A3(_12802_),
    .ZN(_12806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21749_ (.A1(_12805_),
    .A2(_12806_),
    .ZN(_15775_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21750_ (.A1(net21012),
    .A2(_12783_),
    .ZN(_12807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21751_ (.A1(net21436),
    .A2(net21375),
    .ZN(_12808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21752_ (.A1(_12807_),
    .A2(_12808_),
    .ZN(_12809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21753_ (.A1(_12809_),
    .A2(net21272),
    .ZN(_12810_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21754_ (.I(\sa32_sub[0] ),
    .ZN(_12811_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21755_ (.A1(_12807_),
    .A2(net21002),
    .A3(_12808_),
    .ZN(_12812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21756_ (.A1(_12810_),
    .A2(_12812_),
    .ZN(_12813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21757_ (.A1(net21331),
    .A2(net21007),
    .ZN(_12814_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21758_ (.I(\sa21_sub[0] ),
    .ZN(_12815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21759_ (.A1(net21383),
    .A2(net21001),
    .ZN(_12816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21760_ (.A1(net414),
    .A2(_12816_),
    .ZN(_12817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21761_ (.A1(_12813_),
    .A2(_12817_),
    .ZN(_12818_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21762_ (.I(_12817_),
    .ZN(_12819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21763_ (.A1(_12810_),
    .A2(_12812_),
    .A3(_12819_),
    .ZN(_12820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21764_ (.A1(_12818_),
    .A2(_12820_),
    .B(net21486),
    .ZN(_12821_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21765_ (.I(\text_in_r[24] ),
    .ZN(_12822_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21766_ (.A1(_12822_),
    .A2(net21486),
    .Z(_12823_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21767_ (.A1(net20945),
    .A2(net419),
    .B(net21145),
    .ZN(_12824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21768_ (.A1(_12818_),
    .A2(_12820_),
    .ZN(_12825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21769_ (.A1(_12825_),
    .A2(net21094),
    .ZN(_12826_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21770_ (.I(net21145),
    .ZN(_12827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21771_ (.I(_12823_),
    .ZN(_12828_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21772_ (.A1(_12826_),
    .A2(_12827_),
    .A3(_12828_),
    .ZN(_12829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21773_ (.A1(_12824_),
    .A2(_12829_),
    .ZN(_15778_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21774_ (.I(\sa03_sr[1] ),
    .ZN(_12830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21775_ (.A1(_12830_),
    .A2(_12790_),
    .ZN(_12831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21776_ (.A1(net21442),
    .A2(\sa10_sub[1] ),
    .ZN(_12832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21777_ (.A1(_12831_),
    .A2(_12832_),
    .ZN(_12833_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _21778_ (.I(\sa21_sub[2] ),
    .ZN(_12834_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21779_ (.A1(net20891),
    .A2(net20999),
    .ZN(_12835_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17366 (.I(_06829_),
    .Z(net17366));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21781_ (.A1(net20944),
    .A2(net21325),
    .A3(net21000),
    .ZN(_12837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21782_ (.A1(_12835_),
    .A2(_12837_),
    .ZN(_12838_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _21783_ (.I(\sa32_sub[2] ),
    .ZN(_12839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21784_ (.A1(_12839_),
    .A2(net21381),
    .ZN(_12840_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _21785_ (.I(\sa10_sub[2] ),
    .ZN(_12841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21786_ (.A1(_12841_),
    .A2(\sa32_sub[2] ),
    .ZN(_12842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21787_ (.A1(net20943),
    .A2(net20942),
    .ZN(_12843_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21788_ (.I(_12843_),
    .ZN(_12844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21789_ (.A1(_12838_),
    .A2(_12844_),
    .ZN(_12845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21790_ (.A1(_12835_),
    .A2(_12837_),
    .A3(_12843_),
    .ZN(_12846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21791_ (.A1(_12845_),
    .A2(_12846_),
    .B(net21486),
    .ZN(_12847_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21792_ (.I(\text_in_r[26] ),
    .ZN(_12848_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21793_ (.A1(_12848_),
    .A2(net21486),
    .Z(_12849_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21794_ (.I(net21143),
    .ZN(_12850_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21795_ (.A1(_12847_),
    .A2(_12849_),
    .B(_12850_),
    .ZN(_12851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21796_ (.A1(_12845_),
    .A2(_12846_),
    .ZN(_12852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21797_ (.A1(_12852_),
    .A2(net21094),
    .ZN(_12853_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21798_ (.I(_12849_),
    .ZN(_12854_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21799_ (.A1(_12853_),
    .A2(net21143),
    .A3(_12854_),
    .ZN(_12855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21800_ (.A1(_12851_),
    .A2(_12855_),
    .ZN(_12856_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17369 (.I(_06422_),
    .Z(net17369));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21802_ (.A1(_12823_),
    .A2(_12821_),
    .B(_12827_),
    .ZN(_12857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21803_ (.A1(_12826_),
    .A2(net21145),
    .A3(_12828_),
    .ZN(_12858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21804_ (.A1(_12858_),
    .A2(_12857_),
    .ZN(_15769_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21805_ (.A1(_12847_),
    .A2(_12849_),
    .B(net21143),
    .ZN(_12859_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21806_ (.A1(_12853_),
    .A2(_12850_),
    .A3(_12854_),
    .ZN(_12860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21807_ (.A1(_12859_),
    .A2(_12860_),
    .ZN(_12861_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17359 (.I(_07088_),
    .Z(net17359));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17361 (.I(_07027_),
    .Z(net17361));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21810_ (.A1(net19298),
    .A2(net19293),
    .A3(net19286),
    .ZN(_12863_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21811_ (.I(\sa03_sr[2] ),
    .ZN(_12864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21812_ (.A1(net21011),
    .A2(_12864_),
    .ZN(_12865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21813_ (.A1(net21435),
    .A2(net21440),
    .ZN(_12866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21814_ (.A1(_12865_),
    .A2(_12866_),
    .ZN(_12867_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21815_ (.I(\sa32_sub[3] ),
    .ZN(_12868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21816_ (.A1(_12868_),
    .A2(net21323),
    .ZN(_12869_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21817_ (.I(\sa21_sub[3] ),
    .ZN(_12870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21818_ (.A1(_12870_),
    .A2(net21265),
    .ZN(_12871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21819_ (.A1(_12869_),
    .A2(_12871_),
    .ZN(_12872_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21820_ (.A1(_12867_),
    .A2(_12872_),
    .ZN(_12873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21821_ (.A1(_12864_),
    .A2(net21435),
    .ZN(_12874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21822_ (.A1(net21011),
    .A2(net21440),
    .ZN(_12875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21823_ (.A1(_12874_),
    .A2(_12875_),
    .ZN(_12876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21824_ (.A1(_12870_),
    .A2(_12868_),
    .ZN(_12877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21825_ (.A1(\sa21_sub[3] ),
    .A2(\sa32_sub[3] ),
    .ZN(_12878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21826_ (.A1(_12877_),
    .A2(_12878_),
    .ZN(_12879_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21827_ (.A1(_12876_),
    .A2(_12879_),
    .ZN(_12880_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21828_ (.A1(_12873_),
    .A2(_12880_),
    .ZN(_12881_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21829_ (.I(\sa10_sub[3] ),
    .ZN(_12882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21830_ (.A1(net20991),
    .A2(net21373),
    .ZN(_12883_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21831_ (.A1(net21004),
    .A2(net21379),
    .ZN(_12884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21832_ (.A1(_12883_),
    .A2(_12884_),
    .ZN(_12885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21833_ (.A1(_12885_),
    .A2(net21380),
    .ZN(_12886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21834_ (.A1(net21004),
    .A2(_12882_),
    .ZN(_12887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21835_ (.A1(net21373),
    .A2(net21379),
    .ZN(_12888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21836_ (.A1(_12887_),
    .A2(_12888_),
    .ZN(_12889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21837_ (.A1(_12889_),
    .A2(net20996),
    .ZN(_12890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21838_ (.A1(_12886_),
    .A2(_12890_),
    .ZN(_12891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21839_ (.A1(_12881_),
    .A2(_12891_),
    .ZN(_12892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21840_ (.A1(_12876_),
    .A2(_12879_),
    .ZN(_12893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21841_ (.A1(_12867_),
    .A2(_12872_),
    .ZN(_12894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21842_ (.A1(_12893_),
    .A2(_12894_),
    .ZN(_12895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21843_ (.A1(net21004),
    .A2(net20996),
    .ZN(_12896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21844_ (.A1(net21373),
    .A2(net21380),
    .ZN(_12897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21845_ (.A1(_12896_),
    .A2(_12897_),
    .ZN(_12898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21846_ (.A1(_12898_),
    .A2(net21379),
    .ZN(_12899_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21847_ (.A1(net20941),
    .A2(net20991),
    .A3(_12897_),
    .ZN(_12900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21848_ (.A1(_12899_),
    .A2(_12900_),
    .ZN(_12901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21849_ (.A1(_12895_),
    .A2(_12901_),
    .ZN(_12902_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21850_ (.A1(_12892_),
    .A2(_12902_),
    .A3(net21094),
    .ZN(_12903_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21851_ (.I(net21142),
    .ZN(_12904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21852_ (.A1(net21487),
    .A2(\text_in_r[27] ),
    .ZN(_12905_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21853_ (.A1(_12903_),
    .A2(_12904_),
    .A3(_12905_),
    .ZN(_12906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21854_ (.A1(_12881_),
    .A2(_12901_),
    .ZN(_12907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21855_ (.A1(_12895_),
    .A2(_12891_),
    .ZN(_12908_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21856_ (.A1(_12907_),
    .A2(_12908_),
    .A3(net21094),
    .ZN(_12909_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21857_ (.A1(net21094),
    .A2(\text_in_r[27] ),
    .Z(_12910_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21858_ (.A1(_12909_),
    .A2(net21142),
    .A3(_12910_),
    .ZN(_12911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21859_ (.A1(_12906_),
    .A2(_12911_),
    .ZN(_12912_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17374 (.I(_06257_),
    .Z(net17374));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17372 (.I(_06314_),
    .Z(net17372));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21862_ (.A1(_12863_),
    .A2(net19820),
    .ZN(_12915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21863_ (.A1(net21144),
    .A2(_12803_),
    .ZN(_12916_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21864_ (.A1(_12801_),
    .A2(_12804_),
    .A3(_12802_),
    .ZN(_12917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21865_ (.A1(_12917_),
    .A2(_12916_),
    .ZN(_15770_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21866_ (.A1(net19275),
    .A2(net19281),
    .ZN(_12918_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21867_ (.I(_12918_),
    .ZN(_12919_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21868_ (.A1(_12915_),
    .A2(net18310),
    .Z(_12920_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21869_ (.A1(net21378),
    .A2(net21263),
    .ZN(_12921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21870_ (.A1(_12921_),
    .A2(net20887),
    .ZN(_12922_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21871_ (.A1(net21378),
    .A2(net21263),
    .Z(_12923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21872_ (.A1(_12923_),
    .A2(net20888),
    .ZN(_12924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21873_ (.A1(_12922_),
    .A2(_12924_),
    .ZN(_12925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21874_ (.I(_12925_),
    .ZN(_12926_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21875_ (.A1(net21434),
    .A2(net21438),
    .Z(_12927_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21876_ (.I(\sa21_sub[4] ),
    .ZN(_12928_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21877_ (.A1(_12927_),
    .A2(net20990),
    .Z(_12929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21878_ (.A1(_12927_),
    .A2(net20990),
    .ZN(_12930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21879_ (.A1(_12929_),
    .A2(_12930_),
    .ZN(_12931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21880_ (.A1(_12926_),
    .A2(_12931_),
    .ZN(_12932_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21881_ (.A1(_12927_),
    .A2(net20990),
    .Z(_12933_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21882_ (.A1(_12927_),
    .A2(net20990),
    .ZN(_12934_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21883_ (.A1(_12933_),
    .A2(_12934_),
    .ZN(_12935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21884_ (.A1(_12935_),
    .A2(_12925_),
    .ZN(_12936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21885_ (.A1(_12932_),
    .A2(_12936_),
    .A3(net21093),
    .ZN(_12937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21886_ (.A1(net21487),
    .A2(\text_in_r[28] ),
    .ZN(_12938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21887_ (.A1(_12937_),
    .A2(_12938_),
    .ZN(_12939_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21888_ (.I(net21141),
    .ZN(_12940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21889_ (.A1(_12939_),
    .A2(_12940_),
    .ZN(_12941_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21890_ (.A1(_12937_),
    .A2(net21141),
    .A3(_12938_),
    .ZN(_12942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21891_ (.A1(_12941_),
    .A2(_12942_),
    .ZN(_12943_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17358 (.I(_10852_),
    .Z(net17358));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17377 (.I(_06204_),
    .Z(net17377));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21894_ (.A1(net19291),
    .A2(net19286),
    .ZN(_12946_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _21895_ (.I(_12912_),
    .ZN(_12947_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17385 (.I(_05540_),
    .Z(net17385));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21897_ (.A1(_12946_),
    .A2(net19267),
    .ZN(_12949_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21898_ (.I(_15785_[0]),
    .ZN(_12950_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21899_ (.A1(net20038),
    .A2(net19822),
    .A3(_12950_),
    .ZN(_12951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21900_ (.I(_12951_),
    .ZN(_12952_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21901_ (.A1(_12949_),
    .A2(_12952_),
    .Z(_12953_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21902_ (.A1(_12920_),
    .A2(net18858),
    .A3(_12953_),
    .ZN(_12954_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21903_ (.A1(\sa10_sub[4] ),
    .A2(\sa03_sr[4] ),
    .Z(_12955_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21904_ (.A1(\sa21_sub[5] ),
    .A2(\sa32_sub[5] ),
    .Z(_12956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21905_ (.A1(net21319),
    .A2(\sa32_sub[5] ),
    .ZN(_12957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21906_ (.A1(_12956_),
    .A2(_12957_),
    .ZN(_12958_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21907_ (.A1(\sa10_sub[5] ),
    .A2(_12958_),
    .Z(_12959_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21908_ (.A1(net20989),
    .A2(_12959_),
    .Z(_12960_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17356 (.I(_11329_),
    .Z(net17356));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21910_ (.I(net21140),
    .ZN(_12962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21911_ (.A1(net21487),
    .A2(\text_in_r[29] ),
    .ZN(_12963_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21912_ (.A1(_12960_),
    .A2(net21487),
    .B(_12962_),
    .C(_12963_),
    .ZN(_12964_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17384 (.I(_05558_),
    .Z(net17384));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21914_ (.A1(_12960_),
    .A2(net21093),
    .ZN(_12966_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21915_ (.A1(net21093),
    .A2(\text_in_r[29] ),
    .Z(_12967_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21916_ (.A1(_12966_),
    .A2(net21140),
    .A3(_12967_),
    .ZN(_12968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21917_ (.A1(_12964_),
    .A2(_12968_),
    .ZN(_12969_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17373 (.I(net17372),
    .Z(net17373));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19076 (.I(net19075),
    .Z(net19076));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21920_ (.A1(net19281),
    .A2(net18416),
    .Z(_12972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21921_ (.A1(_12972_),
    .A2(net19814),
    .ZN(_12973_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _21922_ (.I(_12943_),
    .ZN(_12974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21923_ (.A1(_12973_),
    .A2(_12974_),
    .ZN(_12975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21924_ (.A1(net19277),
    .A2(net19287),
    .ZN(_12976_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21925_ (.I(_12976_),
    .ZN(_12977_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17354 (.I(_11406_),
    .Z(net17354));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21927_ (.A1(_12977_),
    .A2(net19809),
    .Z(_12979_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21928_ (.A1(_12975_),
    .A2(_12979_),
    .ZN(_12980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21929_ (.A1(_12861_),
    .A2(_15778_[0]),
    .ZN(_12981_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21930_ (.A1(_12981_),
    .A2(net19277),
    .ZN(_12982_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21931_ (.A1(net18298),
    .A2(_12949_),
    .Z(_12983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21932_ (.A1(_12980_),
    .A2(_12983_),
    .ZN(_12984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21933_ (.A1(_12954_),
    .A2(net20264),
    .A3(_12984_),
    .ZN(_12985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21934_ (.A1(_12946_),
    .A2(net19809),
    .ZN(_12986_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21935_ (.A1(_12986_),
    .A2(_12974_),
    .Z(_12987_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21936_ (.I(_15776_[0]),
    .ZN(_12988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21937_ (.A1(net19281),
    .A2(_12988_),
    .ZN(_12989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21938_ (.A1(_12989_),
    .A2(_12947_),
    .Z(_12990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21939_ (.A1(net17550),
    .A2(net18871),
    .ZN(_12991_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17351 (.I(_11474_),
    .Z(net17351));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21941_ (.A1(_12987_),
    .A2(_12991_),
    .B(net20264),
    .ZN(_12993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21942_ (.A1(net19283),
    .A2(net19286),
    .ZN(_12994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21943_ (.A1(_12863_),
    .A2(net19820),
    .A3(net18848),
    .ZN(_12995_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21944_ (.I(_15772_[0]),
    .ZN(_12996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21945_ (.A1(net20038),
    .A2(_12996_),
    .A3(net19822),
    .ZN(_12997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21946_ (.A1(_12947_),
    .A2(_12997_),
    .ZN(_12998_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21947_ (.I(_12998_),
    .ZN(_12999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21948_ (.A1(net19287),
    .A2(_12950_),
    .ZN(_13000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21949_ (.A1(_12999_),
    .A2(net17902),
    .ZN(_13001_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17348 (.I(_11542_),
    .Z(net17348));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21951_ (.A1(_12995_),
    .A2(_13001_),
    .A3(net18855),
    .ZN(_13003_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21952_ (.A1(\sa10_sub[5] ),
    .A2(\sa03_sr[5] ),
    .ZN(_13004_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21953_ (.A1(\sa21_sub[6] ),
    .A2(\sa32_sub[6] ),
    .Z(_13005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21954_ (.A1(\sa21_sub[6] ),
    .A2(net21261),
    .ZN(_13006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21955_ (.A1(_13005_),
    .A2(_13006_),
    .ZN(_13007_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21956_ (.A1(net21376),
    .A2(_13007_),
    .Z(_13008_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21957_ (.A1(_13004_),
    .A2(_13008_),
    .Z(_13009_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17353 (.I(_11456_),
    .Z(net17353));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21959_ (.A1(net21489),
    .A2(\text_in_r[30] ),
    .Z(_13011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21960_ (.A1(_13009_),
    .A2(net21092),
    .B(_13011_),
    .ZN(_13012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21961_ (.A1(_13012_),
    .A2(\u0.tmp_w[30] ),
    .Z(_13013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21962_ (.A1(_13012_),
    .A2(\u0.tmp_w[30] ),
    .ZN(_13014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21963_ (.A1(_13013_),
    .A2(_13014_),
    .Z(_13015_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17349 (.I(_11503_),
    .Z(net17349));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17347 (.I(_11643_),
    .Z(net17347));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21966_ (.A1(_13003_),
    .A2(_12993_),
    .B(net20263),
    .ZN(_13018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21967_ (.A1(_12985_),
    .A2(_13018_),
    .ZN(_13019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21968_ (.A1(_12981_),
    .A2(net19809),
    .ZN(_13020_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21969_ (.I(_13020_),
    .ZN(_13021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21970_ (.A1(net19277),
    .A2(net19286),
    .ZN(_13022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21971_ (.A1(_13021_),
    .A2(net18846),
    .ZN(_13023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21972_ (.A1(net19299),
    .A2(net19286),
    .ZN(_13024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21973_ (.A1(net19287),
    .A2(net19296),
    .ZN(_13025_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17381 (.I(_06057_),
    .Z(net17381));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21975_ (.A1(net18845),
    .A2(_13025_),
    .A3(net19269),
    .ZN(_13027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21976_ (.A1(_13023_),
    .A2(net18864),
    .A3(_13027_),
    .ZN(_13028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21977_ (.A1(net17905),
    .A2(net19819),
    .Z(_13029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21978_ (.A1(net19297),
    .A2(net19293),
    .A3(net19296),
    .ZN(_13030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21979_ (.A1(_13029_),
    .A2(net18840),
    .ZN(_13031_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21980_ (.I(_15771_[0]),
    .ZN(_13032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21981_ (.A1(net19287),
    .A2(net18293),
    .ZN(_13033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21982_ (.I(_15779_[0]),
    .ZN(_13034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21983_ (.A1(net19282),
    .A2(net18291),
    .ZN(_13035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21984_ (.A1(_13033_),
    .A2(_13035_),
    .ZN(_13036_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17355 (.I(_11396_),
    .Z(net17355));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21986_ (.A1(_13036_),
    .A2(net19269),
    .ZN(_13038_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17390 (.I(net17389),
    .Z(net17390));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21988_ (.A1(_13031_),
    .A2(_13038_),
    .A3(net18300),
    .ZN(_13040_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21989_ (.A1(_12960_),
    .A2(net21487),
    .B(net21140),
    .C(_12963_),
    .ZN(_13041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21990_ (.A1(_12966_),
    .A2(_12962_),
    .A3(_12967_),
    .ZN(_13042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21991_ (.A1(_13041_),
    .A2(_13042_),
    .ZN(_13043_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17345 (.I(_11711_),
    .Z(net17345));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21993_ (.A1(_13028_),
    .A2(_13040_),
    .A3(net20260),
    .ZN(_13045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _21994_ (.A1(net20038),
    .A2(net19822),
    .A3(_13032_),
    .ZN(_13046_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21995_ (.I(_13046_),
    .ZN(_13047_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17340 (.I(_12138_),
    .Z(net17340));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21997_ (.A1(_13047_),
    .A2(net19810),
    .B(net18854),
    .ZN(_13049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21998_ (.A1(net19287),
    .A2(net18418),
    .ZN(_13050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21999_ (.A1(_12999_),
    .A2(net18290),
    .ZN(_13051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22000_ (.A1(net19291),
    .A2(_13034_),
    .Z(_13052_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17344 (.I(_11711_),
    .Z(net17344));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22002_ (.A1(net533),
    .A2(net19812),
    .ZN(_13054_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22003_ (.A1(_13049_),
    .A2(_13051_),
    .A3(_13054_),
    .ZN(_13055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22004_ (.A1(net19279),
    .A2(net18417),
    .ZN(_13056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22005_ (.A1(_13056_),
    .A2(net19809),
    .ZN(_13057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22006_ (.A1(net19297),
    .A2(net19293),
    .ZN(_13058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22007_ (.I(net18839),
    .ZN(_13059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22008_ (.A1(net19287),
    .A2(net18296),
    .ZN(_13060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22009_ (.A1(_12947_),
    .A2(_13060_),
    .ZN(_13061_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22010_ (.A1(net17897),
    .A2(_13059_),
    .B(net17547),
    .ZN(_13062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22011_ (.A1(_13062_),
    .A2(net18854),
    .ZN(_13063_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17339 (.I(_12164_),
    .Z(net17339));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22013_ (.A1(_13055_),
    .A2(_13063_),
    .A3(net20268),
    .ZN(_13065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22014_ (.A1(_13045_),
    .A2(_13065_),
    .A3(net20263),
    .ZN(_13066_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17335 (.I(_12233_),
    .Z(net17335));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22016_ (.A1(\sa03_sr[6] ),
    .A2(net21315),
    .Z(_13068_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22017_ (.A1(net21373),
    .A2(net21376),
    .Z(_13069_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _22018_ (.A1(net21259),
    .A2(_13068_),
    .A3(_13069_),
    .Z(_13070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22019_ (.I0(_13070_),
    .I1(\text_in_r[31] ),
    .S(net21489),
    .Z(_13071_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22020_ (.A1(_07739_),
    .A2(_13071_),
    .Z(_13072_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17401 (.I(_04199_),
    .Z(net17401));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22022_ (.A1(_13066_),
    .A2(_13019_),
    .A3(net20806),
    .ZN(_13074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22023_ (.A1(net19287),
    .A2(_12988_),
    .ZN(_13075_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22024_ (.A1(_13024_),
    .A2(net19289),
    .B(_13075_),
    .C(net19811),
    .ZN(_13076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22025_ (.A1(net19287),
    .A2(net18416),
    .ZN(_13077_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22026_ (.I(_13077_),
    .ZN(_13078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22027_ (.A1(_13078_),
    .A2(net19811),
    .Z(_13079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22028_ (.I(_13079_),
    .ZN(_13080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22029_ (.I(_13025_),
    .ZN(_13081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17346 (.I(_11644_),
    .Z(net17346));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22031_ (.A1(_13081_),
    .A2(_13047_),
    .B(net19269),
    .ZN(_13083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22032_ (.A1(_13076_),
    .A2(_13080_),
    .A3(_13083_),
    .ZN(_13084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22033_ (.A1(net19287),
    .A2(net18417),
    .ZN(_13085_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22034_ (.A1(_13085_),
    .A2(net19271),
    .B(net18854),
    .ZN(_13086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22035_ (.A1(net19271),
    .A2(_15792_[0]),
    .Z(_13087_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22036_ (.A1(_13086_),
    .A2(_13087_),
    .Z(_13088_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22037_ (.A1(_13084_),
    .A2(net18862),
    .B(net20268),
    .C(_13088_),
    .ZN(_13089_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22038_ (.I(_12975_),
    .ZN(_13090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22039_ (.A1(net19297),
    .A2(_12861_),
    .ZN(_13091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22040_ (.I(_13091_),
    .ZN(_13092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22041_ (.A1(_13092_),
    .A2(net19286),
    .ZN(_13093_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22042_ (.I(_15781_[0]),
    .ZN(_13094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22043_ (.A1(_12856_),
    .A2(_13094_),
    .ZN(_13095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22044_ (.A1(_13095_),
    .A2(_12947_),
    .ZN(_13096_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22045_ (.I(_13096_),
    .ZN(_13097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22046_ (.A1(_13093_),
    .A2(_13097_),
    .ZN(_13098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22047_ (.A1(_13090_),
    .A2(_13098_),
    .B(net20267),
    .ZN(_13099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22048_ (.A1(_12856_),
    .A2(_15779_[0]),
    .ZN(_13100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22049_ (.A1(_13100_),
    .A2(net19809),
    .ZN(_13101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22050_ (.I(_13101_),
    .ZN(_13102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22051_ (.A1(_13093_),
    .A2(net17545),
    .ZN(_13103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22052_ (.A1(_12972_),
    .A2(net19269),
    .ZN(_13104_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22053_ (.A1(_13103_),
    .A2(net18862),
    .A3(_13104_),
    .ZN(_13105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _22054_ (.I(_13015_),
    .ZN(_13106_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17330 (.I(_12274_),
    .Z(net17330));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22056_ (.A1(_13099_),
    .A2(_13105_),
    .B(net20036),
    .ZN(_13108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22057_ (.A1(_13089_),
    .A2(_13108_),
    .ZN(_13109_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17350 (.I(_11485_),
    .Z(net17350));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22059_ (.A1(_12998_),
    .A2(net18854),
    .Z(_13111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22060_ (.A1(net19287),
    .A2(net18415),
    .ZN(_13112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22061_ (.A1(net19279),
    .A2(net18414),
    .ZN(_13113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22062_ (.A1(_13112_),
    .A2(_13113_),
    .ZN(_13114_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17338 (.I(net17337),
    .Z(net17338));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22064_ (.A1(_13114_),
    .A2(net19813),
    .ZN(_13116_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22065_ (.A1(_13111_),
    .A2(_13116_),
    .B(net20258),
    .ZN(_13117_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _22066_ (.I(_13112_),
    .ZN(_13118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22067_ (.A1(_13118_),
    .A2(net19820),
    .B(net18854),
    .ZN(_13119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22068_ (.A1(_12983_),
    .A2(_13119_),
    .ZN(_13120_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22069_ (.A1(_13117_),
    .A2(_13120_),
    .B(net20263),
    .ZN(_13121_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17332 (.I(_12238_),
    .Z(net17332));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22071_ (.A1(net17550),
    .A2(_12974_),
    .ZN(_13123_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _22072_ (.I(_13033_),
    .ZN(_13124_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22073_ (.A1(_12972_),
    .A2(_13124_),
    .B(net19815),
    .ZN(_13125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22074_ (.A1(_13123_),
    .A2(_13125_),
    .B(net20264),
    .ZN(_13126_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22075_ (.A1(_13091_),
    .A2(net19814),
    .Z(_13127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22076_ (.A1(_13127_),
    .A2(_13085_),
    .ZN(_13128_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22077_ (.A1(net19283),
    .A2(net19296),
    .Z(_13129_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17472 (.I(_01757_),
    .Z(net17472));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22079_ (.A1(net18836),
    .A2(net532),
    .B(net19270),
    .ZN(_13131_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22080_ (.A1(_13128_),
    .A2(_13131_),
    .A3(net18305),
    .ZN(_13132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22081_ (.A1(_13126_),
    .A2(_13132_),
    .ZN(_13133_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22082_ (.A1(_13121_),
    .A2(_13133_),
    .B(net20807),
    .ZN(_13134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22083_ (.A1(_13109_),
    .A2(_13134_),
    .ZN(_13135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22084_ (.A1(_13074_),
    .A2(_13135_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22085_ (.A1(_13000_),
    .A2(_12947_),
    .ZN(_13136_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22086_ (.A1(_13136_),
    .A2(_12919_),
    .ZN(_13137_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22087_ (.A1(_13137_),
    .A2(_12974_),
    .ZN(_13138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22088_ (.A1(net19300),
    .A2(net19296),
    .ZN(_13139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22089_ (.A1(_13139_),
    .A2(net19281),
    .ZN(_13140_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17471 (.I(_01757_),
    .Z(net17471));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22091_ (.A1(_13140_),
    .A2(_12947_),
    .Z(_13142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22092_ (.A1(_13138_),
    .A2(_13142_),
    .ZN(_13143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22093_ (.A1(_13030_),
    .A2(net19269),
    .A3(_13056_),
    .ZN(_13144_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22094_ (.A1(net19280),
    .A2(net18415),
    .Z(_13145_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17317 (.I(_14025_),
    .Z(net17317));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22096_ (.A1(_13145_),
    .A2(net19810),
    .B(net18854),
    .ZN(_13147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22097_ (.A1(_13144_),
    .A2(_13147_),
    .ZN(_13148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22098_ (.A1(_13143_),
    .A2(net20258),
    .A3(_13148_),
    .ZN(_13149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22099_ (.A1(net18834),
    .A2(_12994_),
    .ZN(_13150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22100_ (.A1(_13150_),
    .A2(net19263),
    .ZN(_13151_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22101_ (.A1(net18847),
    .A2(_13085_),
    .A3(net19810),
    .ZN(_13152_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22102_ (.A1(_13151_),
    .A2(_13152_),
    .A3(net18300),
    .ZN(_13153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22103_ (.A1(_13025_),
    .A2(net19810),
    .A3(_13046_),
    .ZN(_13154_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22104_ (.A1(net18281),
    .A2(net17905),
    .A3(net19263),
    .ZN(_13155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22105_ (.A1(_13154_),
    .A2(_13155_),
    .ZN(_13156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22106_ (.A1(_13156_),
    .A2(net18865),
    .ZN(_13157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22107_ (.A1(_13153_),
    .A2(_13157_),
    .A3(net20270),
    .ZN(_13158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22108_ (.A1(_13149_),
    .A2(_13158_),
    .A3(net20035),
    .ZN(_13159_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17342 (.I(_12138_),
    .Z(net17342));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22110_ (.I(_13061_),
    .ZN(_13161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22111_ (.A1(_13161_),
    .A2(net17910),
    .ZN(_13162_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22112_ (.A1(_13076_),
    .A2(net18300),
    .A3(_13162_),
    .ZN(_13163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22113_ (.A1(_13058_),
    .A2(_12947_),
    .ZN(_13164_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22114_ (.A1(_13164_),
    .A2(_12918_),
    .Z(_13165_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _22115_ (.A1(_13118_),
    .A2(net19820),
    .B(_12974_),
    .ZN(_13166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22116_ (.A1(_13165_),
    .A2(_13166_),
    .B(net20258),
    .ZN(_13167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22117_ (.A1(_13163_),
    .A2(_13167_),
    .ZN(_13168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22118_ (.A1(_12999_),
    .A2(net18853),
    .ZN(_13169_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22119_ (.A1(_13025_),
    .A2(net17908),
    .A3(net19817),
    .ZN(_13170_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17341 (.I(net17340),
    .Z(net17341));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22121_ (.A1(_13169_),
    .A2(_13170_),
    .A3(net18858),
    .ZN(_13172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17352 (.I(_11469_),
    .Z(net17352));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _22123_ (.A1(net19808),
    .A2(net19279),
    .ZN(_13174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22124_ (.A1(net18845),
    .A2(net18833),
    .B(net18854),
    .ZN(_13175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22125_ (.A1(net18838),
    .A2(_13022_),
    .A3(net19814),
    .ZN(_13176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22126_ (.A1(_13175_),
    .A2(_13176_),
    .ZN(_13177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22127_ (.A1(_13172_),
    .A2(net20260),
    .A3(_13177_),
    .ZN(_13178_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22128_ (.A1(_13168_),
    .A2(_13178_),
    .A3(net20263),
    .ZN(_13179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22129_ (.A1(_13179_),
    .A2(_13159_),
    .B(net20807),
    .ZN(_13180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22130_ (.A1(_13024_),
    .A2(_13174_),
    .ZN(_13181_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22131_ (.A1(net19809),
    .A2(_13140_),
    .B(_13181_),
    .ZN(_13182_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22132_ (.A1(_12994_),
    .A2(_13050_),
    .A3(net19814),
    .ZN(_13183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22133_ (.I(_13183_),
    .ZN(_13184_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17343 (.I(_12055_),
    .Z(net17343));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22135_ (.A1(_13182_),
    .A2(_13184_),
    .B(net18859),
    .ZN(_13186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22136_ (.I(_12982_),
    .ZN(_13187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22137_ (.A1(_13187_),
    .A2(_13102_),
    .ZN(_13188_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22138_ (.I(_13188_),
    .ZN(_13189_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17329 (.I(_12274_),
    .Z(net17329));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22140_ (.I(_15795_[0]),
    .ZN(_13191_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22141_ (.A1(net19267),
    .A2(_13191_),
    .ZN(_13192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22142_ (.A1(_12974_),
    .A2(_13192_),
    .B(_13043_),
    .ZN(_13193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22143_ (.A1(_13189_),
    .A2(net18303),
    .B(_13193_),
    .ZN(_13194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22144_ (.A1(_13186_),
    .A2(_13194_),
    .ZN(_13195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22145_ (.A1(_13021_),
    .A2(net18839),
    .ZN(_13196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22146_ (.A1(_13196_),
    .A2(_12969_),
    .Z(_13197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22147_ (.A1(_12990_),
    .A2(_12976_),
    .ZN(_13198_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22148_ (.A1(_13198_),
    .A2(net18854),
    .Z(_13199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22149_ (.A1(_13197_),
    .A2(_13199_),
    .B(_13106_),
    .ZN(_13200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22150_ (.A1(_13195_),
    .A2(_13200_),
    .ZN(_13201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22151_ (.A1(_13201_),
    .A2(net20806),
    .ZN(_13202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22152_ (.A1(_13021_),
    .A2(net18290),
    .ZN(_13203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22153_ (.A1(_13203_),
    .A2(_13198_),
    .A3(net18300),
    .ZN(_13204_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22154_ (.A1(_13081_),
    .A2(_12972_),
    .B(net19811),
    .ZN(_13205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22155_ (.A1(_13085_),
    .A2(_13046_),
    .ZN(_13206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22156_ (.A1(_13206_),
    .A2(net19263),
    .ZN(_13207_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22157_ (.A1(_13205_),
    .A2(net18863),
    .A3(_13207_),
    .ZN(_13208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22158_ (.A1(_13204_),
    .A2(_13208_),
    .A3(net20260),
    .ZN(_13209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22159_ (.A1(_12951_),
    .A2(net19809),
    .Z(_13210_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22160_ (.I(_15773_[0]),
    .ZN(_13211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22161_ (.A1(net19287),
    .A2(net18276),
    .ZN(_13212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22162_ (.A1(_13210_),
    .A2(_13212_),
    .ZN(_13213_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22163_ (.A1(_13144_),
    .A2(_13213_),
    .A3(net18854),
    .ZN(_13214_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22164_ (.A1(net18298),
    .A2(_12986_),
    .B(_12974_),
    .C(_12998_),
    .ZN(_13215_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22165_ (.A1(_13214_),
    .A2(_13215_),
    .A3(net20267),
    .ZN(_13216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22166_ (.A1(_13209_),
    .A2(_13216_),
    .B(net20263),
    .ZN(_13217_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22167_ (.A1(_13202_),
    .A2(_13217_),
    .ZN(_13218_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22168_ (.A1(_13180_),
    .A2(_13218_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22169_ (.A1(_12994_),
    .A2(_13075_),
    .ZN(_13219_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22170_ (.A1(_13219_),
    .A2(net19270),
    .A3(_12918_),
    .ZN(_13220_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22171_ (.A1(_13220_),
    .A2(_13128_),
    .A3(net18305),
    .Z(_13221_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22172_ (.A1(net17907),
    .A2(net19817),
    .Z(_13222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22173_ (.A1(_13222_),
    .A2(net17902),
    .ZN(_13223_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22174_ (.A1(net18844),
    .A2(net18837),
    .A3(net19270),
    .ZN(_13224_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22175_ (.A1(_13223_),
    .A2(_13224_),
    .B(net18305),
    .ZN(_13225_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22176_ (.A1(_13221_),
    .A2(_13225_),
    .B(net20264),
    .ZN(_13226_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22177_ (.A1(net18871),
    .A2(net19815),
    .B(net18854),
    .ZN(_13227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22178_ (.A1(net18840),
    .A2(net19269),
    .A3(net17910),
    .ZN(_13228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22179_ (.A1(_13227_),
    .A2(_13228_),
    .B(net20267),
    .ZN(_13229_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _22180_ (.I(_13057_),
    .ZN(_13230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22181_ (.A1(_13230_),
    .A2(_12976_),
    .ZN(_13231_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22182_ (.I(_13231_),
    .ZN(_13232_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22183_ (.A1(net18849),
    .A2(_13077_),
    .A3(net19269),
    .Z(_13233_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22184_ (.A1(_13232_),
    .A2(_13233_),
    .B(net18862),
    .ZN(_13234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22185_ (.A1(_13229_),
    .A2(_13234_),
    .B(net20036),
    .ZN(_13235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22186_ (.A1(_13226_),
    .A2(_13235_),
    .ZN(_13236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22187_ (.A1(net19288),
    .A2(net18413),
    .ZN(_13237_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22188_ (.I(_13237_),
    .ZN(_13238_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22189_ (.A1(net18295),
    .A2(_13238_),
    .B(net18854),
    .ZN(_13239_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22190_ (.A1(net18851),
    .A2(_12947_),
    .A3(_13113_),
    .Z(_13240_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22191_ (.A1(_13239_),
    .A2(_13240_),
    .ZN(_13241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22192_ (.A1(net18847),
    .A2(net17891),
    .A3(net19810),
    .ZN(_13242_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22193_ (.A1(_13085_),
    .A2(net17906),
    .A3(net19264),
    .ZN(_13243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22194_ (.A1(_13242_),
    .A2(_13243_),
    .B(net18866),
    .ZN(_13244_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22195_ (.A1(_13241_),
    .A2(_13244_),
    .B(net20261),
    .ZN(_13245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22196_ (.A1(_13075_),
    .A2(net19269),
    .ZN(_13246_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22197_ (.A1(_13246_),
    .A2(_12919_),
    .Z(_13247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22198_ (.A1(_13247_),
    .A2(net18300),
    .A3(_13116_),
    .ZN(_13248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22199_ (.A1(net18280),
    .A2(_13237_),
    .ZN(_13249_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17306 (.I(_15175_),
    .Z(net17306));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22201_ (.A1(_13249_),
    .A2(net19810),
    .ZN(_13251_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22202_ (.A1(net18847),
    .A2(net17895),
    .A3(net19265),
    .ZN(_13252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22203_ (.A1(_13251_),
    .A2(_13252_),
    .A3(net18865),
    .ZN(_13253_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22204_ (.A1(_13248_),
    .A2(_13253_),
    .A3(net20271),
    .ZN(_13254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22205_ (.A1(_13245_),
    .A2(_13254_),
    .A3(net20035),
    .ZN(_13255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22206_ (.A1(_13236_),
    .A2(_13255_),
    .A3(net20807),
    .ZN(_13256_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22207_ (.A1(_13211_),
    .A2(_12988_),
    .Z(_13257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22208_ (.A1(net19281),
    .A2(_13257_),
    .ZN(_13258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22209_ (.A1(net18840),
    .A2(net19269),
    .A3(net17539),
    .ZN(_13259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22210_ (.A1(net17318),
    .A2(_13259_),
    .A3(net18859),
    .ZN(_13260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22211_ (.A1(_12999_),
    .A2(net17894),
    .ZN(_13261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22212_ (.A1(_13261_),
    .A2(_13049_),
    .B(_13106_),
    .ZN(_13262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22213_ (.A1(_13262_),
    .A2(_13260_),
    .B(net20268),
    .ZN(_13263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22214_ (.A1(_13093_),
    .A2(net17319),
    .ZN(_13264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22215_ (.A1(net18412),
    .A2(net19816),
    .B(net18854),
    .ZN(_13265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22216_ (.A1(_13264_),
    .A2(_13265_),
    .B(net20263),
    .ZN(_13266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22217_ (.A1(net18839),
    .A2(net18849),
    .ZN(_13267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22218_ (.A1(_13267_),
    .A2(net19269),
    .ZN(_13268_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22219_ (.A1(_13128_),
    .A2(net18864),
    .A3(_13268_),
    .ZN(_13269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22220_ (.A1(_13266_),
    .A2(_13269_),
    .ZN(_13270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22221_ (.A1(_13270_),
    .A2(_13263_),
    .B(net20806),
    .ZN(_13271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22222_ (.A1(_13127_),
    .A2(net17900),
    .Z(_13272_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22223_ (.A1(_13085_),
    .A2(_13035_),
    .A3(net19269),
    .Z(_13273_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22224_ (.A1(_13272_),
    .A2(_13273_),
    .B(net18864),
    .ZN(_13274_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22225_ (.A1(_13091_),
    .A2(_13022_),
    .A3(net19271),
    .Z(_13275_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22226_ (.A1(_13275_),
    .A2(net18854),
    .ZN(_13276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22227_ (.A1(net19820),
    .A2(net18277),
    .ZN(_13277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22228_ (.A1(_13276_),
    .A2(_13277_),
    .ZN(_13278_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22229_ (.A1(_13274_),
    .A2(_13278_),
    .A3(net20037),
    .ZN(_13279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22230_ (.A1(net19820),
    .A2(_15799_[0]),
    .ZN(_13280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22231_ (.A1(_13224_),
    .A2(_13280_),
    .B(net18303),
    .ZN(_13281_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _22232_ (.A1(net19820),
    .A2(_15790_[0]),
    .Z(_13282_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22233_ (.A1(_12915_),
    .A2(_13282_),
    .B(net18856),
    .ZN(_13283_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22234_ (.A1(_13281_),
    .A2(_13283_),
    .B(net20263),
    .ZN(_13284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22235_ (.A1(_13279_),
    .A2(_13284_),
    .A3(net20269),
    .ZN(_13285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22236_ (.A1(_13285_),
    .A2(_13271_),
    .ZN(_13286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22237_ (.A1(_13286_),
    .A2(_13256_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _22238_ (.A1(net19269),
    .A2(net18850),
    .A3(net18843),
    .A4(_13035_),
    .ZN(_13287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22239_ (.A1(_13085_),
    .A2(net19811),
    .Z(_13288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22240_ (.A1(_13288_),
    .A2(_13140_),
    .ZN(_13289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22241_ (.A1(_13287_),
    .A2(net18300),
    .A3(_13289_),
    .ZN(_13290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22242_ (.I(_13052_),
    .ZN(_13291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22243_ (.A1(_13029_),
    .A2(_13291_),
    .ZN(_13292_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22244_ (.A1(_13292_),
    .A2(_13027_),
    .A3(net18862),
    .ZN(_13293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22245_ (.A1(_13290_),
    .A2(_13293_),
    .ZN(_13294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22246_ (.A1(_13294_),
    .A2(net20258),
    .ZN(_13295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22247_ (.A1(_12947_),
    .A2(net19280),
    .Z(_13296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22248_ (.I(_13296_),
    .ZN(_13297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22249_ (.A1(_13024_),
    .A2(net18849),
    .ZN(_13298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22250_ (.A1(_13297_),
    .A2(_13298_),
    .Z(_13299_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22251_ (.A1(_13299_),
    .A2(net18300),
    .B(net20258),
    .ZN(_13300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22252_ (.A1(_13230_),
    .A2(net17891),
    .ZN(_13301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22253_ (.A1(_13138_),
    .A2(_13301_),
    .ZN(_13302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22254_ (.A1(_13300_),
    .A2(_13302_),
    .B(net20263),
    .ZN(_13303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22255_ (.A1(_13295_),
    .A2(_13303_),
    .ZN(_13304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22256_ (.A1(net18832),
    .A2(net18294),
    .B(net20270),
    .ZN(_13305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22257_ (.A1(_13174_),
    .A2(net18297),
    .Z(_13306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22258_ (.I(_13306_),
    .ZN(_13307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22259_ (.A1(net18843),
    .A2(_13035_),
    .ZN(_13308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22260_ (.A1(_13308_),
    .A2(net19810),
    .ZN(_13309_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22261_ (.A1(_13305_),
    .A2(_13307_),
    .A3(_13309_),
    .ZN(_13310_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22262_ (.A1(_13061_),
    .A2(net20270),
    .Z(_13311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22263_ (.A1(_13267_),
    .A2(net19810),
    .ZN(_13312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22264_ (.A1(_13311_),
    .A2(_13312_),
    .B(net18300),
    .ZN(_13313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22265_ (.A1(_13310_),
    .A2(_13313_),
    .B(net20035),
    .ZN(_13314_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22266_ (.A1(_13246_),
    .A2(_12952_),
    .Z(_13315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22267_ (.A1(_13315_),
    .A2(_13231_),
    .A3(net20258),
    .ZN(_13316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22268_ (.A1(net17901),
    .A2(net18845),
    .ZN(_13317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22269_ (.A1(_12999_),
    .A2(net18850),
    .ZN(_13318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22270_ (.A1(_13317_),
    .A2(_13318_),
    .A3(net20270),
    .ZN(_13319_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22271_ (.A1(_13316_),
    .A2(_13319_),
    .A3(net18300),
    .ZN(_13320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22272_ (.A1(_13320_),
    .A2(_13314_),
    .ZN(_13321_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22273_ (.I(_13072_),
    .ZN(_13322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22274_ (.A1(_13304_),
    .A2(_13321_),
    .A3(net20636),
    .ZN(_13323_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22275_ (.I(_13113_),
    .ZN(_13324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22276_ (.A1(net19263),
    .A2(_13324_),
    .B(net20270),
    .ZN(_13325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22277_ (.A1(_13325_),
    .A2(_13242_),
    .B(net18866),
    .ZN(_13326_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _22278_ (.I(_12986_),
    .ZN(_13327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22279_ (.A1(_13327_),
    .A2(net17906),
    .ZN(_13328_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22280_ (.A1(_13258_),
    .A2(net19269),
    .Z(_13329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22281_ (.A1(_13329_),
    .A2(net17904),
    .ZN(_13330_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22282_ (.A1(_13328_),
    .A2(_13330_),
    .A3(net20270),
    .ZN(_13331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22283_ (.A1(_13326_),
    .A2(_13331_),
    .B(net20035),
    .ZN(_13332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22284_ (.I(net17905),
    .ZN(_13333_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22285_ (.A1(_13333_),
    .A2(net19810),
    .Z(_13334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22286_ (.A1(_13334_),
    .A2(net20258),
    .B1(net19264),
    .B2(net18308),
    .ZN(_13335_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22287_ (.A1(net17890),
    .A2(net18284),
    .ZN(_13336_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22288_ (.A1(_13336_),
    .A2(_13306_),
    .B(net20266),
    .ZN(_13337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22289_ (.A1(_13335_),
    .A2(_13337_),
    .ZN(_13338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22290_ (.A1(_13338_),
    .A2(net18866),
    .ZN(_13339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22291_ (.A1(_13332_),
    .A2(_13339_),
    .B(_13322_),
    .ZN(_13340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22292_ (.A1(_13329_),
    .A2(net17891),
    .ZN(_13341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22293_ (.A1(net17318),
    .A2(_13341_),
    .B(net18865),
    .ZN(_13342_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22294_ (.I(_13239_),
    .ZN(_13343_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22295_ (.A1(_13342_),
    .A2(_13343_),
    .B(net20270),
    .ZN(_13344_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22296_ (.A1(_13083_),
    .A2(_13176_),
    .A3(net18300),
    .ZN(_13345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22297_ (.A1(_13029_),
    .A2(net669),
    .ZN(_13346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22298_ (.A1(_12946_),
    .A2(_13113_),
    .ZN(_13347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22299_ (.A1(_13347_),
    .A2(net19267),
    .ZN(_13348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22300_ (.A1(_13346_),
    .A2(_13348_),
    .A3(net18861),
    .ZN(_13349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22301_ (.A1(_13345_),
    .A2(_13349_),
    .A3(net20261),
    .ZN(_13350_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22302_ (.A1(_13344_),
    .A2(_13350_),
    .A3(net20035),
    .ZN(_13351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22303_ (.A1(_13340_),
    .A2(_13351_),
    .ZN(_13352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22304_ (.A1(_13323_),
    .A2(_13352_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22305_ (.A1(net17893),
    .A2(net19269),
    .A3(net18850),
    .ZN(_13353_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22306_ (.A1(_13353_),
    .A2(net18863),
    .A3(_13223_),
    .ZN(_13354_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22307_ (.A1(_13059_),
    .A2(_13047_),
    .B(net19266),
    .ZN(_13355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22308_ (.A1(_13076_),
    .A2(net18300),
    .A3(_13355_),
    .ZN(_13356_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22309_ (.A1(_13354_),
    .A2(_13356_),
    .A3(net20268),
    .ZN(_13357_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22310_ (.A1(_13174_),
    .A2(net18417),
    .Z(_13358_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22311_ (.A1(_13358_),
    .A2(_13324_),
    .ZN(_13359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22312_ (.A1(_13359_),
    .A2(_13166_),
    .B(net20267),
    .ZN(_13360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22313_ (.A1(net17541),
    .A2(net17896),
    .ZN(_13361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22314_ (.A1(_13098_),
    .A2(_13361_),
    .A3(net18300),
    .ZN(_13362_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22315_ (.A1(_13360_),
    .A2(_13362_),
    .B(net20036),
    .ZN(_13363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22316_ (.A1(_13357_),
    .A2(_13363_),
    .ZN(_13364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22317_ (.A1(_12918_),
    .A2(_13139_),
    .ZN(_13365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22318_ (.A1(net18868),
    .A2(net18290),
    .A3(net19269),
    .ZN(_13366_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22319_ (.A1(net19269),
    .A2(net18275),
    .B(_13366_),
    .C(net18864),
    .ZN(_13367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22320_ (.A1(_13276_),
    .A2(net17542),
    .ZN(_13368_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22321_ (.A1(_13367_),
    .A2(_13368_),
    .A3(net20269),
    .ZN(_13369_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22322_ (.I(_13164_),
    .ZN(_13370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22323_ (.A1(_13370_),
    .A2(_12994_),
    .ZN(_13371_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22324_ (.A1(_13371_),
    .A2(net17889),
    .A3(net18305),
    .ZN(_13372_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22325_ (.A1(net18307),
    .A2(net18300),
    .ZN(_13373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22326_ (.A1(_13373_),
    .A2(net17546),
    .B(net20269),
    .ZN(_13374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22327_ (.A1(_13372_),
    .A2(_13374_),
    .B(net20263),
    .ZN(_13375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22328_ (.A1(_13369_),
    .A2(_13375_),
    .ZN(_13376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22329_ (.A1(_13364_),
    .A2(_13376_),
    .A3(net20636),
    .ZN(_13377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22330_ (.A1(_12976_),
    .A2(net17899),
    .Z(_13378_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22331_ (.A1(_13378_),
    .A2(net19269),
    .Z(_13379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22332_ (.A1(_13199_),
    .A2(_13379_),
    .ZN(_13380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22333_ (.A1(net17901),
    .A2(net668),
    .ZN(_13381_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22334_ (.A1(net18833),
    .A2(net18854),
    .ZN(_13382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22335_ (.A1(_13381_),
    .A2(_13382_),
    .B(net20258),
    .ZN(_13383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22336_ (.A1(_13380_),
    .A2(_13383_),
    .ZN(_13384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22337_ (.A1(net19818),
    .A2(_13212_),
    .B(net18305),
    .ZN(_13385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22338_ (.A1(net18840),
    .A2(net19270),
    .ZN(_13386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22339_ (.A1(_13385_),
    .A2(_13386_),
    .B(net20264),
    .ZN(_13387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22340_ (.A1(_13222_),
    .A2(net18285),
    .ZN(_13388_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22341_ (.A1(_12983_),
    .A2(_13388_),
    .A3(_12974_),
    .ZN(_13389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22342_ (.A1(_13387_),
    .A2(_13389_),
    .ZN(_13390_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22343_ (.A1(_13384_),
    .A2(_13390_),
    .A3(net20037),
    .ZN(_13391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22344_ (.A1(_13129_),
    .A2(net19809),
    .ZN(_13392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22345_ (.A1(_13392_),
    .A2(net18854),
    .Z(_13393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22346_ (.A1(_13097_),
    .A2(net18869),
    .ZN(_13394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22347_ (.A1(net18309),
    .A2(net19818),
    .ZN(_13395_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22348_ (.A1(_13393_),
    .A2(_13394_),
    .A3(_13395_),
    .ZN(_13396_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22349_ (.I(_15783_[0]),
    .ZN(_13397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22350_ (.A1(_13397_),
    .A2(net19816),
    .B(net18854),
    .ZN(_13398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22351_ (.A1(net18285),
    .A2(net19272),
    .ZN(_13399_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22352_ (.A1(_13398_),
    .A2(_13399_),
    .B(net20264),
    .ZN(_13400_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22353_ (.A1(_13396_),
    .A2(_13400_),
    .B(net20037),
    .ZN(_13401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22354_ (.A1(_13097_),
    .A2(net18849),
    .ZN(_13402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22355_ (.A1(_13365_),
    .A2(net19815),
    .ZN(_13403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22356_ (.A1(_13402_),
    .A2(_13403_),
    .A3(net18854),
    .ZN(_13404_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22357_ (.A1(_13125_),
    .A2(net18306),
    .A3(_13027_),
    .ZN(_13405_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22358_ (.A1(_13404_),
    .A2(_13405_),
    .A3(net20268),
    .ZN(_13406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22359_ (.A1(_13401_),
    .A2(_13406_),
    .ZN(_13407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22360_ (.A1(_13391_),
    .A2(_13407_),
    .A3(net20806),
    .ZN(_13408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22361_ (.A1(_13377_),
    .A2(_13408_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22362_ (.A1(_13140_),
    .A2(net19269),
    .A3(_13291_),
    .Z(_13409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22363_ (.A1(_13327_),
    .A2(net18834),
    .ZN(_13410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22364_ (.A1(_13410_),
    .A2(net18854),
    .ZN(_13411_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22365_ (.A1(_13409_),
    .A2(_13411_),
    .ZN(_13412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22366_ (.A1(_12947_),
    .A2(net19278),
    .ZN(_13413_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22367_ (.A1(_13403_),
    .A2(_12974_),
    .A3(_13413_),
    .Z(_13414_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22368_ (.A1(_13412_),
    .A2(_13414_),
    .B(net20259),
    .ZN(_13415_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _22369_ (.A1(net18837),
    .A2(net19818),
    .A3(_13212_),
    .Z(_13416_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22370_ (.A1(_13416_),
    .A2(_13358_),
    .B(net18861),
    .ZN(_13417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22371_ (.A1(_13237_),
    .A2(net19819),
    .ZN(_13418_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22372_ (.A1(net17544),
    .A2(net17549),
    .B(_13418_),
    .C(net18300),
    .ZN(_13419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22373_ (.A1(_13417_),
    .A2(_13419_),
    .ZN(_13420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22374_ (.A1(_13420_),
    .A2(net20266),
    .ZN(_13421_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22375_ (.A1(_13415_),
    .A2(_13421_),
    .A3(net20263),
    .ZN(_13422_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22376_ (.A1(_13222_),
    .A2(_12974_),
    .ZN(_13423_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22377_ (.A1(_13423_),
    .A2(net18278),
    .B(net20258),
    .ZN(_13424_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22378_ (.I(_13029_),
    .ZN(_13425_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22379_ (.A1(_13348_),
    .A2(net18300),
    .A3(_13425_),
    .ZN(_13426_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22380_ (.A1(_13424_),
    .A2(_13426_),
    .B(net20263),
    .ZN(_13427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22381_ (.I(_13136_),
    .ZN(_13428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22382_ (.A1(_13428_),
    .A2(net17909),
    .ZN(_13429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22383_ (.A1(_12980_),
    .A2(_13429_),
    .ZN(_13430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22384_ (.A1(net17891),
    .A2(net19820),
    .Z(_13431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22385_ (.A1(_13093_),
    .A2(_13431_),
    .ZN(_13432_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22386_ (.A1(_13246_),
    .A2(_13257_),
    .Z(_13433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22387_ (.A1(_13432_),
    .A2(_13433_),
    .A3(net18858),
    .ZN(_13434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22388_ (.A1(_13430_),
    .A2(_13434_),
    .A3(net20259),
    .ZN(_13435_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22389_ (.A1(_13427_),
    .A2(_13435_),
    .B(net20807),
    .ZN(_13436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22390_ (.A1(_13422_),
    .A2(_13436_),
    .ZN(_13437_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22391_ (.I(_13329_),
    .ZN(_13438_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22392_ (.A1(net18312),
    .A2(net18299),
    .B(_13438_),
    .C(net18301),
    .ZN(_13439_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22393_ (.A1(_13166_),
    .A2(net17543),
    .B(net20264),
    .ZN(_13440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22394_ (.A1(_13439_),
    .A2(_13440_),
    .ZN(_13441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22395_ (.A1(net17888),
    .A2(net19821),
    .ZN(_13442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22396_ (.A1(net18292),
    .A2(net19268),
    .B(net18854),
    .ZN(_13443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22397_ (.A1(_13442_),
    .A2(_13443_),
    .B(net20257),
    .ZN(_13444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22398_ (.A1(_13230_),
    .A2(net17903),
    .ZN(_13445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22399_ (.A1(net17320),
    .A2(net18283),
    .ZN(_13446_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22400_ (.A1(_13445_),
    .A2(_13446_),
    .A3(net18854),
    .ZN(_13447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22401_ (.A1(_13444_),
    .A2(_13447_),
    .ZN(_13448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22402_ (.A1(_13441_),
    .A2(_13448_),
    .A3(net20263),
    .ZN(_13449_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22403_ (.A1(net19295),
    .A2(net19268),
    .B(net18854),
    .ZN(_13450_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22404_ (.A1(_13023_),
    .A2(_13450_),
    .B(net20264),
    .ZN(_13451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22405_ (.A1(_13431_),
    .A2(net18867),
    .ZN(_13452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22406_ (.A1(_12999_),
    .A2(net18870),
    .ZN(_13453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22407_ (.A1(_13452_),
    .A2(_13453_),
    .A3(net18855),
    .ZN(_13454_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22408_ (.A1(_13454_),
    .A2(_13451_),
    .B(net20263),
    .ZN(_13455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22409_ (.A1(_12983_),
    .A2(_13119_),
    .A3(net18274),
    .ZN(_13456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22410_ (.A1(net17888),
    .A2(net19821),
    .A3(net17903),
    .ZN(_13457_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22411_ (.A1(net17898),
    .A2(net19268),
    .B(net18302),
    .ZN(_13458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22412_ (.A1(_13457_),
    .A2(_13458_),
    .ZN(_13459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22413_ (.A1(_13456_),
    .A2(_13459_),
    .A3(net20265),
    .ZN(_13460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22414_ (.A1(_13455_),
    .A2(_13460_),
    .ZN(_13461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22415_ (.A1(_13449_),
    .A2(_13461_),
    .A3(net20806),
    .ZN(_13462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22416_ (.A1(_13437_),
    .A2(_13462_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22417_ (.A1(net17891),
    .A2(net17910),
    .A3(net19810),
    .ZN(_13463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22418_ (.A1(net18834),
    .A2(_13174_),
    .ZN(_13464_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22419_ (.A1(_13463_),
    .A2(_13104_),
    .A3(_13464_),
    .ZN(_13465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22420_ (.A1(_13465_),
    .A2(net18300),
    .ZN(_13466_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _22421_ (.A1(net19269),
    .A2(net18282),
    .A3(net18287),
    .A4(net18279),
    .ZN(_13467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22422_ (.I(_13392_),
    .ZN(_13468_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22423_ (.A1(_13086_),
    .A2(_13468_),
    .ZN(_13469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22424_ (.A1(_13467_),
    .A2(_13469_),
    .ZN(_13470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22425_ (.A1(_13466_),
    .A2(_13470_),
    .ZN(_13471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22426_ (.A1(_13471_),
    .A2(net20264),
    .ZN(_13472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22427_ (.A1(net18287),
    .A2(net18279),
    .Z(_13473_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22428_ (.A1(net17548),
    .A2(net19810),
    .ZN(_13474_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22429_ (.A1(_13473_),
    .A2(net19813),
    .B(net18861),
    .C(_13474_),
    .ZN(_13475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22430_ (.A1(_13365_),
    .A2(net19270),
    .ZN(_13476_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22431_ (.A1(_15788_[0]),
    .A2(_15797_[0]),
    .B(net19821),
    .ZN(_13477_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22432_ (.A1(_13476_),
    .A2(net18301),
    .A3(_13477_),
    .ZN(_13478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22433_ (.A1(_13475_),
    .A2(_13478_),
    .A3(net20258),
    .ZN(_13479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22434_ (.A1(_13472_),
    .A2(_13479_),
    .A3(_13106_),
    .ZN(_13480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22435_ (.A1(net19276),
    .A2(net19282),
    .B(net19820),
    .ZN(_13481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22436_ (.A1(_13481_),
    .A2(net18870),
    .ZN(_13482_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22437_ (.A1(net18288),
    .A2(net17887),
    .A3(net19821),
    .ZN(_13483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22438_ (.A1(_13482_),
    .A2(_13483_),
    .B(net18855),
    .ZN(_13484_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22439_ (.A1(net19267),
    .A2(net17905),
    .B(net18854),
    .ZN(_13485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22440_ (.A1(net18312),
    .A2(_13282_),
    .B(_13485_),
    .ZN(_13486_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22441_ (.A1(_13484_),
    .A2(_13486_),
    .B(net20257),
    .ZN(_13487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22442_ (.A1(net17886),
    .A2(net18844),
    .ZN(_13488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22443_ (.A1(net532),
    .A2(net19818),
    .B(net18305),
    .ZN(_13489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22444_ (.A1(_13488_),
    .A2(_13489_),
    .B(net20257),
    .ZN(_13490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22445_ (.A1(_13288_),
    .A2(net17539),
    .B(net18859),
    .ZN(_13491_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22446_ (.A1(_13093_),
    .A2(_12947_),
    .A3(net18842),
    .ZN(_13492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22447_ (.A1(_13491_),
    .A2(_13492_),
    .ZN(_13493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22448_ (.A1(_13490_),
    .A2(_13493_),
    .ZN(_13494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22449_ (.A1(_13487_),
    .A2(net20263),
    .A3(_13494_),
    .ZN(_13495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22450_ (.A1(_13480_),
    .A2(_13495_),
    .A3(net20636),
    .ZN(_13496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22451_ (.A1(_13164_),
    .A2(net18854),
    .Z(_13497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22452_ (.A1(_12995_),
    .A2(_13497_),
    .ZN(_13498_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22453_ (.A1(net18288),
    .A2(net19267),
    .Z(_13499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22454_ (.A1(_13348_),
    .A2(net18301),
    .A3(_13499_),
    .ZN(_13500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22455_ (.A1(_13498_),
    .A2(_13500_),
    .ZN(_13501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22456_ (.A1(_13501_),
    .A2(_13106_),
    .ZN(_13502_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22457_ (.A1(net17546),
    .A2(net18310),
    .B(net17890),
    .ZN(_13503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22458_ (.A1(_13503_),
    .A2(net18857),
    .ZN(_13504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22459_ (.A1(_13220_),
    .A2(net18304),
    .ZN(_13505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22460_ (.A1(_13504_),
    .A2(_13505_),
    .A3(net20263),
    .ZN(_13506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22461_ (.A1(_13502_),
    .A2(_13506_),
    .ZN(_13507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22462_ (.A1(_13507_),
    .A2(net20265),
    .ZN(_13508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22463_ (.A1(net19278),
    .A2(net19817),
    .ZN(_13509_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22464_ (.A1(_13298_),
    .A2(_12974_),
    .A3(_13509_),
    .Z(_13510_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22465_ (.A1(_13510_),
    .A2(net20263),
    .ZN(_13511_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22466_ (.A1(_13022_),
    .A2(net19270),
    .Z(_13512_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22467_ (.A1(_13512_),
    .A2(net17541),
    .B(net18842),
    .ZN(_13513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22468_ (.A1(_13513_),
    .A2(net18859),
    .ZN(_13514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22469_ (.A1(_13511_),
    .A2(_13514_),
    .ZN(_13515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22470_ (.A1(net18286),
    .A2(net19821),
    .B(net18302),
    .ZN(_13516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22471_ (.A1(_13428_),
    .A2(net18288),
    .ZN(_13517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22472_ (.A1(_13516_),
    .A2(_13517_),
    .ZN(_13518_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22473_ (.I(_15789_[0]),
    .ZN(_13519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22474_ (.A1(_13519_),
    .A2(net19268),
    .B(net18856),
    .ZN(_13520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22475_ (.A1(_13452_),
    .A2(_13520_),
    .ZN(_13521_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22476_ (.A1(_13518_),
    .A2(_13521_),
    .A3(net20263),
    .ZN(_13522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22477_ (.A1(_13515_),
    .A2(_13522_),
    .A3(net20257),
    .ZN(_13523_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22478_ (.A1(_13508_),
    .A2(net20806),
    .A3(_13523_),
    .ZN(_13524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22479_ (.A1(_13496_),
    .A2(_13524_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22480_ (.A1(net18832),
    .A2(net18835),
    .B(net18866),
    .ZN(_13525_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22481_ (.I(_13334_),
    .ZN(_13526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22482_ (.A1(_13525_),
    .A2(_13526_),
    .B(net20258),
    .ZN(_13527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22483_ (.A1(net17892),
    .A2(net19265),
    .ZN(_13528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22484_ (.A1(_13230_),
    .A2(net18840),
    .ZN(_13529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22485_ (.A1(_13528_),
    .A2(_13529_),
    .A3(net18865),
    .ZN(_13530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22486_ (.A1(_13527_),
    .A2(_13530_),
    .B(net20035),
    .ZN(_13531_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22487_ (.A1(net18841),
    .A2(net19816),
    .A3(net18868),
    .ZN(_13532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22488_ (.A1(_13276_),
    .A2(_13532_),
    .ZN(_13533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22489_ (.A1(net19818),
    .A2(net19286),
    .ZN(_13534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22490_ (.A1(_13371_),
    .A2(_13534_),
    .ZN(_13535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22491_ (.A1(_13535_),
    .A2(net18860),
    .ZN(_13536_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22492_ (.A1(_13533_),
    .A2(_13536_),
    .A3(net20260),
    .ZN(_13537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22493_ (.A1(_13531_),
    .A2(_13537_),
    .ZN(_13538_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22494_ (.A1(_13328_),
    .A2(net17220),
    .A3(net18865),
    .ZN(_13539_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22495_ (.A1(_13268_),
    .A2(net18300),
    .A3(_13463_),
    .ZN(_13540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22496_ (.A1(_13539_),
    .A2(_13540_),
    .A3(net20271),
    .ZN(_13541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22497_ (.A1(net17892),
    .A2(_13327_),
    .B(net18300),
    .ZN(_13542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22498_ (.A1(net18851),
    .A2(net18852),
    .ZN(_13543_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22499_ (.A1(_13543_),
    .A2(net17548),
    .B(net19266),
    .ZN(_13544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22500_ (.A1(_13542_),
    .A2(_13544_),
    .ZN(_13545_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22501_ (.A1(net17540),
    .A2(net18862),
    .ZN(_13546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22502_ (.A1(_13394_),
    .A2(_13546_),
    .B(net20267),
    .ZN(_13547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22503_ (.A1(_13545_),
    .A2(_13547_),
    .ZN(_13548_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22504_ (.A1(_13541_),
    .A2(_13548_),
    .A3(net20035),
    .ZN(_13549_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22505_ (.A1(_13538_),
    .A2(_13549_),
    .A3(net20808),
    .ZN(_13550_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22506_ (.A1(_13378_),
    .A2(_13327_),
    .Z(_13551_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22507_ (.A1(_12999_),
    .A2(_13291_),
    .Z(_13552_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22508_ (.A1(_13551_),
    .A2(_13552_),
    .B(net20262),
    .ZN(_13553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22509_ (.A1(net20270),
    .A2(net17899),
    .ZN(_13554_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22510_ (.A1(_13079_),
    .A2(_13554_),
    .ZN(_13555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22511_ (.A1(net18833),
    .A2(net19277),
    .ZN(_13556_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22512_ (.A1(_13555_),
    .A2(_13556_),
    .B(net18854),
    .ZN(_13557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22513_ (.A1(_13553_),
    .A2(_13557_),
    .ZN(_13558_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22514_ (.A1(_13543_),
    .A2(net18311),
    .B(net19813),
    .ZN(_13559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22515_ (.A1(_13559_),
    .A2(net20258),
    .A3(_13341_),
    .ZN(_13560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22516_ (.A1(net18415),
    .A2(net19810),
    .B(net20258),
    .ZN(_13561_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22517_ (.A1(_13561_),
    .A2(_13476_),
    .B(net18300),
    .ZN(_13562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22518_ (.A1(_13560_),
    .A2(_13562_),
    .ZN(_13563_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22519_ (.A1(_13558_),
    .A2(_13563_),
    .A3(net20036),
    .ZN(_13564_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22520_ (.A1(net18274),
    .A2(_13509_),
    .Z(_13565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22521_ (.A1(_13199_),
    .A2(_13565_),
    .ZN(_13566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22522_ (.A1(_13397_),
    .A2(net19272),
    .B(net18854),
    .ZN(_13567_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22523_ (.A1(_13080_),
    .A2(_13567_),
    .B(net20268),
    .ZN(_13568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22524_ (.A1(_13566_),
    .A2(_13568_),
    .ZN(_13569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22525_ (.A1(_13327_),
    .A2(net18869),
    .ZN(_13570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22526_ (.A1(net17319),
    .A2(net18289),
    .ZN(_13571_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22527_ (.A1(_13570_),
    .A2(_13571_),
    .A3(net18862),
    .ZN(_13572_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22528_ (.A1(_15797_[0]),
    .A2(net19268),
    .B(net18854),
    .ZN(_13573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22529_ (.A1(net17896),
    .A2(_13113_),
    .ZN(_13574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22530_ (.A1(_13574_),
    .A2(net19813),
    .ZN(_13575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22531_ (.A1(_13573_),
    .A2(_13575_),
    .B(net20258),
    .ZN(_13576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22532_ (.A1(_13572_),
    .A2(_13576_),
    .ZN(_13577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22533_ (.A1(_13569_),
    .A2(_13577_),
    .A3(net20263),
    .ZN(_13578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22534_ (.A1(_13564_),
    .A2(_13578_),
    .A3(net20636),
    .ZN(_13579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22535_ (.A1(_13550_),
    .A2(_13579_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22536_ (.I(\sa20_sr[7] ),
    .ZN(_13580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22537_ (.A1(_13580_),
    .A2(net21371),
    .ZN(_13581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22538_ (.A1(_10394_),
    .A2(net21361),
    .ZN(_13582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22539_ (.A1(_13581_),
    .A2(_13582_),
    .ZN(_13583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22540_ (.A1(_13583_),
    .A2(_10354_),
    .ZN(_13584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22541_ (.A1(_10394_),
    .A2(_13580_),
    .ZN(_13585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22542_ (.A1(net21370),
    .A2(net21361),
    .ZN(_13586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22543_ (.A1(_13585_),
    .A2(_13586_),
    .ZN(_13587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22544_ (.A1(_13587_),
    .A2(_10347_),
    .ZN(_13588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22545_ (.A1(_13584_),
    .A2(_13588_),
    .Z(_13589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22546_ (.A1(net21059),
    .A2(_10362_),
    .ZN(_13590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22547_ (.A1(net21478),
    .A2(_10366_),
    .ZN(_13591_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22548_ (.A1(_13591_),
    .A2(_13590_),
    .Z(_13592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22549_ (.A1(_13592_),
    .A2(_13589_),
    .ZN(_13593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22550_ (.A1(_13584_),
    .A2(_13588_),
    .ZN(_13594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22551_ (.A1(_13590_),
    .A2(_13591_),
    .ZN(_13595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22552_ (.A1(_13594_),
    .A2(_13595_),
    .ZN(_13596_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22553_ (.A1(_13596_),
    .A2(_13593_),
    .A3(_10378_),
    .ZN(_13597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22554_ (.A1(net21484),
    .A2(\text_in_r[113] ),
    .ZN(_13598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22555_ (.A1(_13597_),
    .A2(_13598_),
    .ZN(_13599_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22556_ (.I(net21229),
    .ZN(_13600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22557_ (.A1(_13599_),
    .A2(_13600_),
    .ZN(_13601_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22558_ (.A1(net20256),
    .A2(net21229),
    .A3(net20986),
    .ZN(_13602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22559_ (.A1(_13601_),
    .A2(_13602_),
    .ZN(_15807_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22560_ (.A1(net21097),
    .A2(net21312),
    .ZN(_13603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22561_ (.A1(net21062),
    .A2(net21414),
    .ZN(_13604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22562_ (.A1(_13603_),
    .A2(_13604_),
    .ZN(_13605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22563_ (.A1(_13605_),
    .A2(net21480),
    .ZN(_13606_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22564_ (.A1(_13603_),
    .A2(_13604_),
    .A3(net21101),
    .ZN(_13607_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22565_ (.A1(_13606_),
    .A2(_13607_),
    .A3(net20886),
    .ZN(_13608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22566_ (.A1(net21480),
    .A2(net21414),
    .ZN(_13609_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22567_ (.I(_13609_),
    .ZN(_13610_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22568_ (.A1(net21480),
    .A2(net21414),
    .ZN(_13611_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22569_ (.A1(_13610_),
    .A2(_13611_),
    .B(net21312),
    .ZN(_13612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22570_ (.A1(net21101),
    .A2(net21097),
    .ZN(_13613_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22571_ (.A1(_13613_),
    .A2(net21062),
    .A3(_13609_),
    .ZN(_13614_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22572_ (.A1(_13612_),
    .A2(_13614_),
    .A3(net20885),
    .ZN(_13615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22573_ (.A1(_13615_),
    .A2(_13608_),
    .B(net21493),
    .ZN(_13616_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22574_ (.I(\text_in_r[112] ),
    .ZN(_13617_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22575_ (.A1(_13617_),
    .A2(net21493),
    .Z(_13618_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22576_ (.A1(net20439),
    .A2(_13618_),
    .B(net21230),
    .ZN(_13619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22577_ (.A1(_13608_),
    .A2(_13615_),
    .ZN(_13620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22578_ (.A1(_13620_),
    .A2(net21064),
    .ZN(_13621_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22579_ (.I(net21230),
    .ZN(_13622_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22580_ (.I(_13618_),
    .ZN(_13623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22581_ (.A1(_13621_),
    .A2(_13622_),
    .A3(_13623_),
    .ZN(_13624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22582_ (.A1(_13624_),
    .A2(_13619_),
    .ZN(_15810_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22583_ (.A1(net21367),
    .A2(\sa30_sr[2] ),
    .ZN(_13625_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22584_ (.I(_13625_),
    .ZN(_13626_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22585_ (.A1(net21367),
    .A2(net21307),
    .ZN(_13627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22586_ (.A1(_13626_),
    .A2(_13627_),
    .B(net21476),
    .ZN(_13628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22587_ (.A1(_10417_),
    .A2(_10423_),
    .ZN(_13629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22588_ (.A1(_13629_),
    .A2(_10450_),
    .A3(_13625_),
    .ZN(_13630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22589_ (.A1(_13628_),
    .A2(_13630_),
    .ZN(_13631_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _22590_ (.A1(net21368),
    .A2(net21429),
    .ZN(_13632_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22591_ (.I(_13632_),
    .ZN(_13633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22592_ (.A1(_13633_),
    .A2(_13631_),
    .ZN(_13634_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22593_ (.A1(_13628_),
    .A2(_13630_),
    .A3(_13632_),
    .ZN(_13635_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22594_ (.A1(_13635_),
    .A2(net21066),
    .A3(_13634_),
    .ZN(_13636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22595_ (.A1(net21484),
    .A2(\text_in_r[114] ),
    .ZN(_13637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22596_ (.A1(_13636_),
    .A2(_13637_),
    .ZN(_13638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22597_ (.A1(_13638_),
    .A2(net21228),
    .ZN(_13639_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22598_ (.I(net21228),
    .ZN(_13640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22599_ (.A1(_13640_),
    .A2(net20438),
    .A3(_13637_),
    .ZN(_13641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22600_ (.A1(_13639_),
    .A2(_13641_),
    .ZN(_13642_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17461 (.I(_01963_),
    .Z(net17461));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22602_ (.A1(_13616_),
    .A2(_13618_),
    .B(_13622_),
    .ZN(_13643_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22603_ (.A1(_13621_),
    .A2(net21230),
    .A3(_13623_),
    .ZN(_13644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22604_ (.A1(_13644_),
    .A2(_13643_),
    .ZN(_15801_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22605_ (.A1(_13638_),
    .A2(_13640_),
    .ZN(_13645_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22606_ (.A1(_13636_),
    .A2(net21228),
    .A3(_13637_),
    .ZN(_13646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22607_ (.A1(_13645_),
    .A2(_13646_),
    .ZN(_13647_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17304 (.I(_15207_),
    .Z(net17304));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22609_ (.I(\sa30_sr[4] ),
    .ZN(_13648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22610_ (.A1(_10512_),
    .A2(_13648_),
    .ZN(_13649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22611_ (.A1(\sa20_sr[4] ),
    .A2(\sa30_sr[4] ),
    .ZN(_13650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22612_ (.A1(_13649_),
    .A2(_13650_),
    .ZN(_13651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22613_ (.A1(_10458_),
    .A2(net20987),
    .ZN(_13652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22614_ (.A1(net21365),
    .A2(net21362),
    .ZN(_13653_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22615_ (.A1(_13651_),
    .A2(net20937),
    .A3(net20983),
    .ZN(_13654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22616_ (.A1(_13652_),
    .A2(_13653_),
    .ZN(_13655_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22617_ (.A1(_13655_),
    .A2(net20984),
    .A3(net20938),
    .ZN(_13656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22618_ (.A1(_13654_),
    .A2(_13656_),
    .Z(_13657_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22619_ (.A1(net21473),
    .A2(_10473_),
    .Z(_13658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22620_ (.A1(_13657_),
    .A2(_13658_),
    .ZN(_13659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22621_ (.A1(_13654_),
    .A2(_13656_),
    .ZN(_13660_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22622_ (.A1(net21473),
    .A2(_10469_),
    .Z(_13661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22623_ (.A1(_13660_),
    .A2(_13661_),
    .ZN(_13662_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22624_ (.A1(_13659_),
    .A2(_13662_),
    .A3(net21065),
    .ZN(_13663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22625_ (.A1(net21489),
    .A2(\text_in_r[116] ),
    .ZN(_13664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22626_ (.A1(_13663_),
    .A2(_13664_),
    .ZN(_13665_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22627_ (.I(net21225),
    .ZN(_13666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22628_ (.A1(_13665_),
    .A2(_13666_),
    .ZN(_13667_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22629_ (.A1(_13663_),
    .A2(net21225),
    .A3(_13664_),
    .ZN(_13668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22630_ (.A1(_13667_),
    .A2(_13668_),
    .ZN(_13669_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17312 (.I(_14589_),
    .Z(net17312));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17308 (.I(net17307),
    .Z(net17308));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22633_ (.I(_15803_[0]),
    .ZN(_13672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22634_ (.A1(net19804),
    .A2(net18273),
    .Z(_13673_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _22635_ (.I(_15811_[0]),
    .ZN(_13674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22636_ (.A1(net19800),
    .A2(_13674_),
    .ZN(_13675_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22637_ (.I(_13675_),
    .ZN(_13676_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22638_ (.A1(_10417_),
    .A2(net20987),
    .ZN(_13677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22639_ (.A1(net21367),
    .A2(net21362),
    .ZN(_13678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22640_ (.A1(_13677_),
    .A2(_13678_),
    .ZN(_13679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22641_ (.A1(_10449_),
    .A2(_13679_),
    .ZN(_13680_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22642_ (.A1(net21367),
    .A2(net21362),
    .Z(_13681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22643_ (.A1(_13681_),
    .A2(_10462_),
    .ZN(_13682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22644_ (.A1(_13680_),
    .A2(_13682_),
    .ZN(_13683_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22645_ (.I(_13683_),
    .ZN(_13684_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22646_ (.A1(net504),
    .A2(net21055),
    .ZN(_13685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22647_ (.A1(net21413),
    .A2(net21424),
    .ZN(_13686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22648_ (.A1(_13685_),
    .A2(_13686_),
    .ZN(_13687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22649_ (.A1(_13687_),
    .A2(net21474),
    .ZN(_13688_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22650_ (.I(\sa00_sr[3] ),
    .ZN(_13689_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22651_ (.A1(_13685_),
    .A2(net20982),
    .A3(_13686_),
    .ZN(_13690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22652_ (.A1(_13688_),
    .A2(_13690_),
    .ZN(_13691_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22653_ (.I(_13691_),
    .ZN(_13692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22654_ (.A1(_13684_),
    .A2(_13692_),
    .ZN(_13693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22655_ (.A1(_13683_),
    .A2(_13691_),
    .ZN(_13694_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22656_ (.A1(_13693_),
    .A2(net21066),
    .A3(_13694_),
    .ZN(_13695_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22657_ (.A1(net21484),
    .A2(\text_in_r[115] ),
    .ZN(_13696_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22658_ (.A1(_13695_),
    .A2(_13696_),
    .ZN(_13697_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22659_ (.I(net21227),
    .ZN(_13698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22660_ (.A1(_13697_),
    .A2(_13698_),
    .ZN(_13699_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22661_ (.A1(_13695_),
    .A2(net21227),
    .A3(_13696_),
    .ZN(_13700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22662_ (.A1(_13699_),
    .A2(_13700_),
    .ZN(_13701_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17307 (.I(_15175_),
    .Z(net17307));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17300 (.I(_15266_),
    .Z(net17300));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22665_ (.A1(_13673_),
    .A2(_13676_),
    .B(net18816),
    .ZN(_13704_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22666_ (.I(_15804_[0]),
    .ZN(_13705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22667_ (.A1(net19799),
    .A2(_13705_),
    .ZN(_13706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22668_ (.A1(_13697_),
    .A2(net21227),
    .ZN(_13707_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22669_ (.A1(net20034),
    .A2(_13698_),
    .A3(_13696_),
    .ZN(_13708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22670_ (.A1(_13707_),
    .A2(_13708_),
    .ZN(_13709_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22671_ (.A1(net18806),
    .A2(_13706_),
    .Z(_13710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22672_ (.A1(net19260),
    .A2(net19807),
    .A3(net395),
    .ZN(_13711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22673_ (.A1(net17538),
    .A2(_13711_),
    .ZN(_13712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22674_ (.A1(_13704_),
    .A2(_13712_),
    .ZN(_13713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22675_ (.A1(net19798),
    .A2(net19806),
    .ZN(_13714_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17299 (.I(_15270_),
    .Z(net17299));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22677_ (.A1(net19244),
    .A2(net18806),
    .Z(_13716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22678_ (.A1(net21229),
    .A2(_13599_),
    .ZN(_13717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22679_ (.A1(_13597_),
    .A2(_13600_),
    .A3(_13598_),
    .ZN(_13718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22680_ (.A1(_13717_),
    .A2(_13718_),
    .ZN(_15802_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22681_ (.A1(net19243),
    .A2(net19801),
    .ZN(_13719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22682_ (.A1(_13716_),
    .A2(net18805),
    .ZN(_13720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22683_ (.A1(net19259),
    .A2(net19801),
    .ZN(_13721_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17311 (.I(_14813_),
    .Z(net17311));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17309 (.I(_15175_),
    .Z(net17309));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22686_ (.A1(net19807),
    .A2(net19802),
    .ZN(_13724_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22687_ (.A1(_13721_),
    .A2(net18825),
    .A3(_13724_),
    .ZN(_13725_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17296 (.I(net412),
    .Z(net17296));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22689_ (.A1(_13720_),
    .A2(_13725_),
    .A3(net19252),
    .ZN(_13727_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22690_ (.I(\sa00_sr[5] ),
    .ZN(_13728_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22691_ (.A1(_13728_),
    .A2(_10545_),
    .Z(_13729_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _22692_ (.A1(net21418),
    .A2(net21364),
    .ZN(_13730_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22693_ (.I(_13730_),
    .ZN(_13731_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22694_ (.A1(_13729_),
    .A2(_13731_),
    .Z(_13732_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22695_ (.A1(_13729_),
    .A2(_13731_),
    .ZN(_13733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22696_ (.A1(net21492),
    .A2(\text_in_r[117] ),
    .ZN(_13734_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _22697_ (.A1(_13732_),
    .A2(net21492),
    .A3(_13733_),
    .B(_13734_),
    .ZN(_13735_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22698_ (.A1(_13735_),
    .A2(net21224),
    .Z(_13736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22699_ (.A1(_13735_),
    .A2(net21224),
    .ZN(_13737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22700_ (.A1(_13736_),
    .A2(_13737_),
    .ZN(_13738_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _22701_ (.I(_13738_),
    .ZN(_13739_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17303 (.I(_15243_),
    .Z(net17303));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22703_ (.A1(net19252),
    .A2(_13713_),
    .B(_13727_),
    .C(net20028),
    .ZN(_13741_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22704_ (.I(\sa00_sr[6] ),
    .ZN(_13742_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22705_ (.A1(_13742_),
    .A2(_10582_),
    .Z(_13743_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _22706_ (.A1(net21417),
    .A2(\sa20_sr[5] ),
    .A3(_13743_),
    .Z(_13744_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22707_ (.A1(net21484),
    .A2(\text_in_r[118] ),
    .Z(_13745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22708_ (.A1(_13744_),
    .A2(net21095),
    .B(_13745_),
    .ZN(_13746_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22709_ (.A1(\u0.w[0][22] ),
    .A2(_13746_),
    .Z(_13747_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17301 (.I(_15246_),
    .Z(net17301));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17290 (.I(_00559_),
    .Z(net17290));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22712_ (.A1(net19802),
    .A2(_13705_),
    .ZN(_13750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22713_ (.A1(_13750_),
    .A2(net18813),
    .ZN(_13751_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22714_ (.A1(_13751_),
    .A2(net19251),
    .Z(_13752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22715_ (.A1(net19243),
    .A2(net19802),
    .ZN(_13753_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22716_ (.I(_13753_),
    .ZN(_13754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22717_ (.A1(_13754_),
    .A2(net18810),
    .ZN(_13755_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22718_ (.I(_13706_),
    .ZN(_13756_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17291 (.I(_00559_),
    .Z(net17291));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22720_ (.A1(_13756_),
    .A2(net18806),
    .ZN(_13758_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22721_ (.A1(_13752_),
    .A2(_13755_),
    .A3(_13758_),
    .Z(_13759_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22722_ (.A1(net19803),
    .A2(_13674_),
    .Z(_13760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22723_ (.A1(net19798),
    .A2(_13672_),
    .ZN(_13761_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _22724_ (.I(_13761_),
    .ZN(_13762_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17305 (.I(_15193_),
    .Z(net17305));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22726_ (.A1(_13760_),
    .A2(net17537),
    .B(net18809),
    .ZN(_13764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22727_ (.A1(_13706_),
    .A2(net18813),
    .ZN(_13765_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _22728_ (.I(_13765_),
    .ZN(_13766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22729_ (.A1(net19804),
    .A2(_15803_[0]),
    .ZN(_13767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22730_ (.A1(_13766_),
    .A2(_13767_),
    .ZN(_13768_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17292 (.I(_15388_),
    .Z(net17292));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22732_ (.A1(_13768_),
    .A2(_13764_),
    .B(net19257),
    .ZN(_13770_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17282 (.I(_01761_),
    .Z(net17282));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17288 (.I(_01283_),
    .Z(net17288));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22735_ (.A1(_13770_),
    .A2(_13759_),
    .B(net20252),
    .ZN(_13773_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22736_ (.A1(_13741_),
    .A2(_13773_),
    .A3(net20635),
    .ZN(_13774_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22737_ (.I(_13714_),
    .ZN(_13775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22738_ (.A1(_13775_),
    .A2(net19261),
    .ZN(_13776_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17284 (.I(_01745_),
    .Z(net17284));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17277 (.I(_01839_),
    .Z(net17277));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22741_ (.A1(net19801),
    .A2(net19803),
    .ZN(_13779_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22742_ (.A1(_13776_),
    .A2(net18826),
    .A3(net19241),
    .ZN(_13780_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _22743_ (.I(_15805_[0]),
    .ZN(_13781_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _22744_ (.A1(_13781_),
    .A2(net19802),
    .ZN(_13782_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22745_ (.A1(net18806),
    .A2(net408),
    .B(_13669_),
    .ZN(_13783_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22746_ (.A1(_13780_),
    .A2(net17881),
    .A3(net17535),
    .ZN(_13784_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _22747_ (.I(_15817_[0]),
    .ZN(_13785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22748_ (.A1(net19799),
    .A2(_13785_),
    .ZN(_13786_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22749_ (.A1(_13786_),
    .A2(net18813),
    .Z(_13787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22750_ (.A1(_13665_),
    .A2(net21225),
    .ZN(_13788_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22751_ (.A1(net20255),
    .A2(_13666_),
    .A3(_13664_),
    .ZN(_13789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22752_ (.A1(_13788_),
    .A2(_13789_),
    .ZN(_13790_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17315 (.I(_14469_),
    .Z(net17315));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22754_ (.A1(_13787_),
    .A2(net396),
    .B(net19233),
    .ZN(_13792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22755_ (.A1(net416),
    .A2(net19243),
    .ZN(_13793_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17283 (.I(_01755_),
    .Z(net17283));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22757_ (.A1(net18797),
    .A2(net18812),
    .Z(_13795_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _22758_ (.A1(net19261),
    .A2(net19803),
    .A3(net19801),
    .ZN(_13796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22759_ (.A1(_13795_),
    .A2(net411),
    .ZN(_13797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22760_ (.A1(_13792_),
    .A2(_13797_),
    .ZN(_13798_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22761_ (.A1(_13784_),
    .A2(net20249),
    .A3(_13798_),
    .ZN(_13799_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22762_ (.A1(net19805),
    .A2(net19798),
    .ZN(_13800_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22763_ (.A1(_13800_),
    .A2(net18813),
    .ZN(_13801_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22764_ (.A1(net18268),
    .A2(net19258),
    .ZN(_13802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22765_ (.I(_15808_[0]),
    .ZN(_13803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22766_ (.A1(net417),
    .A2(_13803_),
    .ZN(_13804_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22767_ (.A1(_13804_),
    .A2(net18813),
    .Z(_13805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22768_ (.A1(_13805_),
    .A2(net630),
    .ZN(_13806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22769_ (.A1(_13802_),
    .A2(_13806_),
    .B(net20249),
    .ZN(_13807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22770_ (.A1(net19801),
    .A2(net19799),
    .ZN(_13808_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22771_ (.A1(_13808_),
    .A2(net18806),
    .Z(_13809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22772_ (.A1(_13809_),
    .A2(_13796_),
    .ZN(_13810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22773_ (.A1(net19802),
    .A2(_13785_),
    .ZN(_13811_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22774_ (.A1(_13811_),
    .A2(net18813),
    .Z(_13812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22775_ (.A1(net17534),
    .A2(net17885),
    .ZN(_13813_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22776_ (.A1(_13810_),
    .A2(_13813_),
    .A3(net19258),
    .ZN(_13814_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22777_ (.A1(_13807_),
    .A2(_13814_),
    .B(net20634),
    .ZN(_13815_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _22778_ (.A1(net21470),
    .A2(\sa10_sr[6] ),
    .A3(net21363),
    .Z(_13816_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _22779_ (.A1(net21362),
    .A2(net21298),
    .A3(_13816_),
    .Z(_13817_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22780_ (.A1(net21493),
    .A2(\text_in_r[119] ),
    .Z(_13818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22781_ (.A1(_13817_),
    .A2(net21065),
    .B(_13818_),
    .ZN(_13819_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _22782_ (.A1(\u0.w[0][23] ),
    .A2(_13819_),
    .Z(_13820_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _22783_ (.I(_13820_),
    .ZN(_13821_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19063 (.I(_04769_),
    .Z(net19063));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22785_ (.A1(_13799_),
    .A2(_13815_),
    .B(_13821_),
    .ZN(_13823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22786_ (.A1(_13774_),
    .A2(_13823_),
    .ZN(_13824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22787_ (.A1(_13721_),
    .A2(net19800),
    .A3(net18806),
    .ZN(_13825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22788_ (.A1(net395),
    .A2(net18407),
    .ZN(_13826_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _22789_ (.A1(_13826_),
    .A2(net18813),
    .Z(_13827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22790_ (.A1(_13825_),
    .A2(_13827_),
    .Z(_13828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22791_ (.A1(_13724_),
    .A2(_13761_),
    .Z(_13829_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19267 (.I(_12947_),
    .Z(net19267));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _22793_ (.A1(_13829_),
    .A2(net18809),
    .Z(_13831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22794_ (.A1(net395),
    .A2(net18410),
    .ZN(_13832_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22795_ (.A1(_13832_),
    .A2(net18813),
    .Z(_13833_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22796_ (.A1(_13833_),
    .A2(net19233),
    .Z(_13834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22797_ (.A1(_13828_),
    .A2(_13831_),
    .A3(_13834_),
    .ZN(_13835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22798_ (.A1(net529),
    .A2(net19802),
    .ZN(_13836_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _22799_ (.I(_13836_),
    .ZN(_13837_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22800_ (.A1(net18806),
    .A2(_13837_),
    .B(net19233),
    .ZN(_13838_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19332 (.I(net19331),
    .Z(net19332));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22802_ (.A1(net18825),
    .A2(_15824_[0]),
    .ZN(_13840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22803_ (.A1(_13838_),
    .A2(_13840_),
    .B(net20029),
    .ZN(_13841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22804_ (.A1(_13835_),
    .A2(_13841_),
    .ZN(_13842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22805_ (.A1(net19259),
    .A2(net417),
    .ZN(_13843_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _22806_ (.I(_13843_),
    .ZN(_13844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22807_ (.A1(net19801),
    .A2(_13844_),
    .ZN(_13845_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _22808_ (.I(_15813_[0]),
    .ZN(_13846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22809_ (.A1(_13846_),
    .A2(net19802),
    .ZN(_13847_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22810_ (.A1(net18813),
    .A2(_13847_),
    .Z(_13848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22811_ (.A1(_13845_),
    .A2(_13848_),
    .ZN(_13849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22812_ (.A1(_13849_),
    .A2(net17535),
    .ZN(_13850_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22813_ (.A1(net19802),
    .A2(_15811_[0]),
    .ZN(_13851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22814_ (.A1(_13851_),
    .A2(net18806),
    .ZN(_13852_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22815_ (.I(_13852_),
    .ZN(_13853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22816_ (.A1(net530),
    .A2(_13853_),
    .ZN(_13854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22817_ (.A1(_13782_),
    .A2(net18813),
    .ZN(_13855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22818_ (.A1(_13855_),
    .A2(_13669_),
    .ZN(_13856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22819_ (.I(_13856_),
    .ZN(_13857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22820_ (.A1(_13854_),
    .A2(_13857_),
    .ZN(_13858_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22821_ (.A1(_13850_),
    .A2(_13858_),
    .A3(_13739_),
    .ZN(_13859_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22822_ (.A1(_13842_),
    .A2(_13859_),
    .A3(net20634),
    .ZN(_13860_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _22823_ (.A1(net395),
    .A2(_13846_),
    .ZN(_13861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22824_ (.A1(_13861_),
    .A2(net18806),
    .ZN(_13862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22825_ (.A1(_13862_),
    .A2(net19256),
    .Z(_13863_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22826_ (.A1(_13863_),
    .A2(net17536),
    .A3(net17875),
    .ZN(_13864_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17266 (.I(_02652_),
    .Z(net17266));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22828_ (.A1(_13827_),
    .A2(net19233),
    .Z(_13866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22829_ (.A1(_13780_),
    .A2(_13866_),
    .ZN(_13867_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19306 (.I(net647),
    .Z(net19306));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22831_ (.A1(_13864_),
    .A2(_13867_),
    .A3(net20249),
    .ZN(_13869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22832_ (.A1(_13843_),
    .A2(net18806),
    .ZN(_13870_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22833_ (.I(_13870_),
    .ZN(_13871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22834_ (.A1(_13871_),
    .A2(net18260),
    .ZN(_13872_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17270 (.I(_02066_),
    .Z(net17270));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17264 (.I(_02843_),
    .Z(net17264));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22837_ (.A1(net18798),
    .A2(_13760_),
    .B(net18825),
    .ZN(_13875_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22838_ (.A1(_13872_),
    .A2(net19237),
    .A3(_13875_),
    .ZN(_13876_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22839_ (.A1(_13805_),
    .A2(net19233),
    .ZN(_13877_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22840_ (.A1(_13673_),
    .A2(net17879),
    .B(net18808),
    .ZN(_13878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22841_ (.A1(_13877_),
    .A2(_13878_),
    .B(net20252),
    .ZN(_13879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22842_ (.A1(_13876_),
    .A2(_13879_),
    .ZN(_13880_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _22843_ (.I(net20634),
    .ZN(_13881_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17262 (.I(_02910_),
    .Z(net17262));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22845_ (.A1(_13869_),
    .A2(_13880_),
    .A3(_13881_),
    .ZN(_13883_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22846_ (.A1(_13860_),
    .A2(_13883_),
    .A3(_13821_),
    .ZN(_13884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22847_ (.A1(_13824_),
    .A2(_13884_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22848_ (.A1(net19261),
    .A2(net19801),
    .B(net19241),
    .C(net18825),
    .ZN(_13885_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17261 (.I(_03154_),
    .Z(net17261));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22850_ (.A1(net18260),
    .A2(net18806),
    .Z(_13887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22851_ (.A1(_13887_),
    .A2(net19231),
    .ZN(_13888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22852_ (.A1(_13885_),
    .A2(net19233),
    .A3(_13888_),
    .ZN(_13889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22853_ (.A1(_13829_),
    .A2(net18809),
    .ZN(_13890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22854_ (.A1(_13766_),
    .A2(net18264),
    .ZN(_13891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22855_ (.A1(_13890_),
    .A2(_13891_),
    .ZN(_13892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22856_ (.A1(_13892_),
    .A2(net19254),
    .ZN(_13893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22857_ (.A1(_13889_),
    .A2(_13893_),
    .A3(net20249),
    .ZN(_13894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22858_ (.A1(_13793_),
    .A2(_13808_),
    .ZN(_13895_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17285 (.I(_01721_),
    .Z(net17285));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22860_ (.A1(net18256),
    .A2(net18812),
    .ZN(_13897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22861_ (.A1(_13812_),
    .A2(net18797),
    .ZN(_13898_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17259 (.I(_03170_),
    .Z(net17259));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22863_ (.A1(_13897_),
    .A2(_13898_),
    .A3(net19258),
    .ZN(_13900_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19305 (.I(net19303),
    .Z(net19305));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19177 (.I(_15976_[0]),
    .Z(net19177));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22866_ (.A1(net18411),
    .A2(net19799),
    .ZN(_13903_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22867_ (.A1(_13711_),
    .A2(net18830),
    .A3(net18255),
    .ZN(_13904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22868_ (.A1(net19798),
    .A2(net18408),
    .ZN(_13905_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22869_ (.I(net18253),
    .ZN(_13906_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19282 (.I(net19281),
    .Z(net19282));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22871_ (.A1(_13906_),
    .A2(net18812),
    .B(net19258),
    .ZN(_13908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22872_ (.A1(_13904_),
    .A2(_13908_),
    .ZN(_13909_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22873_ (.A1(_13900_),
    .A2(net20033),
    .A3(_13909_),
    .ZN(_13910_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22874_ (.A1(_13894_),
    .A2(_13910_),
    .A3(_13881_),
    .ZN(_13911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22875_ (.A1(_13766_),
    .A2(net19241),
    .ZN(_13912_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22876_ (.A1(_13804_),
    .A2(net18806),
    .Z(_13913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22877_ (.A1(_13913_),
    .A2(_13724_),
    .ZN(_13914_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22878_ (.A1(_13912_),
    .A2(_13914_),
    .A3(net19254),
    .ZN(_13915_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22879_ (.A1(net18813),
    .A2(net395),
    .Z(_13916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22880_ (.A1(_13916_),
    .A2(net18803),
    .B(net19250),
    .ZN(_13917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22881_ (.A1(_13871_),
    .A2(net18805),
    .ZN(_13918_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22882_ (.A1(_13917_),
    .A2(_13918_),
    .ZN(_13919_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22883_ (.A1(_13915_),
    .A2(_13919_),
    .A3(net20032),
    .ZN(_13920_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22884_ (.A1(_13827_),
    .A2(net18796),
    .Z(_13921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22885_ (.A1(net19260),
    .A2(net395),
    .ZN(_13922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22886_ (.A1(_13922_),
    .A2(net18830),
    .B(net19233),
    .ZN(_13923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22887_ (.A1(_13921_),
    .A2(_13923_),
    .B(net20032),
    .ZN(_13924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22888_ (.A1(_13787_),
    .A2(net17883),
    .ZN(_13925_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22889_ (.A1(_13925_),
    .A2(net19240),
    .Z(_13926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22890_ (.A1(_13926_),
    .A2(_13828_),
    .ZN(_13927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22891_ (.A1(_13924_),
    .A2(_13927_),
    .ZN(_13928_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22892_ (.A1(_13920_),
    .A2(_13928_),
    .A3(net20635),
    .ZN(_13929_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22893_ (.A1(_13911_),
    .A2(_13929_),
    .A3(_13821_),
    .ZN(_13930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22894_ (.A1(net18270),
    .A2(net630),
    .A3(net18831),
    .ZN(_13931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22895_ (.A1(_13809_),
    .A2(_13767_),
    .ZN(_13932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22896_ (.A1(_13931_),
    .A2(net20031),
    .A3(_13932_),
    .ZN(_13933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22897_ (.A1(_13716_),
    .A2(net18792),
    .ZN(_13934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22898_ (.A1(_13805_),
    .A2(net18800),
    .ZN(_13935_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19513 (.I(net19512),
    .Z(net19513));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22900_ (.A1(_13934_),
    .A2(_13935_),
    .A3(net20249),
    .ZN(_13937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22901_ (.A1(_13933_),
    .A2(_13937_),
    .B(net19239),
    .ZN(_13938_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22902_ (.A1(_13739_),
    .A2(_15827_[0]),
    .A3(net18812),
    .Z(_13939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22903_ (.A1(net18270),
    .A2(_13853_),
    .ZN(_13940_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22904_ (.A1(_13939_),
    .A2(net19238),
    .A3(_13940_),
    .Z(_13941_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22905_ (.A1(_13938_),
    .A2(_13941_),
    .B(net20635),
    .ZN(_13942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22906_ (.A1(net18270),
    .A2(net18268),
    .ZN(_13943_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22907_ (.A1(_13765_),
    .A2(net19233),
    .Z(_13944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22908_ (.A1(_13943_),
    .A2(_13944_),
    .B(_13739_),
    .ZN(_13945_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22909_ (.A1(_13786_),
    .A2(net18806),
    .Z(_13946_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22910_ (.A1(net19803),
    .A2(net18269),
    .ZN(_13947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22911_ (.A1(_13946_),
    .A2(net17871),
    .B(net19238),
    .ZN(_13948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22912_ (.A1(_13948_),
    .A2(_13904_),
    .ZN(_13949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22913_ (.A1(_13945_),
    .A2(_13949_),
    .B(net20635),
    .ZN(_13950_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22914_ (.A1(_13724_),
    .A2(net18813),
    .Z(_13951_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22915_ (.A1(_13951_),
    .A2(net19250),
    .Z(_13952_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22916_ (.A1(net18828),
    .A2(_13837_),
    .ZN(_13953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22917_ (.A1(net17879),
    .A2(net18808),
    .ZN(_13954_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22918_ (.A1(_13953_),
    .A2(_13954_),
    .Z(_13955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22919_ (.A1(net17537),
    .A2(net18825),
    .ZN(_13956_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22920_ (.A1(_13952_),
    .A2(_13955_),
    .A3(_13956_),
    .ZN(_13957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22921_ (.A1(_13716_),
    .A2(_13767_),
    .ZN(_13958_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20459 (.I(_09742_),
    .Z(net20459));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22923_ (.A1(_13958_),
    .A2(_13935_),
    .A3(net19240),
    .ZN(_13960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22924_ (.A1(_13957_),
    .A2(net20032),
    .A3(_13960_),
    .ZN(_13961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22925_ (.A1(_13950_),
    .A2(_13961_),
    .B(_13821_),
    .ZN(_13962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22926_ (.A1(_13942_),
    .A2(_13962_),
    .ZN(_13963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22927_ (.A1(_13930_),
    .A2(_13963_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22928_ (.A1(_13808_),
    .A2(_13847_),
    .A3(net18806),
    .ZN(_13964_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22929_ (.A1(net17884),
    .A2(net18262),
    .A3(net18820),
    .ZN(_13965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22930_ (.A1(_13964_),
    .A2(_13965_),
    .ZN(_13966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22931_ (.A1(_13966_),
    .A2(net19235),
    .ZN(_13967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22932_ (.A1(net636),
    .A2(net19799),
    .ZN(_13968_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22933_ (.A1(net18799),
    .A2(net18814),
    .A3(_13968_),
    .ZN(_13969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22934_ (.A1(net395),
    .A2(net18406),
    .ZN(_13970_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22935_ (.A1(net19244),
    .A2(_13970_),
    .A3(net18806),
    .ZN(_13971_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22936_ (.A1(_13969_),
    .A2(net19249),
    .A3(_13971_),
    .ZN(_13972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22937_ (.A1(_13967_),
    .A2(_13972_),
    .ZN(_13973_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22938_ (.A1(_13973_),
    .A2(net20025),
    .B(net20634),
    .ZN(_13974_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22939_ (.A1(_13793_),
    .A2(net18813),
    .Z(_13975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22940_ (.A1(net395),
    .A2(net18266),
    .ZN(_13976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22941_ (.A1(_13975_),
    .A2(_13976_),
    .ZN(_13977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22942_ (.A1(_13977_),
    .A2(_13866_),
    .A3(net17532),
    .ZN(_13978_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _22943_ (.A1(net19247),
    .A2(net525),
    .A3(net18827),
    .Z(_13979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22944_ (.A1(_13970_),
    .A2(net18806),
    .ZN(_13980_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22945_ (.I(_13980_),
    .ZN(_13981_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22946_ (.A1(_13979_),
    .A2(_13981_),
    .B(_13863_),
    .ZN(_13982_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22947_ (.A1(_13978_),
    .A2(_13982_),
    .A3(net20249),
    .ZN(_13983_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22948_ (.A1(_13974_),
    .A2(_13983_),
    .B(_13821_),
    .ZN(_13984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22949_ (.A1(_13872_),
    .A2(net19237),
    .ZN(_13985_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22950_ (.A1(_13979_),
    .A2(_13793_),
    .Z(_13986_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22951_ (.A1(_13985_),
    .A2(_13986_),
    .ZN(_13987_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22952_ (.A1(net18804),
    .A2(net18793),
    .A3(net18825),
    .ZN(_13988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22953_ (.A1(_13970_),
    .A2(_13905_),
    .ZN(_13989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22954_ (.A1(_13989_),
    .A2(net18812),
    .ZN(_13990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22955_ (.A1(_13988_),
    .A2(_13990_),
    .B(net19237),
    .ZN(_13991_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22956_ (.A1(_13987_),
    .A2(_13991_),
    .B(net20249),
    .ZN(_13992_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22957_ (.A1(_13753_),
    .A2(net18806),
    .A3(_13903_),
    .ZN(_13993_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22958_ (.I(_13993_),
    .ZN(_13994_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22959_ (.A1(net19244),
    .A2(net18263),
    .A3(net18822),
    .Z(_13995_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22960_ (.A1(_13994_),
    .A2(_13995_),
    .B(net19253),
    .ZN(_13996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22961_ (.A1(_13711_),
    .A2(net18826),
    .A3(net17877),
    .ZN(_13997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22962_ (.A1(net631),
    .A2(net18811),
    .ZN(_13998_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22963_ (.A1(_13997_),
    .A2(net19237),
    .A3(_13998_),
    .ZN(_13999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22964_ (.A1(_13996_),
    .A2(_13999_),
    .A3(net20032),
    .ZN(_14000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22965_ (.A1(_13992_),
    .A2(net20635),
    .A3(_14000_),
    .ZN(_14001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22966_ (.A1(_13984_),
    .A2(_14001_),
    .ZN(_14002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22967_ (.A1(net18260),
    .A2(net18817),
    .ZN(_14003_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _22968_ (.A1(net18257),
    .A2(_13673_),
    .B1(_13676_),
    .B2(_14003_),
    .ZN(_14004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22969_ (.A1(_14004_),
    .A2(net19252),
    .ZN(_14005_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22970_ (.A1(_13719_),
    .A2(net18817),
    .Z(_14006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22971_ (.A1(_14006_),
    .A2(net18793),
    .ZN(_14007_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22972_ (.A1(net18825),
    .A2(_15827_[0]),
    .Z(_14008_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22973_ (.A1(_14007_),
    .A2(net19236),
    .A3(_14008_),
    .ZN(_14009_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22974_ (.A1(_14005_),
    .A2(net20254),
    .A3(_14009_),
    .ZN(_14010_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22975_ (.I(_13751_),
    .ZN(_14011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22976_ (.A1(_13845_),
    .A2(_14011_),
    .ZN(_14012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22977_ (.A1(_15824_[0]),
    .A2(net18809),
    .B(net19255),
    .ZN(_14013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22978_ (.A1(_14012_),
    .A2(_14013_),
    .B(net20252),
    .ZN(_14014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22979_ (.A1(_13922_),
    .A2(net19245),
    .ZN(_14015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _22980_ (.A1(_14015_),
    .A2(net18829),
    .ZN(_14016_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22981_ (.A1(_13872_),
    .A2(_14016_),
    .A3(net19254),
    .ZN(_14017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22982_ (.A1(_14014_),
    .A2(_14017_),
    .B(net20635),
    .ZN(_14018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22983_ (.A1(_14010_),
    .A2(_14018_),
    .ZN(_14019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22984_ (.A1(_13753_),
    .A2(_13779_),
    .ZN(_14020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22985_ (.I(_13782_),
    .ZN(_14021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22986_ (.A1(_14021_),
    .A2(net18253),
    .ZN(_14022_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22987_ (.A1(_14020_),
    .A2(_14022_),
    .B(net18825),
    .ZN(_14023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22988_ (.A1(_14023_),
    .A2(net19254),
    .A3(_13940_),
    .ZN(_14024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22989_ (.A1(_13762_),
    .A2(net18806),
    .ZN(_14025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22990_ (.A1(_14025_),
    .A2(net19233),
    .Z(_14026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22991_ (.A1(_13766_),
    .A2(_13976_),
    .ZN(_14027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22992_ (.A1(_14027_),
    .A2(_14026_),
    .B(net20252),
    .ZN(_14028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22993_ (.A1(_14028_),
    .A2(_14024_),
    .ZN(_14029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22994_ (.A1(net18809),
    .A2(_15831_[0]),
    .ZN(_14030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22995_ (.A1(_13988_),
    .A2(net19254),
    .A3(_14030_),
    .ZN(_14031_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _22996_ (.A1(net18809),
    .A2(_15822_[0]),
    .Z(_14032_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22997_ (.A1(_13998_),
    .A2(net19237),
    .A3(_14032_),
    .ZN(_14033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22998_ (.A1(_14031_),
    .A2(_14033_),
    .A3(net20254),
    .ZN(_14034_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22999_ (.A1(net20635),
    .A2(_14034_),
    .A3(_14029_),
    .ZN(_14035_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23000_ (.A1(_14035_),
    .A2(_14019_),
    .A3(net20633),
    .ZN(_14036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23001_ (.A1(_14036_),
    .A2(_14002_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23002_ (.A1(net18806),
    .A2(_13847_),
    .Z(_14037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23003_ (.A1(_14037_),
    .A2(net18255),
    .ZN(_14038_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23004_ (.A1(_13898_),
    .A2(_14038_),
    .A3(net19254),
    .ZN(_14039_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _23005_ (.A1(_13719_),
    .A2(_13724_),
    .A3(net19233),
    .Z(_14040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23006_ (.A1(net18817),
    .A2(net19800),
    .ZN(_14041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23007_ (.A1(_14040_),
    .A2(_14041_),
    .ZN(_14042_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23008_ (.A1(_14039_),
    .A2(net20252),
    .A3(_14042_),
    .Z(_14043_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23009_ (.A1(_14043_),
    .A2(net20635),
    .ZN(_14044_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _23010_ (.A1(_13895_),
    .A2(net18824),
    .A3(_13837_),
    .Z(_14045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23011_ (.A1(_13753_),
    .A2(net18816),
    .Z(_14046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23012_ (.A1(_13724_),
    .A2(_13675_),
    .Z(_14047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23013_ (.A1(_14046_),
    .A2(_14047_),
    .ZN(_14048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23014_ (.A1(_14045_),
    .A2(_14048_),
    .A3(net19236),
    .ZN(_14049_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _23015_ (.I(_13710_),
    .ZN(_14050_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23016_ (.A1(_14050_),
    .A2(_13760_),
    .B(_13725_),
    .C(net19252),
    .ZN(_14051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23017_ (.A1(_14049_),
    .A2(_14051_),
    .ZN(_14052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23018_ (.A1(_14052_),
    .A2(net20030),
    .ZN(_14053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23019_ (.A1(_14053_),
    .A2(_14044_),
    .ZN(_14054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23020_ (.A1(net17880),
    .A2(net17883),
    .ZN(_14055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23021_ (.A1(_14055_),
    .A2(net18823),
    .ZN(_14056_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23022_ (.A1(net18823),
    .A2(_14047_),
    .B(_14056_),
    .C(net19250),
    .ZN(_14057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23023_ (.A1(_13787_),
    .A2(_13976_),
    .ZN(_14058_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23024_ (.A1(_14058_),
    .A2(net17870),
    .A3(net19233),
    .ZN(_14059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23025_ (.A1(_14057_),
    .A2(_14059_),
    .A3(net20029),
    .ZN(_14060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23026_ (.A1(_14015_),
    .A2(net18808),
    .ZN(_14061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23027_ (.A1(_14061_),
    .A2(_13752_),
    .B(_13739_),
    .ZN(_14062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23028_ (.A1(_13716_),
    .A2(net18802),
    .ZN(_14063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23029_ (.A1(_13766_),
    .A2(net18801),
    .ZN(_14064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23030_ (.A1(_14063_),
    .A2(_14064_),
    .A3(net19233),
    .ZN(_14065_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23031_ (.A1(_14065_),
    .A2(_14062_),
    .B(_13881_),
    .ZN(_14066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23032_ (.A1(_14060_),
    .A2(_14066_),
    .B(net20805),
    .ZN(_14067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23033_ (.A1(_14054_),
    .A2(_14067_),
    .ZN(_14068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23034_ (.A1(net17872),
    .A2(net18818),
    .ZN(_14069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23035_ (.A1(_13739_),
    .A2(_14069_),
    .Z(_14070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23036_ (.A1(_14070_),
    .A2(net17531),
    .B(net19248),
    .ZN(_14071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23037_ (.A1(_13781_),
    .A2(_13803_),
    .Z(_14072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23038_ (.A1(net19799),
    .A2(_14072_),
    .ZN(_14073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23039_ (.A1(_14073_),
    .A2(net18813),
    .Z(_14074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23040_ (.A1(_14074_),
    .A2(net17876),
    .ZN(_14075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23041_ (.A1(net18268),
    .A2(net17885),
    .ZN(_14076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23042_ (.A1(_14075_),
    .A2(_14076_),
    .A3(net20250),
    .ZN(_14077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23043_ (.A1(_14071_),
    .A2(_14077_),
    .B(_13881_),
    .ZN(_14078_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _23044_ (.A1(net18259),
    .A2(_13852_),
    .B1(net18806),
    .B2(net17882),
    .ZN(_14079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23045_ (.A1(_14079_),
    .A2(net20251),
    .ZN(_14080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23046_ (.I(_13758_),
    .ZN(_14081_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _23047_ (.A1(_14081_),
    .A2(net20025),
    .B1(net18821),
    .B2(net407),
    .ZN(_14082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23048_ (.A1(_14080_),
    .A2(_14082_),
    .ZN(_14083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23049_ (.A1(_14083_),
    .A2(net19248),
    .ZN(_14084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23050_ (.A1(_14078_),
    .A2(_14084_),
    .ZN(_14085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23051_ (.I(_13811_),
    .ZN(_14086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _23052_ (.A1(net19232),
    .A2(_13861_),
    .B(net18818),
    .ZN(_14087_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23053_ (.A1(_14050_),
    .A2(net17529),
    .B(_14087_),
    .C(net19252),
    .ZN(_14088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23054_ (.A1(_13831_),
    .A2(_13918_),
    .A3(net19236),
    .ZN(_14089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23055_ (.A1(_14088_),
    .A2(_14089_),
    .A3(net20026),
    .ZN(_14090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23056_ (.A1(_14074_),
    .A2(net634),
    .ZN(_14091_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23057_ (.A1(_13940_),
    .A2(_14091_),
    .A3(net19234),
    .ZN(_14092_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23058_ (.I(_13971_),
    .ZN(_14093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23059_ (.A1(_14093_),
    .A2(net19248),
    .B(net20027),
    .ZN(_14094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23060_ (.A1(_14092_),
    .A2(_14094_),
    .B(net20634),
    .ZN(_14095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23061_ (.A1(_14090_),
    .A2(_14095_),
    .ZN(_14096_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23062_ (.A1(_14085_),
    .A2(_14096_),
    .A3(net20805),
    .ZN(_14097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23063_ (.A1(_14068_),
    .A2(_14097_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _23064_ (.A1(net19253),
    .A2(_13935_),
    .A3(_13755_),
    .A4(_14025_),
    .ZN(_14098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23065_ (.A1(net18271),
    .A2(net17876),
    .B(net18252),
    .ZN(_14099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23066_ (.A1(_14099_),
    .A2(net19233),
    .ZN(_14100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23067_ (.A1(_14098_),
    .A2(_14100_),
    .A3(net20252),
    .ZN(_14101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23068_ (.A1(_13913_),
    .A2(net18261),
    .ZN(_14102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23069_ (.A1(_13780_),
    .A2(net19237),
    .A3(_14102_),
    .ZN(_14103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23070_ (.A1(_13947_),
    .A2(net18806),
    .ZN(_14104_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23071_ (.A1(_14104_),
    .A2(net19254),
    .Z(_14105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23072_ (.A1(_13711_),
    .A2(net18826),
    .ZN(_14106_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23073_ (.A1(_14105_),
    .A2(_14106_),
    .B(net20249),
    .ZN(_14107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23074_ (.A1(_14103_),
    .A2(_14107_),
    .ZN(_14108_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23075_ (.A1(_14101_),
    .A2(_13881_),
    .A3(_14108_),
    .ZN(_14109_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23076_ (.I(_15815_[0]),
    .ZN(_14110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23077_ (.A1(net18810),
    .A2(_14110_),
    .ZN(_14111_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _23078_ (.A1(_14003_),
    .A2(_14111_),
    .A3(net19233),
    .Z(_14112_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23079_ (.A1(_14112_),
    .A2(net20252),
    .ZN(_14113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23080_ (.A1(_13848_),
    .A2(net18796),
    .ZN(_14114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23081_ (.A1(_14114_),
    .A2(net18265),
    .A3(net19258),
    .ZN(_14115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23082_ (.A1(_14113_),
    .A2(_14115_),
    .B(_13881_),
    .ZN(_14116_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23083_ (.A1(net18802),
    .A2(net18801),
    .A3(net18806),
    .ZN(_14117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23084_ (.A1(_13848_),
    .A2(net19245),
    .ZN(_14118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23085_ (.A1(_14117_),
    .A2(_14118_),
    .A3(net19252),
    .ZN(_14119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23086_ (.A1(_13878_),
    .A2(_13725_),
    .A3(net19233),
    .ZN(_14120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23087_ (.A1(_14119_),
    .A2(_14120_),
    .A3(net20253),
    .ZN(_14121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23088_ (.A1(_14116_),
    .A2(_14121_),
    .B(_13821_),
    .ZN(_14122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23089_ (.A1(_14109_),
    .A2(_14122_),
    .ZN(_14123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23090_ (.A1(_13827_),
    .A2(net19258),
    .Z(_14124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23091_ (.A1(net637),
    .A2(_13953_),
    .Z(_14125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23092_ (.A1(_14125_),
    .A2(_14124_),
    .B(net20249),
    .ZN(_14126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23093_ (.A1(_13946_),
    .A2(net17883),
    .ZN(_14127_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23094_ (.A1(_13849_),
    .A2(net19239),
    .A3(_14127_),
    .ZN(_14128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23095_ (.A1(_14128_),
    .A2(_14126_),
    .B(_13881_),
    .ZN(_14129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23096_ (.A1(_13845_),
    .A2(net18824),
    .A3(net18800),
    .ZN(_14130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23097_ (.A1(_13990_),
    .A2(net19258),
    .Z(_14131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23098_ (.A1(_14130_),
    .A2(_14131_),
    .B(net20032),
    .ZN(_14132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23099_ (.A1(_13922_),
    .A2(net17880),
    .ZN(_14133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23100_ (.A1(_14133_),
    .A2(net18829),
    .ZN(_14134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23101_ (.A1(_13828_),
    .A2(net19240),
    .A3(_14134_),
    .ZN(_14135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23102_ (.A1(_14132_),
    .A2(_14135_),
    .ZN(_14136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23103_ (.A1(_14136_),
    .A2(_14129_),
    .ZN(_14137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23104_ (.A1(_13975_),
    .A2(_13767_),
    .ZN(_14138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23105_ (.A1(net19262),
    .A2(net19805),
    .ZN(_14139_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23106_ (.A1(_14139_),
    .A2(net18795),
    .A3(net18807),
    .ZN(_14140_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23107_ (.A1(_14138_),
    .A2(net19258),
    .A3(_14140_),
    .ZN(_14141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23108_ (.A1(_14007_),
    .A2(net19239),
    .A3(_13934_),
    .ZN(_14142_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23109_ (.A1(_14141_),
    .A2(_14142_),
    .A3(net20249),
    .ZN(_14143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23110_ (.A1(_13922_),
    .A2(net18813),
    .A3(_13808_),
    .ZN(_14144_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23111_ (.A1(_13932_),
    .A2(_14144_),
    .A3(net19239),
    .ZN(_14145_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23112_ (.A1(_14021_),
    .A2(net19258),
    .Z(_14146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23113_ (.I(_13848_),
    .ZN(_14147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23114_ (.A1(_14146_),
    .A2(_14147_),
    .B(net20249),
    .ZN(_14148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23115_ (.A1(_14145_),
    .A2(_14148_),
    .B(net20634),
    .ZN(_14149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23116_ (.A1(_14143_),
    .A2(_14149_),
    .ZN(_14150_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23117_ (.A1(_13821_),
    .A2(_14150_),
    .A3(_14137_),
    .ZN(_14151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23118_ (.A1(_14151_),
    .A2(_14123_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23119_ (.A1(net18813),
    .A2(net18409),
    .Z(_14152_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23120_ (.A1(_13856_),
    .A2(_14152_),
    .ZN(_14153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23121_ (.A1(_13845_),
    .A2(_14037_),
    .ZN(_14154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23122_ (.A1(_14153_),
    .A2(_14154_),
    .ZN(_14155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23123_ (.A1(_13989_),
    .A2(net18831),
    .ZN(_14156_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23124_ (.A1(_13783_),
    .A2(_14156_),
    .A3(_13755_),
    .ZN(_14157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23125_ (.A1(_14155_),
    .A2(_14157_),
    .A3(_13739_),
    .ZN(_14158_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23126_ (.A1(_14087_),
    .A2(_14050_),
    .A3(net19235),
    .ZN(_14159_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23127_ (.A1(_13913_),
    .A2(net19233),
    .ZN(_14160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23128_ (.A1(_13916_),
    .A2(_13721_),
    .ZN(_14161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23129_ (.A1(_14160_),
    .A2(_14161_),
    .ZN(_14162_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23130_ (.A1(_14159_),
    .A2(_14162_),
    .A3(net20250),
    .ZN(_14163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23131_ (.A1(_14163_),
    .A2(_14158_),
    .ZN(_14164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23132_ (.A1(_14164_),
    .A2(_13881_),
    .ZN(_14165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23133_ (.A1(net18813),
    .A2(net19262),
    .ZN(_14166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23134_ (.A1(_14140_),
    .A2(_14166_),
    .ZN(_14167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23135_ (.A1(_14167_),
    .A2(net19234),
    .ZN(_14168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23136_ (.A1(net18267),
    .A2(_14139_),
    .B(net19233),
    .ZN(_14169_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23137_ (.A1(net19246),
    .A2(net19242),
    .B(_13851_),
    .ZN(_14170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23138_ (.A1(_14170_),
    .A2(net18814),
    .ZN(_14171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23139_ (.A1(_14169_),
    .A2(_14171_),
    .ZN(_14172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23140_ (.A1(_14168_),
    .A2(_14172_),
    .A3(net20027),
    .ZN(_14173_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23141_ (.A1(net18259),
    .A2(_14104_),
    .ZN(_14174_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23142_ (.I(_13953_),
    .ZN(_14175_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23143_ (.A1(_14174_),
    .A2(_14175_),
    .B(net19252),
    .ZN(_14176_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23144_ (.A1(_13673_),
    .A2(net17536),
    .B(_13980_),
    .C(net19233),
    .ZN(_14177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23145_ (.A1(_14176_),
    .A2(_14177_),
    .A3(net20250),
    .ZN(_14178_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23146_ (.A1(_14173_),
    .A2(_14178_),
    .A3(net20634),
    .ZN(_14179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23147_ (.A1(_14165_),
    .A2(_14179_),
    .ZN(_14180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23148_ (.A1(_14180_),
    .A2(_13821_),
    .ZN(_14181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23149_ (.A1(_13776_),
    .A2(net18809),
    .ZN(_14182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23150_ (.A1(_13760_),
    .A2(net18825),
    .ZN(_14183_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23151_ (.A1(_14182_),
    .A2(net17529),
    .B(net19254),
    .C(_14183_),
    .ZN(_14184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23152_ (.A1(net18798),
    .A2(net18809),
    .ZN(_14185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23153_ (.A1(_13780_),
    .A2(_13866_),
    .A3(_14185_),
    .ZN(_14186_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23154_ (.A1(_14184_),
    .A2(_14186_),
    .A3(net20250),
    .ZN(_14187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23155_ (.A1(net19805),
    .A2(net18819),
    .B(_13669_),
    .ZN(_14188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23156_ (.A1(_13720_),
    .A2(_14188_),
    .B(net20250),
    .ZN(_14189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23157_ (.A1(_13766_),
    .A2(net410),
    .ZN(_14190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23158_ (.A1(_14037_),
    .A2(net18795),
    .ZN(_14191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23159_ (.A1(_14190_),
    .A2(_14191_),
    .A3(net19257),
    .ZN(_14192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23160_ (.A1(_14189_),
    .A2(_14192_),
    .B(net20634),
    .ZN(_14193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23161_ (.A1(_14187_),
    .A2(_14193_),
    .ZN(_14194_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23162_ (.I(_13812_),
    .ZN(_14195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23163_ (.A1(_14124_),
    .A2(_14195_),
    .B(net20249),
    .ZN(_14196_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23164_ (.I(net18270),
    .ZN(_14197_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23165_ (.A1(_14074_),
    .A2(net19252),
    .ZN(_14198_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23166_ (.A1(_14197_),
    .A2(_13998_),
    .B(_14198_),
    .ZN(_14199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23167_ (.A1(_14196_),
    .A2(_14199_),
    .ZN(_14200_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23168_ (.I(_13903_),
    .ZN(_14201_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _23169_ (.A1(_14201_),
    .A2(_14086_),
    .A3(net18826),
    .Z(_14202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23170_ (.A1(_13766_),
    .A2(net18258),
    .ZN(_14203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23171_ (.A1(_14202_),
    .A2(net19254),
    .A3(_14203_),
    .ZN(_14204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23172_ (.A1(net18272),
    .A2(net18825),
    .B(net19255),
    .ZN(_14205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23173_ (.A1(_14182_),
    .A2(_14205_),
    .B(_13739_),
    .ZN(_14206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23174_ (.A1(_14204_),
    .A2(_14206_),
    .ZN(_14207_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23175_ (.A1(_14200_),
    .A2(_14207_),
    .A3(net20635),
    .ZN(_14208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23176_ (.A1(_14194_),
    .A2(_14208_),
    .A3(net20805),
    .ZN(_14209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23177_ (.A1(_14181_),
    .A2(_14209_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23178_ (.A1(_14006_),
    .A2(_13946_),
    .B(_13724_),
    .ZN(_14210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23179_ (.A1(_14210_),
    .A2(net19250),
    .ZN(_14211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23180_ (.A1(net18806),
    .A2(net430),
    .ZN(_14212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23181_ (.A1(_14040_),
    .A2(net18251),
    .B(net20251),
    .ZN(_14213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23182_ (.A1(_14211_),
    .A2(_14213_),
    .ZN(_14214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23183_ (.A1(net17869),
    .A2(net18811),
    .ZN(_14215_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23184_ (.A1(_14087_),
    .A2(net19238),
    .A3(_14215_),
    .ZN(_14216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23185_ (.A1(_13923_),
    .A2(_13810_),
    .ZN(_14217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23186_ (.A1(_14216_),
    .A2(_14217_),
    .A3(net20249),
    .ZN(_14218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23187_ (.A1(_14218_),
    .A2(_14214_),
    .B(net20635),
    .ZN(_14219_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23188_ (.A1(_13979_),
    .A2(net19239),
    .A3(net18796),
    .ZN(_14220_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23189_ (.A1(_14114_),
    .A2(net19258),
    .A3(net17873),
    .ZN(_14221_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23190_ (.A1(_14220_),
    .A2(_14221_),
    .A3(net20249),
    .ZN(_14222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23191_ (.A1(net17533),
    .A2(net18255),
    .ZN(_14223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23192_ (.A1(_13952_),
    .A2(_14223_),
    .ZN(_14224_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23193_ (.I(_15821_[0]),
    .ZN(_14225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23194_ (.A1(_14225_),
    .A2(net18814),
    .B(net19249),
    .ZN(_14226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23195_ (.A1(_14226_),
    .A2(_14191_),
    .ZN(_14227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23196_ (.A1(_14224_),
    .A2(net20032),
    .A3(_14227_),
    .ZN(_14228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23197_ (.A1(_14228_),
    .A2(_14222_),
    .B(_13881_),
    .ZN(_14229_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23198_ (.A1(_14219_),
    .A2(_14229_),
    .B(net20805),
    .ZN(_14230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23199_ (.A1(_13916_),
    .A2(_14139_),
    .ZN(_14231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23200_ (.A1(net17878),
    .A2(_13847_),
    .A3(net18806),
    .ZN(_14232_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23201_ (.A1(_14231_),
    .A2(_13855_),
    .A3(_14232_),
    .ZN(_14233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23202_ (.A1(_14233_),
    .A2(net19233),
    .ZN(_14234_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23203_ (.A1(_13968_),
    .A2(net18263),
    .Z(_14235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23204_ (.A1(_14235_),
    .A2(net18822),
    .A3(_13826_),
    .ZN(_14236_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23205_ (.A1(_14185_),
    .A2(_13838_),
    .A3(_14236_),
    .ZN(_14237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23206_ (.A1(_14234_),
    .A2(_14237_),
    .ZN(_14238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23207_ (.A1(_14238_),
    .A2(net20252),
    .ZN(_14239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23208_ (.A1(_14046_),
    .A2(net18802),
    .ZN(_14240_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23209_ (.A1(_15820_[0]),
    .A2(_15829_[0]),
    .Z(_14241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23210_ (.A1(net18810),
    .A2(_14241_),
    .B(net19250),
    .ZN(_14242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23211_ (.A1(_14242_),
    .A2(_14240_),
    .B(net20251),
    .ZN(_14243_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23212_ (.A1(net18806),
    .A2(_14235_),
    .B(net17317),
    .C(net19252),
    .ZN(_14244_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23213_ (.A1(_14243_),
    .A2(_14244_),
    .B(net20635),
    .ZN(_14245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23214_ (.A1(_14245_),
    .A2(_14239_),
    .ZN(_14246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23215_ (.A1(_13916_),
    .A2(net19801),
    .B(net19250),
    .ZN(_14247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23216_ (.A1(_13887_),
    .A2(net17530),
    .ZN(_14248_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23217_ (.A1(_14247_),
    .A2(_13725_),
    .A3(_14248_),
    .ZN(_14249_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23218_ (.A1(net18804),
    .A2(net18791),
    .A3(net18825),
    .ZN(_14250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23219_ (.A1(_13760_),
    .A2(net18809),
    .B(net19233),
    .ZN(_14251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23220_ (.A1(_14250_),
    .A2(_14251_),
    .B(net20030),
    .ZN(_14252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23221_ (.A1(_14249_),
    .A2(_14252_),
    .B(_13881_),
    .ZN(_14253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23222_ (.A1(_13975_),
    .A2(net18794),
    .ZN(_14254_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23223_ (.A1(_14104_),
    .A2(_14201_),
    .Z(_14255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23224_ (.A1(_14255_),
    .A2(net19237),
    .A3(_14254_),
    .ZN(_14256_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23225_ (.A1(net631),
    .A2(net18811),
    .A3(net17885),
    .ZN(_14257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23226_ (.A1(_14257_),
    .A2(net19254),
    .A3(_14032_),
    .ZN(_14258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23227_ (.A1(_14256_),
    .A2(_14258_),
    .A3(net20032),
    .ZN(_14259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23228_ (.A1(_14259_),
    .A2(_14253_),
    .ZN(_14260_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23229_ (.A1(_14246_),
    .A2(_14260_),
    .A3(net20633),
    .ZN(_14261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23230_ (.A1(_14261_),
    .A2(_14230_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23231_ (.A1(net19805),
    .A2(net18819),
    .B(_14144_),
    .ZN(_14262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23232_ (.A1(_14262_),
    .A2(net19257),
    .ZN(_14263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23233_ (.A1(_13795_),
    .A2(_13711_),
    .ZN(_14264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23234_ (.A1(_14264_),
    .A2(_14007_),
    .A3(net19238),
    .ZN(_14265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23235_ (.A1(_14263_),
    .A2(_14265_),
    .A3(net20024),
    .ZN(_14266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23236_ (.A1(net603),
    .A2(net18831),
    .ZN(_14267_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23237_ (.A1(_13711_),
    .A2(net18808),
    .A3(net18254),
    .ZN(_14268_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23238_ (.A1(_14267_),
    .A2(_14268_),
    .A3(net19258),
    .ZN(_14269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23239_ (.A1(_13758_),
    .A2(net19233),
    .Z(_14270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23240_ (.A1(_13895_),
    .A2(net18830),
    .ZN(_14271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23241_ (.A1(_14270_),
    .A2(_14271_),
    .B(net20031),
    .ZN(_14272_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23242_ (.A1(_14272_),
    .A2(_14269_),
    .B(_13881_),
    .ZN(_14273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23243_ (.A1(_14266_),
    .A2(_14273_),
    .B(_13821_),
    .ZN(_14274_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _23244_ (.A1(_14020_),
    .A2(_13762_),
    .Z(_14275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23245_ (.A1(_14275_),
    .A2(net18821),
    .ZN(_14276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23246_ (.A1(net17874),
    .A2(net18268),
    .B(net19239),
    .ZN(_14277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23247_ (.A1(_14276_),
    .A2(_14277_),
    .ZN(_14278_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23248_ (.I(_13946_),
    .ZN(_14279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23249_ (.A1(_14114_),
    .A2(net19239),
    .A3(_14279_),
    .ZN(_14280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23250_ (.A1(_14278_),
    .A2(_13739_),
    .A3(_14280_),
    .ZN(_14281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23251_ (.A1(_14016_),
    .A2(net19233),
    .A3(net17528),
    .ZN(_14282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23252_ (.A1(_13925_),
    .A2(_14076_),
    .A3(net19257),
    .ZN(_14283_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23253_ (.A1(_14282_),
    .A2(_14283_),
    .A3(net20249),
    .ZN(_14284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23254_ (.A1(_14281_),
    .A2(_13881_),
    .A3(_14284_),
    .ZN(_14285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23255_ (.A1(_14274_),
    .A2(_14285_),
    .ZN(_14286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23256_ (.A1(net18815),
    .A2(_14110_),
    .ZN(_14287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23257_ (.A1(_13834_),
    .A2(_14287_),
    .B(net20251),
    .ZN(_14288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23258_ (.A1(_14212_),
    .A2(_13669_),
    .Z(_14289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23259_ (.A1(_13935_),
    .A2(_14289_),
    .A3(_14185_),
    .ZN(_14290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23260_ (.A1(_14288_),
    .A2(_14290_),
    .B(_13881_),
    .ZN(_14291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23261_ (.A1(_14011_),
    .A2(net18254),
    .ZN(_14292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23262_ (.A1(net18268),
    .A2(net18795),
    .ZN(_14293_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23263_ (.A1(_14292_),
    .A2(_14293_),
    .A3(net19248),
    .ZN(_14294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23264_ (.A1(net17882),
    .A2(_13968_),
    .Z(_14295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23265_ (.A1(net18815),
    .A2(_15829_[0]),
    .ZN(_14296_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23266_ (.A1(_14295_),
    .A2(net18814),
    .B(net19235),
    .C(_14296_),
    .ZN(_14297_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23267_ (.A1(_14294_),
    .A2(_14297_),
    .A3(net20251),
    .ZN(_14298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23268_ (.A1(_14291_),
    .A2(_14298_),
    .B(net20805),
    .ZN(_14299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23269_ (.A1(_14275_),
    .A2(net18806),
    .ZN(_14300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23270_ (.A1(net18254),
    .A2(net18258),
    .A3(net18822),
    .ZN(_14301_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23271_ (.A1(_14300_),
    .A2(net19235),
    .A3(_14301_),
    .ZN(_14302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23272_ (.A1(net19232),
    .A2(net18807),
    .ZN(_14303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23273_ (.A1(_14289_),
    .A2(_14303_),
    .Z(_14304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23274_ (.A1(_14304_),
    .A2(_14091_),
    .B(net20251),
    .ZN(_14305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23275_ (.A1(_14302_),
    .A2(_14305_),
    .ZN(_14306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23276_ (.A1(net18806),
    .A2(net18409),
    .ZN(_14307_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23277_ (.A1(_14240_),
    .A2(net19250),
    .A3(_14307_),
    .ZN(_14308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23278_ (.A1(_13754_),
    .A2(net18815),
    .ZN(_14309_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23279_ (.A1(_13834_),
    .A2(net17880),
    .A3(_14309_),
    .ZN(_14310_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23280_ (.A1(_14308_),
    .A2(_14310_),
    .A3(net20251),
    .ZN(_14311_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23281_ (.A1(_14306_),
    .A2(_14311_),
    .A3(_13881_),
    .ZN(_14312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23282_ (.A1(_14299_),
    .A2(_14312_),
    .ZN(_14313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23283_ (.A1(_14286_),
    .A2(_14313_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23284_ (.I(\sa21_sr[7] ),
    .ZN(_14314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23285_ (.A1(_14314_),
    .A2(net21359),
    .ZN(_14315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23286_ (.A1(net21346),
    .A2(_11194_),
    .ZN(_14316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23287_ (.A1(_14316_),
    .A2(_14315_),
    .ZN(_14317_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23288_ (.A1(_14317_),
    .A2(_11161_),
    .Z(_14318_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23289_ (.A1(_11161_),
    .A2(_14317_),
    .ZN(_14319_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23290_ (.A1(_14318_),
    .A2(_14319_),
    .ZN(_14320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23291_ (.A1(_11174_),
    .A2(net21040),
    .ZN(_14321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23292_ (.A1(_11170_),
    .A2(net21466),
    .ZN(_14322_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23293_ (.A1(_14321_),
    .A2(_14322_),
    .Z(_14323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23294_ (.A1(_14320_),
    .A2(_14323_),
    .ZN(_14324_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23295_ (.A1(_11194_),
    .A2(_14314_),
    .ZN(_14325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23296_ (.A1(net21359),
    .A2(\sa21_sr[7] ),
    .ZN(_14326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23297_ (.A1(_14325_),
    .A2(_14326_),
    .ZN(_14327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23298_ (.A1(_11147_),
    .A2(_14327_),
    .ZN(_14328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23299_ (.A1(_11161_),
    .A2(_14317_),
    .ZN(_14329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23300_ (.A1(_14328_),
    .A2(_14329_),
    .ZN(_14330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23301_ (.A1(_14321_),
    .A2(_14322_),
    .ZN(_14331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23302_ (.A1(_14330_),
    .A2(_14331_),
    .ZN(_14332_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17248 (.I(_03501_),
    .Z(net17248));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23304_ (.A1(_14324_),
    .A2(_14332_),
    .A3(_10378_),
    .ZN(_14334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23305_ (.A1(net21493),
    .A2(\text_in_r[81] ),
    .ZN(_14335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23306_ (.A1(_14334_),
    .A2(_14335_),
    .ZN(_14336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23307_ (.A1(net20023),
    .A2(_07874_),
    .ZN(_14337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23308_ (.A1(net20247),
    .A2(net21202),
    .A3(net20980),
    .ZN(_14338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23309_ (.A1(_14338_),
    .A2(_14337_),
    .ZN(_15839_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23310_ (.A1(net21044),
    .A2(net21297),
    .ZN(_14339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23311_ (.A1(net21042),
    .A2(net21401),
    .ZN(_14340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23312_ (.A1(_14339_),
    .A2(_14340_),
    .ZN(_14341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23313_ (.A1(_14341_),
    .A2(net21467),
    .ZN(_14342_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23314_ (.A1(_14339_),
    .A2(_14340_),
    .A3(net21047),
    .ZN(_14343_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23315_ (.A1(_14342_),
    .A2(_14343_),
    .A3(net20884),
    .ZN(_14344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23316_ (.A1(net21467),
    .A2(net21401),
    .ZN(_14345_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23317_ (.I(_14345_),
    .ZN(_14346_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23318_ (.A1(net21467),
    .A2(net21402),
    .ZN(_14347_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23319_ (.A1(_14346_),
    .A2(_14347_),
    .B(net21297),
    .ZN(_14348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23320_ (.A1(net21047),
    .A2(net21044),
    .ZN(_14349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23321_ (.A1(_14349_),
    .A2(net21042),
    .A3(_14345_),
    .ZN(_14350_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23322_ (.A1(_14348_),
    .A2(_14350_),
    .A3(_14327_),
    .ZN(_14351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23323_ (.A1(_14344_),
    .A2(_14351_),
    .B(net21493),
    .ZN(_14352_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23324_ (.I(\text_in_r[80] ),
    .ZN(_14353_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23325_ (.A1(_14353_),
    .A2(net21493),
    .Z(_14354_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23326_ (.A1(net20437),
    .A2(net20936),
    .B(net21203),
    .ZN(_14355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23327_ (.A1(_14344_),
    .A2(_14351_),
    .ZN(_14356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23328_ (.A1(_14356_),
    .A2(_10378_),
    .ZN(_14357_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23329_ (.I(_14354_),
    .ZN(_14358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23330_ (.A1(net20246),
    .A2(_07869_),
    .A3(net20883),
    .ZN(_14359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23331_ (.A1(_14355_),
    .A2(_14359_),
    .ZN(_15842_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23332_ (.A1(net21355),
    .A2(\sa30_sub[2] ),
    .Z(_14360_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23333_ (.A1(net21355),
    .A2(net21293),
    .ZN(_14361_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23334_ (.A1(_14360_),
    .A2(_14361_),
    .B(net21463),
    .ZN(_14362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23335_ (.A1(_11216_),
    .A2(_11221_),
    .ZN(_14363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23336_ (.A1(net21356),
    .A2(net21293),
    .ZN(_14364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23337_ (.A1(_14363_),
    .A2(_11250_),
    .A3(_14364_),
    .ZN(_14365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23338_ (.A1(_14362_),
    .A2(_14365_),
    .ZN(_14366_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23339_ (.A1(net21409),
    .A2(net21357),
    .ZN(_14367_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23340_ (.I(_14367_),
    .ZN(_14368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23341_ (.A1(_14366_),
    .A2(_14368_),
    .ZN(_14369_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23342_ (.A1(_14362_),
    .A2(_14365_),
    .A3(_14367_),
    .ZN(_14370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23343_ (.A1(_14369_),
    .A2(_14370_),
    .B(net21499),
    .ZN(_14371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23344_ (.I(\text_in_r[82] ),
    .ZN(_14372_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23345_ (.A1(_14372_),
    .A2(net21493),
    .Z(_14373_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23346_ (.A1(_14371_),
    .A2(_14373_),
    .B(_07879_),
    .ZN(_14374_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23347_ (.A1(_14369_),
    .A2(_14370_),
    .ZN(_14375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23348_ (.A1(_14375_),
    .A2(net21073),
    .ZN(_14376_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23349_ (.I(_14373_),
    .ZN(_14377_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23350_ (.A1(_14376_),
    .A2(net21201),
    .A3(_14377_),
    .ZN(_14378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23351_ (.A1(_14374_),
    .A2(_14378_),
    .ZN(_14379_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17243 (.I(_04007_),
    .Z(net17243));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23353_ (.A1(_14352_),
    .A2(_14354_),
    .B(_07869_),
    .ZN(_14380_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23354_ (.A1(_14357_),
    .A2(net21203),
    .A3(_14358_),
    .ZN(_14381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23355_ (.A1(_14380_),
    .A2(_14381_),
    .ZN(_15833_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23356_ (.A1(_14371_),
    .A2(_14373_),
    .B(net21201),
    .ZN(_14382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23357_ (.A1(_14376_),
    .A2(_07879_),
    .A3(_14377_),
    .ZN(_14383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23358_ (.A1(_14382_),
    .A2(_14383_),
    .ZN(_14384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17241 (.I(_04086_),
    .Z(net17241));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17246 (.I(_03570_),
    .Z(net17246));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23361_ (.I(_15836_[0]),
    .ZN(_14386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23362_ (.A1(net19788),
    .A2(net18250),
    .ZN(_14387_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23363_ (.I(_14387_),
    .ZN(_14388_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23364_ (.A1(net21354),
    .A2(net21347),
    .Z(_14389_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23365_ (.A1(_14389_),
    .A2(_11262_),
    .ZN(_14390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23366_ (.A1(_11216_),
    .A2(net20981),
    .ZN(_14391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23367_ (.A1(\sa21_sr[2] ),
    .A2(net21347),
    .ZN(_14392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23368_ (.A1(_14391_),
    .A2(_14392_),
    .ZN(_14393_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23369_ (.A1(_11249_),
    .A2(_14393_),
    .ZN(_14394_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23370_ (.A1(_14390_),
    .A2(_14394_),
    .ZN(_14395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23371_ (.A1(net21044),
    .A2(net21036),
    .ZN(_14396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23372_ (.A1(net21402),
    .A2(net21408),
    .ZN(_14397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23373_ (.A1(_14396_),
    .A2(_14397_),
    .ZN(_14398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23374_ (.A1(_14398_),
    .A2(net21462),
    .ZN(_14399_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23375_ (.I(\sa01_sr[3] ),
    .ZN(_14400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23376_ (.A1(_14396_),
    .A2(net20979),
    .A3(_14397_),
    .ZN(_14401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23377_ (.A1(_14399_),
    .A2(_14401_),
    .ZN(_14402_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23378_ (.I(_14402_),
    .ZN(_14403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23379_ (.A1(_14395_),
    .A2(_14403_),
    .ZN(_14404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23380_ (.A1(_11249_),
    .A2(_14393_),
    .ZN(_14405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23381_ (.A1(_14389_),
    .A2(_11262_),
    .ZN(_14406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23382_ (.A1(_14405_),
    .A2(_14406_),
    .ZN(_14407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23383_ (.A1(_14407_),
    .A2(_14402_),
    .ZN(_14408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23384_ (.A1(_14404_),
    .A2(_14408_),
    .A3(net21071),
    .ZN(_14409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23385_ (.A1(net21496),
    .A2(\text_in_r[83] ),
    .ZN(_14410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23386_ (.A1(_14409_),
    .A2(_14410_),
    .ZN(_14411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23387_ (.A1(_14411_),
    .A2(_07884_),
    .ZN(_14412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23388_ (.A1(_14409_),
    .A2(net21200),
    .A3(_14410_),
    .ZN(_14413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23389_ (.A1(_14412_),
    .A2(_14413_),
    .ZN(_14414_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17250 (.I(_03449_),
    .Z(net17250));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23391_ (.A1(_14388_),
    .A2(net18771),
    .ZN(_14416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23392_ (.A1(_11258_),
    .A2(net20981),
    .ZN(_14417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23393_ (.A1(\sa21_sr[3] ),
    .A2(net21347),
    .ZN(_14418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23394_ (.A1(_14417_),
    .A2(_14418_),
    .ZN(_14419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23395_ (.A1(_11305_),
    .A2(_14419_),
    .ZN(_14420_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23396_ (.I(_14419_),
    .ZN(_14421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23397_ (.A1(_14421_),
    .A2(net20951),
    .ZN(_14422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23398_ (.A1(_14420_),
    .A2(_14422_),
    .ZN(_14423_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23399_ (.A1(_11273_),
    .A2(net21461),
    .Z(_14424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23400_ (.A1(_11273_),
    .A2(net21461),
    .ZN(_14425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23401_ (.A1(_14424_),
    .A2(_14425_),
    .ZN(_14426_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23402_ (.A1(_14423_),
    .A2(_14426_),
    .Z(_14427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23403_ (.A1(_14423_),
    .A2(_14426_),
    .ZN(_14428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23404_ (.A1(_14427_),
    .A2(net21071),
    .A3(_14428_),
    .ZN(_14429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23405_ (.A1(net21496),
    .A2(\text_in_r[84] ),
    .ZN(_14430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23406_ (.A1(_14429_),
    .A2(_14430_),
    .ZN(_14431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23407_ (.A1(_14431_),
    .A2(net21198),
    .ZN(_14432_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23408_ (.A1(_14429_),
    .A2(_07888_),
    .A3(_14430_),
    .ZN(_14433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23409_ (.A1(_14432_),
    .A2(_14433_),
    .ZN(_14434_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _23410_ (.I(_14434_),
    .ZN(_14435_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17253 (.I(_03411_),
    .Z(net17253));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23412_ (.A1(_14416_),
    .A2(net18240),
    .Z(_14437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23413_ (.A1(net20245),
    .A2(_14386_),
    .A3(net20022),
    .ZN(_14438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23414_ (.A1(_14411_),
    .A2(net21200),
    .ZN(_14439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23415_ (.A1(net20020),
    .A2(_07884_),
    .A3(net20978),
    .ZN(_14440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23416_ (.A1(_14439_),
    .A2(_14440_),
    .ZN(_14441_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19450 (.I(net19446),
    .Z(net19450));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23418_ (.A1(net17867),
    .A2(net18763),
    .Z(_14443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23419_ (.A1(net21202),
    .A2(_14336_),
    .ZN(_14444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23420_ (.A1(_14334_),
    .A2(_07874_),
    .A3(_14335_),
    .ZN(_14445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23421_ (.A1(_14445_),
    .A2(_14444_),
    .ZN(_15834_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23422_ (.A1(net19228),
    .A2(_14379_),
    .ZN(_14446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23423_ (.A1(_14443_),
    .A2(net18749),
    .ZN(_14447_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23424_ (.A1(net21460),
    .A2(_11339_),
    .ZN(_14448_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23425_ (.A1(net21406),
    .A2(net21351),
    .ZN(_14449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23426_ (.I(_14449_),
    .ZN(_14450_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23427_ (.A1(_14448_),
    .A2(_14450_),
    .Z(_14451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23428_ (.A1(_14448_),
    .A2(_14450_),
    .ZN(_14452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23429_ (.A1(_14451_),
    .A2(_14452_),
    .A3(net21067),
    .ZN(_14453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23430_ (.A1(net21495),
    .A2(\text_in_r[85] ),
    .ZN(_14454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23431_ (.A1(_14453_),
    .A2(_14454_),
    .ZN(_14455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23432_ (.A1(_14455_),
    .A2(net21197),
    .ZN(_14456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23433_ (.A1(_14453_),
    .A2(_07893_),
    .A3(_14454_),
    .ZN(_14457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23434_ (.A1(_14456_),
    .A2(_14457_),
    .ZN(_14458_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _23435_ (.I(_14458_),
    .ZN(_14459_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19492 (.I(net19487),
    .Z(net19492));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23437_ (.A1(_14437_),
    .A2(_14447_),
    .B(_14459_),
    .ZN(_14461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23438_ (.I(_15835_[0]),
    .ZN(_14462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23439_ (.A1(net19780),
    .A2(_14462_),
    .ZN(_14463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23440_ (.I(_14463_),
    .ZN(_14464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23441_ (.A1(_14464_),
    .A2(net18750),
    .ZN(_14465_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17236 (.I(_05727_),
    .Z(net17236));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23443_ (.A1(_14465_),
    .A2(net18764),
    .Z(_14467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23444_ (.A1(_14414_),
    .A2(_14438_),
    .ZN(_14468_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _23445_ (.I(_14468_),
    .ZN(_14469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23446_ (.A1(net19790),
    .A2(net18405),
    .ZN(_14470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23447_ (.A1(net17314),
    .A2(net18234),
    .ZN(_14471_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _23448_ (.I(_15843_[0]),
    .ZN(_14472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23449_ (.A1(net19793),
    .A2(_14472_),
    .Z(_14473_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17238 (.I(_04273_),
    .Z(net17238));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23451_ (.A1(_14473_),
    .A2(net18760),
    .ZN(_14475_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23452_ (.A1(_14467_),
    .A2(_14471_),
    .A3(_14475_),
    .ZN(_14476_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23453_ (.A1(net21405),
    .A2(net21350),
    .ZN(_14477_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23454_ (.I(\sa01_sr[6] ),
    .ZN(_14478_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23455_ (.A1(_14478_),
    .A2(_11382_),
    .Z(_14479_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _23456_ (.A1(_14477_),
    .A2(_14479_),
    .ZN(_14480_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23457_ (.A1(net21496),
    .A2(\text_in_r[86] ),
    .Z(_14481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23458_ (.A1(_14480_),
    .A2(net21071),
    .B(_14481_),
    .ZN(_14482_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23459_ (.A1(net21196),
    .A2(_14482_),
    .Z(_14483_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19491 (.I(net19487),
    .Z(net19491));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _23461_ (.I(_14483_),
    .ZN(_14485_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17235 (.I(_06173_),
    .Z(net17235));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23463_ (.A1(_14461_),
    .A2(_14476_),
    .B(net20242),
    .ZN(_14487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23464_ (.A1(_14384_),
    .A2(net19796),
    .ZN(_14488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23465_ (.A1(net19221),
    .A2(net18750),
    .ZN(_14489_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _23466_ (.I(_14489_),
    .ZN(_14490_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23467_ (.A1(net19225),
    .A2(net19787),
    .ZN(_14491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23468_ (.A1(_14490_),
    .A2(_14491_),
    .ZN(_14492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23469_ (.A1(net19230),
    .A2(net19787),
    .ZN(_14493_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17237 (.I(_05598_),
    .Z(net17237));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23471_ (.A1(_14379_),
    .A2(net19795),
    .ZN(_14495_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23472_ (.A1(_14493_),
    .A2(net18782),
    .A3(net19220),
    .ZN(_14496_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17234 (.I(_06315_),
    .Z(net17234));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23474_ (.A1(_14492_),
    .A2(_14496_),
    .A3(net18240),
    .ZN(_14498_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23475_ (.A1(net19230),
    .A2(net19797),
    .A3(net19793),
    .ZN(_14499_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23476_ (.A1(_14499_),
    .A2(_14443_),
    .ZN(_14500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23477_ (.A1(net19791),
    .A2(net18235),
    .ZN(_14501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23478_ (.A1(net19782),
    .A2(_14472_),
    .ZN(_14502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23479_ (.A1(_14501_),
    .A2(_14502_),
    .ZN(_14503_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17232 (.I(_11613_),
    .Z(net17232));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23481_ (.A1(_14503_),
    .A2(net18779),
    .ZN(_14505_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17233 (.I(_06514_),
    .Z(net17233));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23483_ (.A1(_14500_),
    .A2(_14505_),
    .A3(net18770),
    .ZN(_14507_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17244 (.I(_03883_),
    .Z(net17244));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17242 (.I(_04086_),
    .Z(net17242));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23486_ (.A1(_14498_),
    .A2(_14507_),
    .A3(net19779),
    .ZN(_14510_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23487_ (.A1(net21459),
    .A2(net21404),
    .Z(_14511_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23488_ (.A1(net21349),
    .A2(_14511_),
    .Z(_14512_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _23489_ (.A1(net443),
    .A2(net21285),
    .A3(_14512_),
    .Z(_14513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _23490_ (.I0(_14513_),
    .I1(\text_in_r[87] ),
    .S(net21493),
    .Z(_14514_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _23491_ (.A1(_07904_),
    .A2(_14514_),
    .Z(_14515_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17252 (.I(_03420_),
    .Z(net17252));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23493_ (.I(_14515_),
    .ZN(_14517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23494_ (.A1(_14487_),
    .A2(_14510_),
    .B(_14517_),
    .ZN(_14518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23495_ (.A1(net19225),
    .A2(net19780),
    .ZN(_14519_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _23496_ (.I(_14519_),
    .ZN(_14520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23497_ (.A1(_14379_),
    .A2(net19787),
    .ZN(_14521_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17230 (.I(_12266_),
    .Z(net17230));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _23499_ (.A1(_14521_),
    .A2(net19225),
    .B(net18750),
    .ZN(_14523_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23500_ (.I(_15849_[0]),
    .ZN(_14524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23501_ (.A1(net19780),
    .A2(_14524_),
    .ZN(_14525_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19462 (.I(_06762_),
    .Z(net19462));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23503_ (.A1(net19217),
    .A2(net17860),
    .A3(net18788),
    .ZN(_14527_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17228 (.I(_12355_),
    .Z(net17228));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23505_ (.A1(net18231),
    .A2(_14523_),
    .B(_14527_),
    .C(net18238),
    .ZN(_14529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23506_ (.I(_14488_),
    .ZN(_14530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23507_ (.A1(_14530_),
    .A2(net19230),
    .ZN(_14531_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17227 (.I(_12385_),
    .Z(net17227));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23509_ (.A1(_14531_),
    .A2(net18786),
    .A3(net19217),
    .ZN(_14533_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23510_ (.I(_14446_),
    .ZN(_14534_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _23511_ (.I(_15837_[0]),
    .ZN(_14535_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _23512_ (.A1(net19792),
    .A2(_14535_),
    .ZN(_14536_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17255 (.I(_03338_),
    .Z(net17255));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23514_ (.A1(_14534_),
    .A2(net17858),
    .B(net18761),
    .ZN(_14538_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23515_ (.A1(_14533_),
    .A2(_14538_),
    .A3(net18768),
    .ZN(_14539_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17229 (.I(_12296_),
    .Z(net17229));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23517_ (.A1(_14529_),
    .A2(_14539_),
    .A3(net20019),
    .ZN(_14541_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _23518_ (.A1(net19217),
    .A2(net19226),
    .ZN(_14542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23519_ (.I(_15840_[0]),
    .ZN(_14543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23520_ (.A1(net19783),
    .A2(net18226),
    .ZN(_14544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23521_ (.A1(_14544_),
    .A2(net18782),
    .ZN(_14545_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23522_ (.A1(_14542_),
    .A2(_14545_),
    .ZN(_14546_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19456 (.I(net19455),
    .Z(net19456));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23524_ (.A1(_14521_),
    .A2(net18750),
    .ZN(_14548_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _23525_ (.I(_14548_),
    .ZN(_14549_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _23526_ (.A1(_14546_),
    .A2(net18239),
    .A3(_14549_),
    .Z(_14550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23527_ (.A1(net19793),
    .A2(_14524_),
    .ZN(_14551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23528_ (.A1(_14551_),
    .A2(net18783),
    .ZN(_14552_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _23529_ (.I(_14552_),
    .ZN(_14553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23530_ (.A1(_14553_),
    .A2(net17867),
    .ZN(_14554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23531_ (.A1(net19784),
    .A2(net19787),
    .ZN(_14555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23532_ (.A1(net18746),
    .A2(net18750),
    .A3(net19215),
    .ZN(_14556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23533_ (.A1(_14554_),
    .A2(_14556_),
    .A3(net18239),
    .ZN(_14557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23534_ (.A1(_14550_),
    .A2(_14459_),
    .A3(_14557_),
    .ZN(_14558_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23535_ (.A1(_14541_),
    .A2(_14558_),
    .A3(net20242),
    .ZN(_14559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23536_ (.A1(_14518_),
    .A2(_14559_),
    .ZN(_14560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23537_ (.A1(net19230),
    .A2(net19784),
    .ZN(_14561_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23538_ (.A1(_14561_),
    .A2(net18750),
    .Z(_14562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23539_ (.A1(net20244),
    .A2(net20021),
    .A3(net18403),
    .ZN(_14563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23540_ (.A1(_14562_),
    .A2(net18224),
    .ZN(_14564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23541_ (.A1(net19794),
    .A2(_15843_[0]),
    .ZN(_14565_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23542_ (.A1(net18222),
    .A2(net18771),
    .Z(_14566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23543_ (.A1(_14566_),
    .A2(net19215),
    .ZN(_14567_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17239 (.I(_04267_),
    .Z(net17239));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23545_ (.A1(_14564_),
    .A2(_14567_),
    .B(net18240),
    .ZN(_14569_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23546_ (.I(_14536_),
    .ZN(_14570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23547_ (.A1(_14570_),
    .A2(_14501_),
    .ZN(_14571_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17219 (.I(_14858_),
    .Z(net17219));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23549_ (.A1(_14571_),
    .A2(net18760),
    .ZN(_14573_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19455 (.I(_16169_[0]),
    .Z(net19455));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23551_ (.A1(_14573_),
    .A2(_14545_),
    .B(net18765),
    .ZN(_14575_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23552_ (.A1(_14569_),
    .A2(_14575_),
    .B(net20242),
    .ZN(_14576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23553_ (.A1(_14536_),
    .A2(net18785),
    .ZN(_14577_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23554_ (.A1(_14577_),
    .A2(net18245),
    .Z(_14578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23555_ (.A1(_14565_),
    .A2(net18750),
    .ZN(_14579_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23556_ (.I(_14579_),
    .ZN(_14580_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23557_ (.A1(_14379_),
    .A2(net19795),
    .ZN(_14581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23558_ (.A1(_14581_),
    .A2(net19229),
    .ZN(_14582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23559_ (.A1(_14580_),
    .A2(net18741),
    .ZN(_14583_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19461 (.I(net19460),
    .Z(net19461));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23561_ (.A1(_14578_),
    .A2(_14583_),
    .B(_14485_),
    .ZN(_14585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23562_ (.I(_15845_[0]),
    .ZN(_14586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23563_ (.A1(_14379_),
    .A2(_14586_),
    .ZN(_14587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23564_ (.A1(_14587_),
    .A2(_14414_),
    .ZN(_14588_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23565_ (.I(_14588_),
    .ZN(_14589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23566_ (.A1(net17312),
    .A2(net18741),
    .ZN(_14590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23567_ (.A1(net17858),
    .A2(net18760),
    .ZN(_14591_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23568_ (.A1(_14590_),
    .A2(net18765),
    .A3(_14591_),
    .ZN(_14592_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17215 (.I(_15431_),
    .Z(net17215));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23570_ (.A1(_14585_),
    .A2(_14592_),
    .B(net20019),
    .ZN(_14594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23571_ (.A1(_14576_),
    .A2(_14594_),
    .ZN(_14595_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23572_ (.A1(net19780),
    .A2(net18226),
    .ZN(_14596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23573_ (.A1(net18756),
    .A2(net17849),
    .B(net18236),
    .ZN(_14597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23574_ (.A1(_14533_),
    .A2(_14597_),
    .ZN(_14598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23575_ (.A1(net19792),
    .A2(net18401),
    .ZN(_14599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23576_ (.A1(net19780),
    .A2(net18400),
    .ZN(_14600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23577_ (.A1(_14599_),
    .A2(_14600_),
    .ZN(_14601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23578_ (.A1(_14601_),
    .A2(net18752),
    .ZN(_14602_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23579_ (.A1(_14602_),
    .A2(net17526),
    .A3(net18245),
    .ZN(_14603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23580_ (.A1(_14598_),
    .A2(_14603_),
    .A3(net20243),
    .ZN(_14604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23581_ (.A1(net19219),
    .A2(net17864),
    .ZN(_14605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23582_ (.A1(_14605_),
    .A2(net18774),
    .B(net18249),
    .ZN(_14606_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17220 (.I(_13162_),
    .Z(net17220));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23584_ (.A1(net19792),
    .A2(net18226),
    .ZN(_14608_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23585_ (.A1(_14582_),
    .A2(net18753),
    .A3(_14608_),
    .ZN(_14609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23586_ (.A1(net19792),
    .A2(net18402),
    .ZN(_14610_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23587_ (.I(_14610_),
    .ZN(_14611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23588_ (.A1(_14611_),
    .A2(net18750),
    .Z(_14612_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _23589_ (.I(_14612_),
    .ZN(_14613_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23590_ (.A1(_14606_),
    .A2(_14609_),
    .A3(_14613_),
    .ZN(_14614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23591_ (.A1(net18782),
    .A2(_15856_[0]),
    .ZN(_14615_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23592_ (.I(_14563_),
    .ZN(_14616_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17216 (.I(_15299_),
    .Z(net17216));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23594_ (.A1(_14616_),
    .A2(net18761),
    .B(net18764),
    .ZN(_14618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23595_ (.A1(_14615_),
    .A2(_14618_),
    .B(_14485_),
    .ZN(_14619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23596_ (.A1(_14614_),
    .A2(_14619_),
    .ZN(_14620_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23597_ (.A1(_14604_),
    .A2(_14620_),
    .A3(net20019),
    .ZN(_14621_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23598_ (.A1(_14595_),
    .A2(_14621_),
    .A3(net20431),
    .ZN(_14622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23599_ (.A1(_14560_),
    .A2(_14622_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23600_ (.A1(_14552_),
    .A2(_14520_),
    .B(net18245),
    .ZN(_14623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23601_ (.A1(_14519_),
    .A2(_14555_),
    .ZN(_14624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23602_ (.A1(_14624_),
    .A2(net18758),
    .Z(_14625_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23603_ (.A1(_14623_),
    .A2(_14625_),
    .ZN(_14626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23604_ (.A1(_14446_),
    .A2(net19216),
    .A3(net17866),
    .ZN(_14627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23605_ (.A1(net19783),
    .A2(net18401),
    .ZN(_14628_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23606_ (.A1(_14628_),
    .A2(net18776),
    .B(net18764),
    .ZN(_14629_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23607_ (.A1(_14627_),
    .A2(net18773),
    .B(_14629_),
    .ZN(_14630_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23608_ (.A1(_14626_),
    .A2(_14630_),
    .B(_14459_),
    .ZN(_14631_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23609_ (.A1(net19220),
    .A2(net17864),
    .A3(net18752),
    .ZN(_14632_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23610_ (.A1(_14599_),
    .A2(net17866),
    .A3(net18771),
    .ZN(_14633_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20436 (.I(net20433),
    .Z(net20436));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23612_ (.A1(_14632_),
    .A2(_14633_),
    .B(net18764),
    .ZN(_14635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23613_ (.A1(_14563_),
    .A2(net18750),
    .ZN(_14636_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23614_ (.A1(_14636_),
    .A2(net19214),
    .B(net18764),
    .ZN(_14637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23615_ (.A1(net19230),
    .A2(net19797),
    .ZN(_14638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23616_ (.A1(_14638_),
    .A2(_14555_),
    .B(net18759),
    .ZN(_14639_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23617_ (.A1(_14637_),
    .A2(_14639_),
    .ZN(_14640_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23618_ (.A1(_14635_),
    .A2(_14640_),
    .B(net20017),
    .ZN(_14641_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23619_ (.A1(_14631_),
    .A2(net20240),
    .A3(_14641_),
    .ZN(_14642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23620_ (.A1(net19780),
    .A2(net18399),
    .ZN(_14643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23621_ (.A1(_14643_),
    .A2(_14563_),
    .ZN(_14644_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23622_ (.A1(_14644_),
    .A2(net18784),
    .B(_14435_),
    .ZN(_14645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23623_ (.A1(_14645_),
    .A2(_14609_),
    .ZN(_14646_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23624_ (.A1(_14596_),
    .A2(net18750),
    .B(net18764),
    .ZN(_14647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23625_ (.A1(net19230),
    .A2(net19793),
    .ZN(_14648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23626_ (.A1(_14648_),
    .A2(net18786),
    .ZN(_14649_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23627_ (.A1(_14647_),
    .A2(net18744),
    .A3(_14649_),
    .ZN(_14650_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23628_ (.A1(_14646_),
    .A2(_14650_),
    .A3(net20016),
    .ZN(_14651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23629_ (.A1(_14469_),
    .A2(net19216),
    .ZN(_14652_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23630_ (.A1(net19220),
    .A2(_14544_),
    .A3(net18758),
    .ZN(_14653_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19849 (.I(net19840),
    .Z(net19849));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23632_ (.A1(_14652_),
    .A2(_14653_),
    .A3(net18246),
    .ZN(_14655_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23633_ (.A1(net18750),
    .A2(net19780),
    .ZN(_14656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23634_ (.A1(_14656_),
    .A2(_14493_),
    .B(net18247),
    .ZN(_14657_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23635_ (.A1(_14561_),
    .A2(_14491_),
    .A3(net18750),
    .ZN(_14658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23636_ (.A1(_14657_),
    .A2(_14658_),
    .ZN(_14659_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23637_ (.A1(_14655_),
    .A2(_14659_),
    .A3(_14459_),
    .ZN(_14660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23638_ (.A1(_14660_),
    .A2(_14651_),
    .ZN(_14661_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20629 (.I(_04579_),
    .Z(net20629));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23640_ (.A1(_14661_),
    .A2(net20435),
    .ZN(_14663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23641_ (.A1(_14663_),
    .A2(_14642_),
    .ZN(_14664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23642_ (.A1(_14664_),
    .A2(net20432),
    .ZN(_14665_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23643_ (.A1(_14495_),
    .A2(net18781),
    .ZN(_14666_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23644_ (.A1(_14563_),
    .A2(net18750),
    .ZN(_14667_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23645_ (.A1(_14666_),
    .A2(_14667_),
    .ZN(_14668_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23646_ (.A1(net17857),
    .A2(net18750),
    .B(net18764),
    .ZN(_14669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23647_ (.A1(_14464_),
    .A2(net18771),
    .ZN(_14670_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23648_ (.A1(_14668_),
    .A2(_14669_),
    .A3(_14670_),
    .ZN(_14671_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _23649_ (.A1(_14446_),
    .A2(net18771),
    .A3(_14544_),
    .ZN(_14672_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23650_ (.A1(net19223),
    .A2(_14470_),
    .A3(net18751),
    .ZN(_14673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23651_ (.A1(_14672_),
    .A2(_14673_),
    .A3(net18770),
    .ZN(_14674_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23652_ (.A1(_14671_),
    .A2(_14674_),
    .A3(_14459_),
    .ZN(_14675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23653_ (.A1(net18230),
    .A2(_14549_),
    .ZN(_14676_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23654_ (.A1(_14468_),
    .A2(net18764),
    .Z(_14677_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23655_ (.A1(_14676_),
    .A2(_14677_),
    .B(_14459_),
    .ZN(_14678_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23656_ (.A1(_14525_),
    .A2(net18750),
    .Z(_14679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23657_ (.A1(net19792),
    .A2(net18227),
    .ZN(_14680_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23658_ (.A1(_14679_),
    .A2(net17844),
    .B(net18766),
    .ZN(_14681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23659_ (.A1(_14627_),
    .A2(net18790),
    .ZN(_14682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23660_ (.A1(_14681_),
    .A2(_14682_),
    .ZN(_14683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23661_ (.A1(_14678_),
    .A2(_14683_),
    .ZN(_14684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23662_ (.A1(_14675_),
    .A2(_14684_),
    .B(net20435),
    .ZN(_14685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23663_ (.A1(_14490_),
    .A2(net18738),
    .ZN(_14686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23664_ (.A1(_14686_),
    .A2(_14672_),
    .ZN(_14687_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23665_ (.A1(_14687_),
    .A2(net20017),
    .B(net18770),
    .ZN(_14688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23666_ (.A1(_14495_),
    .A2(net19229),
    .ZN(_14689_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20737 (.I(net20721),
    .Z(net20737));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23668_ (.A1(_14689_),
    .A2(net19214),
    .B(net18777),
    .ZN(_14691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23669_ (.A1(net19215),
    .A2(_14470_),
    .A3(net18751),
    .ZN(_14692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23670_ (.A1(_14691_),
    .A2(_14692_),
    .ZN(_14693_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23671_ (.A1(_14693_),
    .A2(_14459_),
    .ZN(_14694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23672_ (.I(_15859_[0]),
    .ZN(_14695_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23673_ (.A1(net18771),
    .A2(_14695_),
    .Z(_14696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23674_ (.A1(_14696_),
    .A2(net20018),
    .B(net18248),
    .ZN(_14697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23675_ (.A1(_14531_),
    .A2(_14580_),
    .ZN(_14698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23676_ (.A1(_14697_),
    .A2(_14698_),
    .ZN(_14699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23677_ (.A1(_14699_),
    .A2(net20433),
    .ZN(_14700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23678_ (.A1(_14688_),
    .A2(_14694_),
    .B(_14700_),
    .ZN(_14701_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23679_ (.A1(_14685_),
    .A2(_14701_),
    .B(net20632),
    .ZN(_14702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23680_ (.A1(_14665_),
    .A2(_14702_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23681_ (.A1(_14525_),
    .A2(net18786),
    .Z(_14703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23682_ (.A1(_14703_),
    .A2(_14499_),
    .ZN(_14704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23683_ (.A1(_14704_),
    .A2(_14523_),
    .ZN(_14705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23684_ (.A1(_14705_),
    .A2(net18764),
    .ZN(_14706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23685_ (.A1(net19780),
    .A2(net18404),
    .ZN(_14707_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23686_ (.A1(net18748),
    .A2(net18758),
    .A3(_14707_),
    .ZN(_14708_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23687_ (.A1(net19223),
    .A2(net18219),
    .A3(net18775),
    .ZN(_14709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23688_ (.A1(_14708_),
    .A2(_14709_),
    .A3(net18248),
    .ZN(_14710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23689_ (.A1(_14706_),
    .A2(_14459_),
    .A3(_14710_),
    .ZN(_14711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23690_ (.A1(_14689_),
    .A2(net18778),
    .ZN(_14712_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23691_ (.A1(_14544_),
    .A2(net17852),
    .A3(net18750),
    .ZN(_14713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23692_ (.A1(_14712_),
    .A2(_14713_),
    .ZN(_14714_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23693_ (.A1(_14714_),
    .A2(net18242),
    .B(_14459_),
    .ZN(_14715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23694_ (.A1(_14582_),
    .A2(_14608_),
    .ZN(_14716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23695_ (.A1(_14716_),
    .A2(net18774),
    .ZN(_14717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23696_ (.A1(_14717_),
    .A2(_14564_),
    .A3(net18770),
    .ZN(_14718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23697_ (.A1(_14715_),
    .A2(_14718_),
    .ZN(_14719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23698_ (.A1(_14711_),
    .A2(_14719_),
    .ZN(_14720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23699_ (.A1(_14720_),
    .A2(net20434),
    .ZN(_14721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23700_ (.A1(net19793),
    .A2(net18399),
    .ZN(_14722_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23701_ (.I(_14722_),
    .ZN(_14723_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23702_ (.A1(net18232),
    .A2(_14723_),
    .B(net18247),
    .ZN(_14724_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23703_ (.A1(net18749),
    .A2(net18772),
    .A3(net18221),
    .Z(_14725_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23704_ (.A1(_14724_),
    .A2(_14725_),
    .ZN(_14726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23705_ (.A1(_14563_),
    .A2(net18771),
    .Z(_14727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23706_ (.A1(_14727_),
    .A2(net17866),
    .ZN(_14728_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23707_ (.A1(net19215),
    .A2(net17850),
    .A3(net18763),
    .ZN(_14729_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23708_ (.A1(_14728_),
    .A2(_14729_),
    .B(net18240),
    .ZN(_14730_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23709_ (.A1(_14726_),
    .A2(_14730_),
    .B(net19779),
    .ZN(_14731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23710_ (.A1(net18744),
    .A2(net18773),
    .A3(net17848),
    .ZN(_14732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23711_ (.A1(_14732_),
    .A2(_14602_),
    .A3(net18764),
    .ZN(_14733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23712_ (.A1(net19222),
    .A2(net18786),
    .ZN(_14734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23713_ (.A1(_14722_),
    .A2(net18750),
    .ZN(_14735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23714_ (.A1(_14734_),
    .A2(net17849),
    .B(_14735_),
    .ZN(_14736_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23715_ (.I(_14600_),
    .ZN(_14737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23716_ (.A1(_14737_),
    .A2(net18750),
    .ZN(_14738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23717_ (.A1(_14738_),
    .A2(net18246),
    .Z(_14739_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23718_ (.A1(_14736_),
    .A2(_14739_),
    .ZN(_14740_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23719_ (.A1(_14733_),
    .A2(_14740_),
    .A3(net20017),
    .ZN(_14741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23720_ (.A1(_14731_),
    .A2(_14741_),
    .A3(net20239),
    .ZN(_14742_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23721_ (.A1(_14721_),
    .A2(_14742_),
    .A3(net20632),
    .ZN(_14743_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23722_ (.A1(_14446_),
    .A2(net18771),
    .Z(_14744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23723_ (.A1(_14744_),
    .A2(net19215),
    .ZN(_14745_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20696 (.I(_07706_),
    .Z(net20696));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23725_ (.A1(_14564_),
    .A2(_14745_),
    .B(net20017),
    .ZN(_14747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23726_ (.A1(_14727_),
    .A2(net17861),
    .B(_14459_),
    .ZN(_14748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23727_ (.A1(net18225),
    .A2(_14501_),
    .ZN(_14749_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23728_ (.A1(_14748_),
    .A2(_14749_),
    .Z(_14750_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23729_ (.A1(_14747_),
    .A2(_14750_),
    .B(net18244),
    .ZN(_14751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23730_ (.A1(_15856_[0]),
    .A2(net18758),
    .B(_14458_),
    .ZN(_14752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23731_ (.A1(_14387_),
    .A2(net18771),
    .Z(_14753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23732_ (.A1(_14753_),
    .A2(_14582_),
    .ZN(_14754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23733_ (.A1(_14752_),
    .A2(_14754_),
    .B(_14435_),
    .ZN(_14755_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23734_ (.A1(_14561_),
    .A2(_14491_),
    .A3(net18771),
    .ZN(_14756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23735_ (.A1(net18759),
    .A2(net18213),
    .ZN(_14757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23736_ (.A1(_14756_),
    .A2(net20018),
    .A3(_14757_),
    .ZN(_14758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23737_ (.A1(_14755_),
    .A2(_14758_),
    .B(net20433),
    .ZN(_14759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23738_ (.A1(_14751_),
    .A2(_14759_),
    .ZN(_14760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23739_ (.A1(_14656_),
    .A2(net18739),
    .ZN(_14761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23740_ (.A1(_14761_),
    .A2(net18246),
    .Z(_14762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23741_ (.A1(net18786),
    .A2(net19780),
    .ZN(_14763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23742_ (.A1(_14535_),
    .A2(_14543_),
    .Z(_14764_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23743_ (.A1(_14763_),
    .A2(_14764_),
    .Z(_14765_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23744_ (.A1(_14762_),
    .A2(_14698_),
    .A3(_14765_),
    .ZN(_14766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23745_ (.A1(net17315),
    .A2(net17848),
    .ZN(_14767_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23746_ (.A1(_14767_),
    .A2(_14467_),
    .B(net20017),
    .ZN(_14768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23747_ (.A1(_14768_),
    .A2(_14766_),
    .ZN(_14769_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _23748_ (.A1(net18750),
    .A2(_15854_[0]),
    .Z(_14770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23749_ (.A1(_14523_),
    .A2(_14770_),
    .ZN(_14771_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23750_ (.A1(_14771_),
    .A2(net18240),
    .Z(_14772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23751_ (.A1(_15863_[0]),
    .A2(net18751),
    .B(net18770),
    .ZN(_14773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23752_ (.A1(_14773_),
    .A2(_14712_),
    .B(_14459_),
    .ZN(_14774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23753_ (.A1(_14772_),
    .A2(_14774_),
    .ZN(_14775_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23754_ (.A1(_14769_),
    .A2(net20434),
    .A3(_14775_),
    .ZN(_14776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23755_ (.A1(_14776_),
    .A2(_14760_),
    .A3(net20432),
    .ZN(_14777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23756_ (.A1(_14743_),
    .A2(_14777_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23757_ (.A1(net18218),
    .A2(_14636_),
    .Z(_14778_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23758_ (.A1(net19219),
    .A2(_14502_),
    .Z(_14779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23759_ (.A1(net18211),
    .A2(_14779_),
    .ZN(_14780_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23760_ (.A1(_14778_),
    .A2(_14780_),
    .A3(net18770),
    .ZN(_14781_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23761_ (.I(_14438_),
    .ZN(_14782_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _23762_ (.A1(_14473_),
    .A2(net18780),
    .A3(_14782_),
    .Z(_14783_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23763_ (.A1(_14783_),
    .A2(net18241),
    .A3(_14496_),
    .ZN(_14784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23764_ (.A1(_14781_),
    .A2(_14784_),
    .ZN(_14785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23765_ (.A1(_14785_),
    .A2(net19779),
    .ZN(_14786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23766_ (.A1(_14493_),
    .A2(net19222),
    .ZN(_14787_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23767_ (.A1(_14787_),
    .A2(net18764),
    .Z(_14788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23768_ (.A1(_14788_),
    .A2(_14763_),
    .B(_14459_),
    .ZN(_14789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23769_ (.A1(_14587_),
    .A2(net18750),
    .Z(_14790_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23770_ (.A1(_14790_),
    .A2(_14707_),
    .Z(_14791_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23771_ (.A1(_14623_),
    .A2(_14791_),
    .Z(_14792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23772_ (.A1(_14789_),
    .A2(_14792_),
    .B(net20435),
    .ZN(_14793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23773_ (.A1(_14786_),
    .A2(_14793_),
    .ZN(_14794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23774_ (.A1(_14779_),
    .A2(net18751),
    .ZN(_14795_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23775_ (.A1(net17868),
    .A2(net17865),
    .A3(net18778),
    .ZN(_14796_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23776_ (.A1(_14795_),
    .A2(_14459_),
    .A3(_14796_),
    .ZN(_14797_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23777_ (.A1(_14686_),
    .A2(net20017),
    .A3(_14416_),
    .ZN(_14798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23778_ (.A1(_14797_),
    .A2(_14798_),
    .ZN(_14799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23779_ (.A1(_14799_),
    .A2(net18243),
    .ZN(_14800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23780_ (.A1(net17863),
    .A2(net18747),
    .ZN(_14801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23781_ (.A1(net17315),
    .A2(net18749),
    .ZN(_14802_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23782_ (.A1(_14801_),
    .A2(_14802_),
    .A3(net20017),
    .ZN(_14803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23783_ (.A1(_14703_),
    .A2(net17848),
    .ZN(_14804_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23784_ (.A1(_14804_),
    .A2(_14708_),
    .A3(_14459_),
    .ZN(_14805_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23785_ (.A1(_14803_),
    .A2(_14805_),
    .A3(net18770),
    .ZN(_14806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23786_ (.A1(_14800_),
    .A2(_14806_),
    .A3(net20434),
    .ZN(_14807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23787_ (.A1(_14794_),
    .A2(_14807_),
    .A3(net20432),
    .ZN(_14808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23788_ (.A1(net17843),
    .A2(net18772),
    .B(_14458_),
    .ZN(_14809_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23789_ (.A1(_14809_),
    .A2(_14729_),
    .B(net18240),
    .ZN(_14810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23790_ (.A1(_14549_),
    .A2(net17867),
    .ZN(_14811_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23791_ (.A1(net19780),
    .A2(_14764_),
    .ZN(_14812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23792_ (.A1(_14812_),
    .A2(net18785),
    .Z(_14813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23793_ (.A1(net17311),
    .A2(net17854),
    .ZN(_14814_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23794_ (.A1(_14811_),
    .A2(_14814_),
    .A3(net20016),
    .ZN(_14815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23795_ (.A1(_14810_),
    .A2(_14815_),
    .B(net20242),
    .ZN(_14816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23796_ (.A1(net18763),
    .A2(_14782_),
    .ZN(_14817_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23797_ (.I(_14817_),
    .ZN(_14818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _23798_ (.A1(_14818_),
    .A2(_14459_),
    .B1(net18772),
    .B2(net17857),
    .ZN(_14819_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _23799_ (.I(_14561_),
    .ZN(_14820_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23800_ (.A1(_14820_),
    .A2(_14579_),
    .B(_14416_),
    .ZN(_14821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23801_ (.A1(_14821_),
    .A2(_14458_),
    .ZN(_14822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23802_ (.A1(_14819_),
    .A2(_14822_),
    .ZN(_14823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23803_ (.A1(_14823_),
    .A2(net18239),
    .ZN(_14824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23804_ (.A1(_14816_),
    .A2(_14824_),
    .B(_14517_),
    .ZN(_14825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23805_ (.A1(_14813_),
    .A2(net17850),
    .ZN(_14826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23806_ (.A1(_14698_),
    .A2(_14826_),
    .B(net18246),
    .ZN(_14827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23807_ (.I(_14724_),
    .ZN(_14828_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23808_ (.A1(_14827_),
    .A2(_14828_),
    .B(net20016),
    .ZN(_14829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23809_ (.A1(_14606_),
    .A2(net18214),
    .ZN(_14830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23810_ (.A1(_14443_),
    .A2(net17854),
    .ZN(_14831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23811_ (.A1(net19216),
    .A2(_14600_),
    .ZN(_14832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _23812_ (.A1(_14832_),
    .A2(net18780),
    .ZN(_14833_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23813_ (.A1(_14831_),
    .A2(_14833_),
    .A3(net18240),
    .ZN(_14834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23814_ (.A1(_14830_),
    .A2(_14834_),
    .A3(net19779),
    .ZN(_14835_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23815_ (.A1(_14829_),
    .A2(_14835_),
    .A3(net20239),
    .ZN(_14836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23816_ (.A1(_14825_),
    .A2(_14836_),
    .ZN(_14837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23817_ (.A1(_14808_),
    .A2(_14837_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23818_ (.A1(net17859),
    .A2(net18769),
    .ZN(_14838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23819_ (.A1(net17856),
    .A2(net18762),
    .ZN(_14839_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23820_ (.A1(_14839_),
    .A2(net17847),
    .ZN(_14840_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23821_ (.A1(_14680_),
    .A2(net18754),
    .ZN(_14841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23822_ (.A1(_14841_),
    .A2(net18236),
    .Z(_14842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23823_ (.A1(_14499_),
    .A2(net18782),
    .ZN(_14843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23824_ (.A1(_14842_),
    .A2(_14843_),
    .B(net20019),
    .ZN(_14844_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23825_ (.A1(_14838_),
    .A2(_14840_),
    .B(_14844_),
    .ZN(_14845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23826_ (.A1(net17862),
    .A2(net17853),
    .ZN(_14846_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23827_ (.A1(net18215),
    .A2(net18236),
    .ZN(_14847_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23828_ (.A1(_14846_),
    .A2(_14847_),
    .B(_14459_),
    .ZN(_14848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23829_ (.A1(_14446_),
    .A2(_14463_),
    .ZN(_14849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23830_ (.A1(_14849_),
    .A2(net18753),
    .ZN(_14850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23831_ (.A1(_14850_),
    .A2(_14672_),
    .A3(net18246),
    .ZN(_14851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23832_ (.A1(_14848_),
    .A2(_14851_),
    .ZN(_14852_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23833_ (.A1(_14845_),
    .A2(_14852_),
    .A3(net20243),
    .ZN(_14853_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23834_ (.I(_15847_[0]),
    .ZN(_14854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23835_ (.A1(_14854_),
    .A2(net18758),
    .B(net18249),
    .ZN(_14855_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23836_ (.I(_14727_),
    .ZN(_14856_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23837_ (.A1(_14855_),
    .A2(_14856_),
    .B(net20017),
    .ZN(_14857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23838_ (.A1(_14589_),
    .A2(net18743),
    .ZN(_14858_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23839_ (.A1(_14493_),
    .A2(net19781),
    .A3(net18761),
    .ZN(_14859_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23840_ (.A1(net17219),
    .A2(net18210),
    .A3(net18236),
    .ZN(_14860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23841_ (.A1(_14857_),
    .A2(_14860_),
    .B(net20242),
    .ZN(_14861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23842_ (.A1(_14519_),
    .A2(_14638_),
    .ZN(_14862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23843_ (.A1(_14862_),
    .A2(net18754),
    .ZN(_14863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23844_ (.A1(net17312),
    .A2(net19222),
    .ZN(_14864_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23845_ (.A1(_14863_),
    .A2(_14864_),
    .A3(net18236),
    .ZN(_14865_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23846_ (.A1(_14573_),
    .A2(net18765),
    .A3(_14496_),
    .ZN(_14866_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23847_ (.A1(_14865_),
    .A2(_14866_),
    .A3(net20019),
    .ZN(_14867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23848_ (.A1(_14861_),
    .A2(_14867_),
    .ZN(_14868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23849_ (.A1(_14853_),
    .A2(net20632),
    .A3(_14868_),
    .ZN(_14869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23850_ (.A1(_14756_),
    .A2(net18764),
    .Z(_14870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23851_ (.A1(_14870_),
    .A2(_14686_),
    .ZN(_14871_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _23852_ (.A1(_14862_),
    .A2(net18787),
    .Z(_14872_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23853_ (.A1(net18744),
    .A2(net18784),
    .A3(net18234),
    .ZN(_14873_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23854_ (.A1(_14872_),
    .A2(_14873_),
    .A3(net18245),
    .ZN(_14874_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23855_ (.A1(_14871_),
    .A2(_14874_),
    .A3(net20019),
    .ZN(_14875_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _23856_ (.A1(_14649_),
    .A2(net19213),
    .Z(_14876_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23857_ (.A1(_14876_),
    .A2(net18770),
    .A3(_14692_),
    .ZN(_14877_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23858_ (.A1(_14570_),
    .A2(net18239),
    .Z(_14878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23859_ (.A1(_14878_),
    .A2(net17524),
    .B(net20019),
    .ZN(_14879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23860_ (.A1(_14877_),
    .A2(_14879_),
    .B(net20435),
    .ZN(_14880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23861_ (.A1(_14875_),
    .A2(_14880_),
    .ZN(_14881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23862_ (.A1(_14582_),
    .A2(net18790),
    .ZN(_14882_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23863_ (.A1(_14882_),
    .A2(net18228),
    .B(_14713_),
    .C(net18240),
    .ZN(_14883_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23864_ (.A1(_14670_),
    .A2(net18764),
    .Z(_14884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23865_ (.A1(net18215),
    .A2(net19230),
    .ZN(_14885_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23866_ (.A1(_14884_),
    .A2(_14609_),
    .A3(_14885_),
    .ZN(_14886_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23867_ (.A1(_14883_),
    .A2(_14886_),
    .A3(net20016),
    .ZN(_14887_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23868_ (.A1(_14667_),
    .A2(net17843),
    .ZN(_14888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23869_ (.A1(net17522),
    .A2(_14888_),
    .B(net20019),
    .ZN(_14889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23870_ (.A1(net17846),
    .A2(net18760),
    .ZN(_14890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23871_ (.A1(_14590_),
    .A2(net18764),
    .A3(_14890_),
    .ZN(_14891_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23872_ (.A1(_14889_),
    .A2(_14891_),
    .B(net20242),
    .ZN(_14892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23873_ (.A1(_14887_),
    .A2(_14892_),
    .ZN(_14893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23874_ (.A1(_14881_),
    .A2(_14893_),
    .A3(net20431),
    .ZN(_14894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23875_ (.A1(_14869_),
    .A2(_14894_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23876_ (.A1(_14531_),
    .A2(net18223),
    .ZN(_14895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23877_ (.A1(_14895_),
    .A2(net18789),
    .ZN(_14896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23878_ (.A1(net17855),
    .A2(net18740),
    .ZN(_14897_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23879_ (.A1(_14896_),
    .A2(net18236),
    .A3(_14897_),
    .Z(_14898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23880_ (.A1(net18789),
    .A2(net19226),
    .ZN(_14899_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _23881_ (.A1(_14863_),
    .A2(net18768),
    .A3(_14899_),
    .Z(_14900_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23882_ (.A1(_14898_),
    .A2(_14900_),
    .B(net19776),
    .ZN(_14901_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23883_ (.A1(_14841_),
    .A2(_14820_),
    .ZN(_14902_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23884_ (.A1(_14902_),
    .A2(net17845),
    .B(net18237),
    .ZN(_14903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23885_ (.A1(net17313),
    .A2(_14501_),
    .ZN(_14904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23886_ (.A1(_14904_),
    .A2(net18768),
    .A3(_14735_),
    .ZN(_14905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23887_ (.A1(_14905_),
    .A2(_14903_),
    .ZN(_14906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23888_ (.A1(_14906_),
    .A2(net20019),
    .B(net20243),
    .ZN(_14907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23889_ (.A1(_14907_),
    .A2(_14901_),
    .ZN(_14908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23890_ (.A1(_14553_),
    .A2(net17856),
    .ZN(_14909_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23891_ (.A1(_14538_),
    .A2(net18769),
    .A3(_14909_),
    .ZN(_14910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23892_ (.A1(net17521),
    .A2(net18741),
    .ZN(_14911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23893_ (.A1(net18787),
    .A2(net18401),
    .ZN(_14912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23894_ (.A1(_14578_),
    .A2(_14911_),
    .A3(_14912_),
    .ZN(_14913_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23895_ (.A1(_14910_),
    .A2(_14913_),
    .A3(net19775),
    .ZN(_14914_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23896_ (.A1(_14443_),
    .A2(net18239),
    .ZN(_14915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23897_ (.A1(_14915_),
    .A2(_14833_),
    .B(_14459_),
    .ZN(_14916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23898_ (.A1(net18215),
    .A2(net18745),
    .ZN(_14917_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23899_ (.A1(_14917_),
    .A2(net18237),
    .A3(_14839_),
    .ZN(_14918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23900_ (.A1(_14916_),
    .A2(_14918_),
    .B(net20436),
    .ZN(_14919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23901_ (.A1(_14914_),
    .A2(_14919_),
    .B(net20632),
    .ZN(_14920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23902_ (.A1(_14908_),
    .A2(_14920_),
    .ZN(_14921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23903_ (.A1(net18742),
    .A2(net18754),
    .ZN(_14922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23904_ (.I(net18209),
    .ZN(_14923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23905_ (.A1(net18229),
    .A2(net18755),
    .A3(net17853),
    .ZN(_14924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23906_ (.A1(_14473_),
    .A2(net18786),
    .B(net18768),
    .ZN(_14925_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23907_ (.A1(_14924_),
    .A2(_14925_),
    .B(_14459_),
    .ZN(_14926_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23908_ (.A1(_14598_),
    .A2(_14923_),
    .B(_14926_),
    .ZN(_14927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23909_ (.A1(net19797),
    .A2(net18786),
    .B(net18247),
    .ZN(_14928_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23910_ (.A1(_14928_),
    .A2(_14492_),
    .B(net20018),
    .ZN(_14929_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23911_ (.A1(_14542_),
    .A2(net17526),
    .Z(_14930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23912_ (.A1(_14790_),
    .A2(net18743),
    .ZN(_14931_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23913_ (.A1(_14930_),
    .A2(_14931_),
    .A3(net18236),
    .ZN(_14932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23914_ (.A1(_14929_),
    .A2(_14932_),
    .B(net20433),
    .ZN(_14933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23915_ (.A1(_14927_),
    .A2(_14933_),
    .ZN(_14934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23916_ (.A1(net17313),
    .A2(net18223),
    .ZN(_14935_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23917_ (.A1(net17853),
    .A2(net18212),
    .A3(net18755),
    .ZN(_14936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23918_ (.A1(_14935_),
    .A2(_14936_),
    .A3(net18236),
    .ZN(_14937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23919_ (.A1(net18233),
    .A2(net18789),
    .B(net18236),
    .ZN(_14938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23920_ (.A1(net18229),
    .A2(net18754),
    .ZN(_14939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23921_ (.A1(_14938_),
    .A2(_14939_),
    .ZN(_14940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23922_ (.A1(_14937_),
    .A2(_14940_),
    .A3(net20019),
    .ZN(_14941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23923_ (.A1(net17522),
    .A2(net17525),
    .B(net20019),
    .ZN(_14942_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23924_ (.A1(_14689_),
    .A2(net19213),
    .B(net18752),
    .ZN(_14943_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23925_ (.A1(net17311),
    .A2(net18245),
    .ZN(_14944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23926_ (.A1(_14943_),
    .A2(_14944_),
    .ZN(_14945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23927_ (.A1(_14942_),
    .A2(_14945_),
    .ZN(_14946_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23928_ (.A1(_14941_),
    .A2(net20436),
    .A3(_14946_),
    .ZN(_14947_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23929_ (.A1(_14934_),
    .A2(net20632),
    .A3(_14947_),
    .ZN(_14948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23930_ (.A1(_14921_),
    .A2(_14948_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23931_ (.A1(_14790_),
    .A2(net17860),
    .ZN(_14949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23932_ (.A1(_14949_),
    .A2(_14577_),
    .A3(_14761_),
    .ZN(_14950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23933_ (.A1(_14950_),
    .A2(net18766),
    .ZN(_14951_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _23934_ (.A1(net18775),
    .A2(_14599_),
    .A3(net18219),
    .A4(net18220),
    .ZN(_14952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23935_ (.A1(_14952_),
    .A2(_14618_),
    .A3(_14922_),
    .ZN(_14953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23936_ (.A1(_14951_),
    .A2(_14953_),
    .ZN(_14954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23937_ (.A1(_14954_),
    .A2(net20019),
    .ZN(_14955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23938_ (.A1(_14862_),
    .A2(net18787),
    .ZN(_14956_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23939_ (.A1(_15852_[0]),
    .A2(_15861_[0]),
    .Z(_14957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23940_ (.A1(net18757),
    .A2(_14957_),
    .B(net18236),
    .ZN(_14958_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23941_ (.A1(_14956_),
    .A2(_14958_),
    .B(net20019),
    .ZN(_14959_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23942_ (.A1(net18219),
    .A2(_14600_),
    .Z(_14960_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _23943_ (.A1(net18758),
    .A2(_14960_),
    .B(net17316),
    .C(net18249),
    .ZN(_14961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23944_ (.A1(_14959_),
    .A2(_14961_),
    .B(net20433),
    .ZN(_14962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23945_ (.A1(_14955_),
    .A2(_14962_),
    .ZN(_14963_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23946_ (.A1(_14771_),
    .A2(net18239),
    .A3(net17310),
    .ZN(_14964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23947_ (.A1(net18743),
    .A2(net18782),
    .ZN(_14965_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23948_ (.A1(_14965_),
    .A2(_14542_),
    .B(_14841_),
    .ZN(_14966_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23949_ (.I(_14707_),
    .ZN(_14967_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23950_ (.A1(_14967_),
    .A2(net18760),
    .B(net18236),
    .ZN(_14968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23951_ (.A1(_14966_),
    .A2(_14968_),
    .ZN(_14969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23952_ (.A1(_14964_),
    .A2(_14969_),
    .ZN(_14970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23953_ (.A1(_14970_),
    .A2(net19777),
    .ZN(_14971_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23954_ (.A1(net18741),
    .A2(net18782),
    .A3(net19220),
    .ZN(_14972_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23955_ (.A1(net17520),
    .A2(_14563_),
    .A3(net18761),
    .ZN(_14973_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23956_ (.A1(_14972_),
    .A2(net18767),
    .A3(_14973_),
    .ZN(_14974_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23957_ (.A1(net18742),
    .A2(net19226),
    .B(net18789),
    .ZN(_14975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23958_ (.A1(_14473_),
    .A2(net18760),
    .B(net18767),
    .ZN(_14976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23959_ (.A1(_14975_),
    .A2(_14976_),
    .B(_14459_),
    .ZN(_14977_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23960_ (.A1(_14974_),
    .A2(_14977_),
    .B(net20242),
    .ZN(_14978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23961_ (.A1(_14971_),
    .A2(_14978_),
    .ZN(_14979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23962_ (.A1(_14963_),
    .A2(net20431),
    .A3(_14979_),
    .ZN(_14980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23963_ (.A1(_14717_),
    .A2(net18768),
    .ZN(_14981_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _23964_ (.A1(net17523),
    .A2(_14520_),
    .B(net17851),
    .ZN(_14982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23965_ (.A1(_14982_),
    .A2(net18236),
    .ZN(_14983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23966_ (.A1(_14981_),
    .A2(_14983_),
    .ZN(_14984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23967_ (.A1(_14984_),
    .A2(net20019),
    .ZN(_14985_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _23968_ (.A1(net18754),
    .A2(_15853_[0]),
    .Z(_14986_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23969_ (.A1(_14931_),
    .A2(net18768),
    .A3(_14986_),
    .ZN(_14987_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23970_ (.I(_14666_),
    .ZN(_14988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _23971_ (.A1(_14988_),
    .A2(net18236),
    .Z(_14989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23972_ (.A1(_14553_),
    .A2(net18212),
    .ZN(_14990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23973_ (.A1(_14989_),
    .A2(_14990_),
    .ZN(_14991_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23974_ (.A1(_14987_),
    .A2(_14991_),
    .A3(net19775),
    .ZN(_14992_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23975_ (.A1(_14985_),
    .A2(_14992_),
    .A3(net20436),
    .ZN(_14993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23976_ (.A1(_14787_),
    .A2(net18788),
    .ZN(_14994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23977_ (.A1(net19218),
    .A2(net18217),
    .ZN(_14995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23978_ (.A1(_14995_),
    .A2(net18750),
    .ZN(_14996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23979_ (.A1(_14994_),
    .A2(_14996_),
    .A3(net18238),
    .ZN(_14997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23980_ (.A1(net18750),
    .A2(net19225),
    .ZN(_14998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23981_ (.A1(_14788_),
    .A2(net18208),
    .ZN(_14999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23982_ (.A1(_14997_),
    .A2(_14999_),
    .A3(net19778),
    .ZN(_15000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23983_ (.A1(_14556_),
    .A2(net18239),
    .A3(net18216),
    .ZN(_15001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23984_ (.A1(_14968_),
    .A2(_14833_),
    .ZN(_15002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23985_ (.A1(_15001_),
    .A2(_15002_),
    .A3(net20019),
    .ZN(_15003_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23986_ (.A1(_15000_),
    .A2(_15003_),
    .A3(net20242),
    .ZN(_15004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23987_ (.A1(_14993_),
    .A2(_15004_),
    .A3(net20632),
    .ZN(_15005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23988_ (.A1(_14980_),
    .A2(_15005_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23989_ (.A1(net18750),
    .A2(net19787),
    .Z(_15006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _23990_ (.I(_15006_),
    .ZN(_15007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23991_ (.A1(_14876_),
    .A2(_15007_),
    .ZN(_15008_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _23992_ (.A1(_15008_),
    .A2(net18240),
    .B(_14485_),
    .ZN(_15009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23993_ (.A1(_14820_),
    .A2(net18750),
    .ZN(_15010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23994_ (.A1(_14870_),
    .A2(_14872_),
    .A3(_15010_),
    .ZN(_15011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23995_ (.A1(_15009_),
    .A2(_15011_),
    .ZN(_15012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23996_ (.A1(_14446_),
    .A2(_14463_),
    .A3(_14521_),
    .ZN(_15013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _23997_ (.A1(_15013_),
    .A2(net18782),
    .ZN(_15014_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _23998_ (.A1(_15014_),
    .A2(_14989_),
    .A3(_14859_),
    .ZN(_15015_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _23999_ (.A1(_14679_),
    .A2(net18236),
    .ZN(_15016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24000_ (.A1(_15016_),
    .A2(_14858_),
    .B(net20433),
    .ZN(_15017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24001_ (.A1(_15015_),
    .A2(_15017_),
    .B(net20019),
    .ZN(_15018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24002_ (.A1(_15012_),
    .A2(_15018_),
    .ZN(_15019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24003_ (.A1(_14745_),
    .A2(_14949_),
    .B(net18240),
    .ZN(_15020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24004_ (.A1(_14644_),
    .A2(net18780),
    .ZN(_15021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24005_ (.A1(_14811_),
    .A2(_15021_),
    .B(net18764),
    .ZN(_15022_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24006_ (.A1(_15020_),
    .A2(_15022_),
    .B(net20241),
    .ZN(_15023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24007_ (.A1(_14627_),
    .A2(net18758),
    .ZN(_15024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24008_ (.A1(_15024_),
    .A2(net18240),
    .A3(_14882_),
    .ZN(_15025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24009_ (.A1(_14817_),
    .A2(net18764),
    .Z(_15026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24010_ (.A1(net18218),
    .A2(net18772),
    .ZN(_15027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24011_ (.A1(_15026_),
    .A2(_15027_),
    .B(_14485_),
    .ZN(_15028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24012_ (.A1(_15028_),
    .A2(_15025_),
    .B(_14459_),
    .ZN(_15029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24013_ (.A1(_15023_),
    .A2(_15029_),
    .ZN(_15030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24014_ (.A1(_15019_),
    .A2(_15030_),
    .A3(net20632),
    .ZN(_15031_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24015_ (.A1(_14854_),
    .A2(net18774),
    .B(net18249),
    .ZN(_15032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24016_ (.A1(_15032_),
    .A2(_14613_),
    .B(_14485_),
    .ZN(_15033_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24017_ (.A1(_14998_),
    .A2(_14435_),
    .Z(_15034_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24018_ (.A1(_14672_),
    .A2(net17842),
    .A3(_14922_),
    .ZN(_15035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24019_ (.A1(_15033_),
    .A2(_15035_),
    .B(net20018),
    .ZN(_15036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24020_ (.A1(_15006_),
    .A2(net19793),
    .ZN(_15037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24021_ (.A1(_15034_),
    .A2(_15037_),
    .Z(_15038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24022_ (.A1(_15038_),
    .A2(_14826_),
    .B(net20433),
    .ZN(_15039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24023_ (.A1(_15013_),
    .A2(net18751),
    .ZN(_15040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24024_ (.A1(_14566_),
    .A2(_14707_),
    .ZN(_15041_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24025_ (.A1(_15040_),
    .A2(net18770),
    .A3(_15041_),
    .ZN(_15042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24026_ (.A1(_15039_),
    .A2(_15042_),
    .ZN(_15043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24027_ (.A1(_15036_),
    .A2(_15043_),
    .B(_14515_),
    .ZN(_15044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24028_ (.A1(net18786),
    .A2(_15861_[0]),
    .ZN(_15045_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24029_ (.A1(_14738_),
    .A2(net18764),
    .A3(_15045_),
    .Z(_15046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24030_ (.A1(net17527),
    .A2(net18758),
    .ZN(_15047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24031_ (.A1(_15046_),
    .A2(_15047_),
    .B(_14485_),
    .ZN(_15048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _24032_ (.A1(net18744),
    .A2(_14549_),
    .B1(_14753_),
    .B2(_14707_),
    .ZN(_15049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24033_ (.A1(_15049_),
    .A2(net18246),
    .ZN(_15050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24034_ (.A1(_15048_),
    .A2(_15050_),
    .ZN(_15051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24035_ (.A1(net18401),
    .A2(net18754),
    .B(net18764),
    .ZN(_15052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24036_ (.A1(_14956_),
    .A2(_15052_),
    .B(net20433),
    .ZN(_15053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24037_ (.A1(_14849_),
    .A2(net18774),
    .ZN(_15054_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24038_ (.A1(_14467_),
    .A2(_14613_),
    .A3(_15054_),
    .ZN(_15055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24039_ (.A1(_15053_),
    .A2(_15055_),
    .ZN(_15056_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24040_ (.A1(_15051_),
    .A2(net20017),
    .A3(_15056_),
    .ZN(_15057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24041_ (.A1(_15044_),
    .A2(_15057_),
    .ZN(_15058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24042_ (.A1(_15031_),
    .A2(_15058_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24043_ (.I(\sa20_sub[7] ),
    .ZN(_15059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24044_ (.A1(_12006_),
    .A2(_15059_),
    .ZN(_15060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24045_ (.A1(net21344),
    .A2(net21334),
    .ZN(_15061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24046_ (.A1(_15060_),
    .A2(_15061_),
    .ZN(_15062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24047_ (.A1(_11964_),
    .A2(_15062_),
    .ZN(_15063_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24048_ (.A1(\sa20_sub[0] ),
    .A2(\sa20_sub[7] ),
    .Z(_15064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24049_ (.A1(_15064_),
    .A2(net20904),
    .ZN(_15065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24050_ (.A1(_15065_),
    .A2(_15063_),
    .ZN(_15066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24051_ (.I(_15066_),
    .ZN(_15067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24052_ (.A1(_11977_),
    .A2(net21019),
    .ZN(_15068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24053_ (.A1(_11984_),
    .A2(net21453),
    .ZN(_15069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24054_ (.A1(_15068_),
    .A2(_15069_),
    .ZN(_15070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24055_ (.I(_15070_),
    .ZN(_15071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24056_ (.A1(_15071_),
    .A2(_15067_),
    .ZN(_15072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24057_ (.A1(_15066_),
    .A2(_15070_),
    .ZN(_15073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24058_ (.A1(_15072_),
    .A2(_10378_),
    .A3(_15073_),
    .ZN(_15074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24059_ (.A1(net21501),
    .A2(\text_in_r[49] ),
    .ZN(_15075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24060_ (.A1(_15074_),
    .A2(_15075_),
    .ZN(_15076_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24061_ (.I(net21175),
    .ZN(_15077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24062_ (.A1(net19212),
    .A2(_15077_),
    .ZN(_15078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24063_ (.A1(net19774),
    .A2(net21175),
    .A3(net20975),
    .ZN(_15079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24064_ (.A1(_15079_),
    .A2(_15078_),
    .ZN(_15871_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24065_ (.A1(net21028),
    .A2(net21026),
    .ZN(_15080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24066_ (.A1(net21456),
    .A2(net21384),
    .ZN(_15081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24067_ (.A1(_15080_),
    .A2(_15081_),
    .ZN(_15082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24068_ (.A1(_15082_),
    .A2(net21284),
    .ZN(_15083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24069_ (.A1(_15080_),
    .A2(net21022),
    .A3(_15081_),
    .ZN(_15084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24070_ (.A1(_15083_),
    .A2(_15084_),
    .ZN(_15085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24071_ (.A1(_15085_),
    .A2(net20976),
    .ZN(_15086_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24072_ (.A1(_15083_),
    .A2(_15084_),
    .A3(net20882),
    .ZN(_15087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _24073_ (.A1(_15087_),
    .A2(_15086_),
    .B(net21501),
    .ZN(_15088_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24074_ (.I(\text_in_r[48] ),
    .ZN(_15089_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24075_ (.A1(_15089_),
    .A2(net21501),
    .Z(_15090_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24076_ (.A1(net20238),
    .A2(_15090_),
    .B(net21176),
    .ZN(_15091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24077_ (.A1(_15086_),
    .A2(_15087_),
    .ZN(_15092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24078_ (.A1(net21084),
    .A2(_15092_),
    .ZN(_15093_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24079_ (.I(net21176),
    .ZN(_15094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24080_ (.I(_15090_),
    .ZN(_15095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24081_ (.A1(_15093_),
    .A2(_15094_),
    .A3(_15095_),
    .ZN(_15096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24082_ (.A1(_15091_),
    .A2(_15096_),
    .ZN(_15874_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24083_ (.A1(\sa20_sub[2] ),
    .A2(\sa31_sub[2] ),
    .Z(_15097_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24084_ (.A1(\sa20_sub[2] ),
    .A2(\sa31_sub[2] ),
    .ZN(_15098_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24085_ (.A1(_15097_),
    .A2(_15098_),
    .B(net21452),
    .ZN(_15099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24086_ (.A1(_12025_),
    .A2(_12030_),
    .ZN(_15100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24087_ (.A1(net21339),
    .A2(\sa31_sub[2] ),
    .ZN(_15101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24088_ (.A1(_15100_),
    .A2(_12057_),
    .A3(_15101_),
    .ZN(_15102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24089_ (.A1(_15099_),
    .A2(_15102_),
    .ZN(_15103_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24090_ (.A1(net21396),
    .A2(net21342),
    .ZN(_15104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24091_ (.I(_15104_),
    .ZN(_15105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24092_ (.A1(_15103_),
    .A2(_15105_),
    .ZN(_15106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24093_ (.A1(_15099_),
    .A2(_15102_),
    .A3(_15104_),
    .ZN(_15107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24094_ (.A1(_15106_),
    .A2(_15107_),
    .B(net21506),
    .ZN(_15108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24095_ (.I(\text_in_r[50] ),
    .ZN(_15109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24096_ (.A1(_15109_),
    .A2(net21506),
    .Z(_15110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24097_ (.I(net21174),
    .ZN(_15111_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24098_ (.A1(_15108_),
    .A2(_15110_),
    .B(_15111_),
    .ZN(_15112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24099_ (.A1(_15106_),
    .A2(_15107_),
    .ZN(_15113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24100_ (.A1(_15113_),
    .A2(net21076),
    .ZN(_15114_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24101_ (.I(_15110_),
    .ZN(_15115_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24102_ (.A1(_15114_),
    .A2(net21174),
    .A3(_15115_),
    .ZN(_15116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24103_ (.A1(_15112_),
    .A2(_15116_),
    .ZN(_15117_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17205 (.I(_03450_),
    .Z(net17205));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24105_ (.A1(_15088_),
    .A2(_15090_),
    .B(_15094_),
    .ZN(_15118_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24106_ (.A1(_15093_),
    .A2(net21176),
    .A3(_15095_),
    .ZN(_15119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24107_ (.A1(_15118_),
    .A2(_15119_),
    .ZN(_15865_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24108_ (.A1(_15108_),
    .A2(net20935),
    .B(net21174),
    .ZN(_15120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24109_ (.A1(_15114_),
    .A2(_15111_),
    .A3(_15115_),
    .ZN(_15121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24110_ (.A1(_15120_),
    .A2(_15121_),
    .ZN(_15122_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20762 (.I(net20757),
    .Z(net20762));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24112_ (.A1(net19769),
    .A2(net17602),
    .ZN(_15123_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24113_ (.A1(net17601),
    .A2(net20015),
    .A3(net20237),
    .ZN(_15124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24114_ (.A1(net21025),
    .A2(_12032_),
    .ZN(_15125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24115_ (.A1(net21385),
    .A2(net21393),
    .ZN(_15126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24116_ (.A1(_15125_),
    .A2(_15126_),
    .ZN(_15127_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24117_ (.A1(net21450),
    .A2(_15127_),
    .Z(_15128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24118_ (.A1(_12025_),
    .A2(net20977),
    .ZN(_15129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24119_ (.A1(net21339),
    .A2(net21333),
    .ZN(_15130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24120_ (.A1(_15129_),
    .A2(_15130_),
    .ZN(_15131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24121_ (.A1(_12056_),
    .A2(_15131_),
    .ZN(_15132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24122_ (.A1(net20977),
    .A2(net21339),
    .ZN(_15133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24123_ (.A1(_12025_),
    .A2(net21333),
    .ZN(_15134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24124_ (.A1(_15133_),
    .A2(_15134_),
    .ZN(_15135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24125_ (.A1(_12069_),
    .A2(_15135_),
    .ZN(_15136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24126_ (.A1(_15132_),
    .A2(_15136_),
    .ZN(_15137_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24127_ (.I(_15137_),
    .ZN(_15138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24128_ (.A1(_15128_),
    .A2(_15138_),
    .ZN(_15139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24129_ (.A1(_15127_),
    .A2(net21450),
    .Z(_15140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24130_ (.A1(_15127_),
    .A2(net21450),
    .ZN(_15141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24131_ (.A1(_15140_),
    .A2(_15141_),
    .ZN(_15142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24132_ (.A1(_15142_),
    .A2(_15137_),
    .ZN(_15143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24133_ (.A1(_15139_),
    .A2(net21086),
    .A3(_15143_),
    .ZN(_15144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24134_ (.A1(net21506),
    .A2(\text_in_r[51] ),
    .ZN(_15145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24135_ (.A1(_15144_),
    .A2(_15145_),
    .ZN(_15146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24136_ (.I(net21173),
    .ZN(_15147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24137_ (.A1(_15146_),
    .A2(_15147_),
    .ZN(_15148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24138_ (.A1(_15144_),
    .A2(net21173),
    .A3(_15145_),
    .ZN(_15149_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24139_ (.A1(_15148_),
    .A2(_15149_),
    .ZN(_15150_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17203 (.I(_06491_),
    .Z(net17203));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17206 (.I(_03394_),
    .Z(net17206));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24142_ (.A1(_15123_),
    .A2(net454),
    .B(net18724),
    .ZN(_15153_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24143_ (.A1(\sa20_sub[4] ),
    .A2(\sa31_sub[4] ),
    .Z(_15154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24144_ (.I(_15154_),
    .ZN(_15155_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24145_ (.A1(\sa20_sub[3] ),
    .A2(net21332),
    .Z(_15156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24146_ (.A1(_15155_),
    .A2(_15156_),
    .ZN(_15157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24147_ (.I(_15156_),
    .ZN(_15158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24148_ (.A1(_15158_),
    .A2(_15154_),
    .ZN(_15159_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24149_ (.A1(_15157_),
    .A2(_15159_),
    .Z(_15160_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24150_ (.A1(net21449),
    .A2(net20897),
    .Z(_15161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24151_ (.A1(_15160_),
    .A2(_15161_),
    .ZN(_15162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24152_ (.A1(_15157_),
    .A2(_15159_),
    .ZN(_15163_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24153_ (.A1(net21449),
    .A2(net20898),
    .Z(_15164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24154_ (.A1(_15163_),
    .A2(_15164_),
    .ZN(_15165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24155_ (.A1(_15162_),
    .A2(_15165_),
    .A3(net21085),
    .ZN(_15166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24156_ (.A1(net21501),
    .A2(\text_in_r[52] ),
    .ZN(_15167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24157_ (.A1(_15166_),
    .A2(_15167_),
    .ZN(_15168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24158_ (.A1(_15168_),
    .A2(net21171),
    .ZN(_15169_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24159_ (.I(net21171),
    .ZN(_15170_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24160_ (.A1(_15166_),
    .A2(_15170_),
    .A3(_15167_),
    .ZN(_15171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24161_ (.A1(_15169_),
    .A2(_15171_),
    .ZN(_15172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20761 (.I(net20757),
    .Z(net20761));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24163_ (.I(_15868_[0]),
    .ZN(_15174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24164_ (.A1(_15174_),
    .A2(net19768),
    .ZN(_15175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24165_ (.A1(_15150_),
    .A2(_15175_),
    .ZN(_15176_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _24166_ (.I(_15176_),
    .ZN(_15177_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _24167_ (.A1(_15153_),
    .A2(net19759),
    .A3(_15177_),
    .Z(_15178_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24168_ (.A1(net21390),
    .A2(net21337),
    .ZN(_15179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24169_ (.I(\sa02_sr[5] ),
    .ZN(_15180_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24170_ (.A1(_15180_),
    .A2(_12151_),
    .Z(_15181_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24171_ (.A1(_15179_),
    .A2(_15181_),
    .Z(_15182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24172_ (.A1(_15182_),
    .A2(net21067),
    .ZN(_15183_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _24173_ (.A1(net21067),
    .A2(\text_in_r[53] ),
    .Z(_15184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24174_ (.A1(_15183_),
    .A2(_15184_),
    .ZN(_15185_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24175_ (.I(net21170),
    .ZN(_15186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24176_ (.A1(_15185_),
    .A2(_15186_),
    .ZN(_15187_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24177_ (.A1(_15183_),
    .A2(net21170),
    .A3(_15184_),
    .ZN(_15188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24178_ (.A1(_15187_),
    .A2(_15188_),
    .ZN(_15189_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17287 (.I(_01291_),
    .Z(net17287));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17201 (.I(_15268_),
    .Z(net17201));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24181_ (.I(_15872_[0]),
    .ZN(_15192_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _24182_ (.A1(net19768),
    .A2(_15192_),
    .ZN(_15193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24183_ (.A1(_15146_),
    .A2(net21173),
    .ZN(_15194_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24184_ (.A1(_15144_),
    .A2(_15147_),
    .A3(_15145_),
    .ZN(_15195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24185_ (.A1(_15194_),
    .A2(_15195_),
    .ZN(_15196_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17276 (.I(_01842_),
    .Z(net17276));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24187_ (.A1(_15193_),
    .A2(net18708),
    .ZN(_15198_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20913 (.I(_10515_),
    .Z(net20913));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24189_ (.A1(_15198_),
    .A2(net19759),
    .Z(_15200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24190_ (.A1(net19208),
    .A2(_15117_),
    .ZN(_15201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24191_ (.A1(_15201_),
    .A2(net18734),
    .Z(_15202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24192_ (.A1(net18207),
    .A2(net19211),
    .A3(net19768),
    .ZN(_15203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24193_ (.A1(_15202_),
    .A2(_15203_),
    .ZN(_15204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24194_ (.A1(_15200_),
    .A2(_15204_),
    .ZN(_15205_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24195_ (.A1(_15178_),
    .A2(net20011),
    .A3(_15205_),
    .ZN(_15206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24196_ (.A1(net19768),
    .A2(_15192_),
    .ZN(_15207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24197_ (.A1(_15207_),
    .A2(net18731),
    .Z(_15208_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24198_ (.A1(_15208_),
    .A2(net19759),
    .ZN(_15209_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _24199_ (.I(_15867_[0]),
    .ZN(_15210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24200_ (.A1(net19773),
    .A2(_15210_),
    .Z(_15211_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output387 (.I(net387),
    .Z(text_out[9]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24202_ (.A1(net19768),
    .A2(net17603),
    .Z(_15213_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output386 (.I(net386),
    .Z(text_out[99]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output385 (.I(net385),
    .Z(text_out[98]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24205_ (.A1(_15211_),
    .A2(_15213_),
    .B(net18717),
    .ZN(_15216_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output384 (.I(net384),
    .Z(text_out[97]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24207_ (.A1(_15209_),
    .A2(_15216_),
    .B(net20009),
    .ZN(_15218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24208_ (.A1(net19209),
    .A2(net19768),
    .ZN(_15219_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24209_ (.I(_15219_),
    .ZN(_15220_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _24210_ (.A1(net19768),
    .A2(_15875_[0]),
    .ZN(_15221_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output383 (.I(net383),
    .Z(text_out[96]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output382 (.I(net382),
    .Z(text_out[95]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24213_ (.A1(_15220_),
    .A2(net17514),
    .B(net18733),
    .ZN(_15224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24214_ (.A1(net18207),
    .A2(net19768),
    .ZN(_15225_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output381 (.I(net381),
    .Z(text_out[94]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24216_ (.A1(net402),
    .A2(net20013),
    .A3(net20235),
    .ZN(_15227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24217_ (.A1(_15225_),
    .A2(net18713),
    .A3(net17511),
    .ZN(_15228_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output380 (.I(net380),
    .Z(text_out[93]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24219_ (.A1(_15224_),
    .A2(_15228_),
    .A3(net19762),
    .ZN(_15230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24220_ (.A1(_15218_),
    .A2(_15230_),
    .ZN(_15231_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24221_ (.A1(\sa12_sr[5] ),
    .A2(net21336),
    .ZN(_15232_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24222_ (.I(\sa02_sr[6] ),
    .ZN(_15233_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24223_ (.A1(_15233_),
    .A2(_12190_),
    .Z(_15234_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24224_ (.A1(_15232_),
    .A2(_15234_),
    .ZN(_15235_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24225_ (.A1(net21511),
    .A2(\text_in_r[54] ),
    .Z(_15236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _24226_ (.A1(_15235_),
    .A2(net21086),
    .B(_15236_),
    .ZN(_15237_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24227_ (.A1(\u0.w[2][22] ),
    .A2(_15237_),
    .Z(_15238_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24228_ (.I(_15238_),
    .ZN(_15239_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output379 (.I(net379),
    .Z(text_out[92]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24230_ (.A1(_15206_),
    .A2(_15231_),
    .A3(net20232),
    .ZN(_15241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24231_ (.A1(net18207),
    .A2(net19208),
    .A3(net19768),
    .ZN(_15242_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24232_ (.A1(_15192_),
    .A2(net20014),
    .A3(net20236),
    .ZN(_15243_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24233_ (.A1(_15242_),
    .A2(net18711),
    .A3(_15243_),
    .ZN(_15244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24234_ (.A1(net19211),
    .A2(_15117_),
    .ZN(_15245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24235_ (.A1(net19768),
    .A2(_15210_),
    .ZN(_15246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24236_ (.A1(_15245_),
    .A2(_15246_),
    .ZN(_15247_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output378 (.I(net378),
    .Z(text_out[91]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24238_ (.A1(_15168_),
    .A2(_15170_),
    .ZN(_15249_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24239_ (.A1(_15166_),
    .A2(net21171),
    .A3(_15167_),
    .ZN(_15250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24240_ (.A1(_15249_),
    .A2(_15250_),
    .ZN(_15251_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output377 (.I(net377),
    .Z(text_out[90]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24242_ (.A1(_15247_),
    .A2(net18731),
    .B(net19747),
    .ZN(_15253_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24243_ (.A1(net19771),
    .A2(net17603),
    .Z(_15254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24244_ (.A1(_15254_),
    .A2(net18708),
    .ZN(_15255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24245_ (.A1(_15244_),
    .A2(_15253_),
    .A3(_15255_),
    .ZN(_15256_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24246_ (.I(_15227_),
    .ZN(_15257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _24247_ (.A1(net18708),
    .A2(_15257_),
    .B(_15172_),
    .ZN(_15258_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output376 (.I(net376),
    .Z(text_out[8]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24249_ (.A1(net18732),
    .A2(_15888_[0]),
    .ZN(_15260_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24250_ (.I(_15189_),
    .ZN(_15261_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output375 (.I(net375),
    .Z(text_out[89]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24252_ (.A1(_15258_),
    .A2(_15260_),
    .B(net19742),
    .ZN(_15263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24253_ (.A1(_15256_),
    .A2(_15263_),
    .ZN(_15264_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24254_ (.I(_15877_[0]),
    .ZN(_15265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24255_ (.A1(_15265_),
    .A2(net20013),
    .A3(net20234),
    .ZN(_15266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24256_ (.A1(_15150_),
    .A2(_15266_),
    .ZN(_15267_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24257_ (.I(_15267_),
    .ZN(_15268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24258_ (.A1(net17841),
    .A2(net17200),
    .ZN(_15269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24259_ (.A1(_15213_),
    .A2(net18718),
    .ZN(_15270_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24260_ (.A1(_15269_),
    .A2(net19760),
    .A3(net17299),
    .ZN(_15271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24261_ (.A1(_15213_),
    .A2(net18727),
    .ZN(_15272_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24262_ (.A1(_15272_),
    .A2(net19747),
    .Z(_15273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24263_ (.A1(_15117_),
    .A2(_15875_[0]),
    .ZN(_15274_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24264_ (.A1(_15274_),
    .A2(net18708),
    .Z(_15275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24265_ (.A1(net17841),
    .A2(_15275_),
    .ZN(_15276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24266_ (.A1(_15273_),
    .A2(_15276_),
    .ZN(_15277_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output374 (.I(net374),
    .Z(text_out[88]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24268_ (.A1(_15271_),
    .A2(_15277_),
    .A3(net19744),
    .ZN(_15279_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output373 (.I(net373),
    .Z(text_out[87]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24270_ (.A1(_15264_),
    .A2(_15279_),
    .A3(net20429),
    .ZN(_15281_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24271_ (.A1(net21445),
    .A2(net21387),
    .Z(_15282_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24272_ (.A1(net21335),
    .A2(_15282_),
    .Z(_15283_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _24273_ (.A1(net21332),
    .A2(net21274),
    .A3(_15283_),
    .Z(_15284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _24274_ (.I0(_15284_),
    .I1(\text_in_r[55] ),
    .S(net21505),
    .Z(_15285_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24275_ (.A1(\u0.w[2][23] ),
    .A2(_15285_),
    .ZN(_15286_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output372 (.I(net372),
    .Z(text_out[86]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24277_ (.I(_15286_),
    .ZN(_15288_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24278_ (.A1(_15241_),
    .A2(_15281_),
    .A3(net20428),
    .ZN(_15289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24279_ (.A1(_15117_),
    .A2(_15174_),
    .ZN(_15290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24280_ (.A1(_15290_),
    .A2(net18729),
    .Z(_15291_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24281_ (.A1(_15291_),
    .A2(net19759),
    .ZN(_15292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24282_ (.A1(_15076_),
    .A2(net21175),
    .ZN(_15293_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24283_ (.A1(_15074_),
    .A2(_15077_),
    .A3(_15075_),
    .ZN(_15294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24284_ (.A1(_15293_),
    .A2(_15294_),
    .ZN(_15866_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24285_ (.A1(net18201),
    .A2(_15117_),
    .ZN(_15295_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output371 (.I(net371),
    .Z(text_out[85]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24287_ (.A1(_15295_),
    .A2(net18727),
    .ZN(_15297_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24288_ (.I(_15297_),
    .ZN(_15298_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24289_ (.I(_15175_),
    .ZN(_15299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24290_ (.A1(_15299_),
    .A2(net18715),
    .ZN(_15300_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24291_ (.A1(_15292_),
    .A2(_15298_),
    .A3(_15300_),
    .Z(_15301_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _24292_ (.A1(_15246_),
    .A2(net18727),
    .Z(_15302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24293_ (.A1(_15221_),
    .A2(net18708),
    .ZN(_15303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24294_ (.A1(_15302_),
    .A2(_15303_),
    .Z(_15304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24295_ (.A1(net19772),
    .A2(net17605),
    .ZN(_15305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24296_ (.A1(_15177_),
    .A2(_15305_),
    .ZN(_15306_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output370 (.I(net370),
    .Z(text_out[84]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24298_ (.A1(_15304_),
    .A2(_15306_),
    .B(net19747),
    .ZN(_15308_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24299_ (.A1(_15301_),
    .A2(_15308_),
    .B(net20009),
    .ZN(_15309_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24300_ (.I(_15875_[0]),
    .ZN(_15310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24301_ (.A1(net19768),
    .A2(_15310_),
    .ZN(_15311_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24302_ (.A1(net17605),
    .A2(net19768),
    .B(_15311_),
    .ZN(_15312_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output369 (.I(net369),
    .Z(text_out[83]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24304_ (.A1(_15312_),
    .A2(net18735),
    .B(net19747),
    .ZN(_15314_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24305_ (.A1(net18206),
    .A2(net19211),
    .A3(net19772),
    .ZN(_15315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24306_ (.A1(net17307),
    .A2(net18717),
    .Z(_15316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24307_ (.A1(_15315_),
    .A2(_15316_),
    .ZN(_15317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24308_ (.A1(_15314_),
    .A2(_15317_),
    .ZN(_15318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24309_ (.A1(_15219_),
    .A2(net18708),
    .Z(_15319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24310_ (.A1(net18203),
    .A2(net19208),
    .ZN(_15320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24311_ (.A1(_15319_),
    .A2(_15320_),
    .ZN(_15321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24312_ (.A1(net18207),
    .A2(net19208),
    .ZN(_15322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24313_ (.A1(net17832),
    .A2(net18731),
    .A3(_15245_),
    .ZN(_15323_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output368 (.I(net368),
    .Z(text_out[82]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24315_ (.A1(_15321_),
    .A2(_15323_),
    .A3(net19752),
    .ZN(_15325_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24316_ (.A1(_15318_),
    .A2(net19744),
    .A3(_15325_),
    .ZN(_15326_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24317_ (.A1(_15309_),
    .A2(_15326_),
    .A3(net20429),
    .ZN(_15327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24318_ (.A1(_15201_),
    .A2(net18708),
    .ZN(_15328_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24319_ (.A1(_15328_),
    .A2(net19759),
    .Z(_15329_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24320_ (.A1(net18207),
    .A2(net19208),
    .A3(net19772),
    .ZN(_15330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24321_ (.A1(_15330_),
    .A2(_15208_),
    .ZN(_15331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24322_ (.A1(_15329_),
    .A2(_15331_),
    .B(net20009),
    .ZN(_15332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24323_ (.A1(net19208),
    .A2(net19768),
    .ZN(_15333_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24324_ (.A1(_15333_),
    .A2(net18720),
    .Z(_15334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24325_ (.A1(_15334_),
    .A2(_15330_),
    .ZN(_15335_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _24326_ (.I(_15881_[0]),
    .ZN(_15336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24327_ (.A1(_15117_),
    .A2(_15336_),
    .ZN(_15337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24328_ (.A1(_15177_),
    .A2(net17296),
    .ZN(_15338_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24329_ (.A1(_15335_),
    .A2(_15338_),
    .A3(net19752),
    .ZN(_15339_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output367 (.I(net367),
    .Z(text_out[81]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24331_ (.A1(_15332_),
    .A2(_15339_),
    .B(net20429),
    .ZN(_15341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24332_ (.A1(_15270_),
    .A2(net19759),
    .ZN(_15342_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24333_ (.A1(_15342_),
    .A2(_15297_),
    .ZN(_15343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24334_ (.A1(_15343_),
    .A2(_15204_),
    .ZN(_15344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24335_ (.A1(net19768),
    .A2(_15336_),
    .ZN(_15345_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24336_ (.A1(_15345_),
    .A2(_15150_),
    .Z(_15346_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output366 (.I(net366),
    .Z(text_out[80]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24338_ (.A1(_15346_),
    .A2(net18707),
    .B(net19759),
    .ZN(_15348_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output365 (.I(net365),
    .Z(text_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24340_ (.A1(net18203),
    .A2(net19768),
    .ZN(_15350_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24341_ (.A1(_15330_),
    .A2(net18721),
    .A3(net17829),
    .ZN(_15351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24342_ (.A1(_15348_),
    .A2(_15351_),
    .ZN(_15352_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output364 (.I(net364),
    .Z(text_out[79]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24344_ (.A1(_15344_),
    .A2(_15352_),
    .A3(net20009),
    .ZN(_15354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24345_ (.A1(_15354_),
    .A2(_15341_),
    .B(_15288_),
    .ZN(_15355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24346_ (.A1(_15327_),
    .A2(_15355_),
    .ZN(_15356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24347_ (.A1(_15289_),
    .A2(_15356_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24348_ (.A1(_15208_),
    .A2(net17837),
    .ZN(_15357_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output363 (.I(net363),
    .Z(text_out[78]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24350_ (.A1(net18706),
    .A2(_15305_),
    .A3(net18719),
    .ZN(_15359_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24351_ (.A1(_15357_),
    .A2(net19759),
    .A3(_15359_),
    .ZN(_15360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24352_ (.A1(net17516),
    .A2(net18717),
    .B(net19759),
    .ZN(_15361_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _24353_ (.A1(_15245_),
    .A2(net18731),
    .Z(_15362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24354_ (.A1(net17302),
    .A2(net17511),
    .ZN(_15363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24355_ (.A1(_15363_),
    .A2(net18732),
    .ZN(_15364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24356_ (.A1(_15361_),
    .A2(_15362_),
    .A3(_15364_),
    .ZN(_15365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24357_ (.A1(_15360_),
    .A2(_15365_),
    .A3(net19745),
    .ZN(_15366_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24358_ (.I(_15328_),
    .ZN(_15367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24359_ (.A1(_15367_),
    .A2(_15203_),
    .ZN(_15368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24360_ (.A1(_15176_),
    .A2(net19765),
    .Z(_15369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24361_ (.A1(_15368_),
    .A2(_15369_),
    .B(net19742),
    .ZN(_15370_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24362_ (.A1(_15345_),
    .A2(net18709),
    .Z(_15371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24363_ (.I(_15869_[0]),
    .ZN(_15372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24364_ (.A1(net19770),
    .A2(_15372_),
    .ZN(_15373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24365_ (.A1(_15371_),
    .A2(_15373_),
    .B(net19765),
    .ZN(_15374_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24366_ (.A1(net19768),
    .A2(net17604),
    .Z(_15375_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24367_ (.I(_15375_),
    .ZN(_15376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24368_ (.A1(_15315_),
    .A2(net18734),
    .A3(_15376_),
    .ZN(_15377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24369_ (.A1(_15374_),
    .A2(_15377_),
    .ZN(_15378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24370_ (.A1(_15370_),
    .A2(_15378_),
    .ZN(_15379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24371_ (.A1(_15366_),
    .A2(_15379_),
    .B(net20429),
    .ZN(_15380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24372_ (.A1(_15334_),
    .A2(_15305_),
    .ZN(_15381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24373_ (.A1(net18726),
    .A2(net19768),
    .Z(_15382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24374_ (.A1(net18206),
    .A2(net19211),
    .ZN(_15383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24375_ (.A1(_15382_),
    .A2(_15383_),
    .ZN(_15384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24376_ (.A1(_15381_),
    .A2(_15384_),
    .ZN(_15385_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _24377_ (.A1(net18708),
    .A2(net19768),
    .ZN(_15386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24378_ (.A1(_15386_),
    .A2(_15322_),
    .ZN(_15387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24379_ (.A1(_15387_),
    .A2(net19747),
    .ZN(_15388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24380_ (.A1(_15203_),
    .A2(_15275_),
    .ZN(_15389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24381_ (.A1(_15389_),
    .A2(net19763),
    .ZN(_15390_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24382_ (.A1(_15385_),
    .A2(net17292),
    .B(_15390_),
    .ZN(_15391_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24383_ (.I(_15891_[0]),
    .ZN(_15392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24384_ (.A1(net18734),
    .A2(_15392_),
    .Z(_15393_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output362 (.I(net362),
    .Z(text_out[77]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24386_ (.A1(_15393_),
    .A2(net19754),
    .B(net20009),
    .ZN(_15395_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24387_ (.A1(net20009),
    .A2(net19747),
    .Z(_15396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24388_ (.A1(_15357_),
    .A2(_15396_),
    .ZN(_15397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24389_ (.A1(net18207),
    .A2(net19772),
    .ZN(_15398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24390_ (.A1(_15319_),
    .A2(_15398_),
    .ZN(_15399_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24391_ (.I(_15399_),
    .ZN(_15400_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24392_ (.A1(_15397_),
    .A2(_15400_),
    .B(net20429),
    .ZN(_15401_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24393_ (.A1(_15391_),
    .A2(_15395_),
    .B(_15401_),
    .ZN(_15402_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24394_ (.A1(_15380_),
    .A2(_15402_),
    .B(net20631),
    .ZN(_15403_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output361 (.I(net361),
    .Z(text_out[76]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24396_ (.A1(net17828),
    .A2(net19768),
    .A3(net18710),
    .ZN(_15405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24397_ (.A1(_15337_),
    .A2(net18731),
    .Z(_15406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24398_ (.A1(_15406_),
    .A2(_15350_),
    .ZN(_15407_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24399_ (.A1(_15405_),
    .A2(_15407_),
    .A3(net19747),
    .ZN(_15408_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24400_ (.A1(net19768),
    .A2(net17602),
    .Z(_15409_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output360 (.I(net360),
    .Z(text_out[75]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24402_ (.A1(_15409_),
    .A2(net18710),
    .B(net19747),
    .ZN(_15411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24403_ (.A1(_15377_),
    .A2(_15411_),
    .ZN(_15412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24404_ (.A1(_15408_),
    .A2(_15412_),
    .A3(net19746),
    .ZN(_15413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24405_ (.A1(net18203),
    .A2(net19211),
    .ZN(_15414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24406_ (.A1(_15202_),
    .A2(_15414_),
    .ZN(_15415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24407_ (.A1(net18708),
    .A2(_15227_),
    .Z(_15416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24408_ (.A1(_15416_),
    .A2(net18703),
    .ZN(_15417_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24409_ (.A1(_15415_),
    .A2(net19766),
    .A3(_15417_),
    .ZN(_15418_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24410_ (.A1(net17216),
    .A2(net17305),
    .B(net18731),
    .ZN(_15419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24411_ (.A1(_15247_),
    .A2(net18708),
    .ZN(_15420_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24412_ (.A1(_15419_),
    .A2(_15420_),
    .A3(net19747),
    .ZN(_15421_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24413_ (.A1(_15418_),
    .A2(_15421_),
    .A3(net20009),
    .ZN(_15422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24414_ (.A1(_15413_),
    .A2(_15422_),
    .A3(net20233),
    .ZN(_15423_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24415_ (.A1(_15346_),
    .A2(net17298),
    .B(net19747),
    .ZN(_15424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24416_ (.A1(_15424_),
    .A2(_15244_),
    .ZN(_15425_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24417_ (.A1(_15198_),
    .A2(net19747),
    .Z(_15426_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output359 (.I(net359),
    .Z(text_out[74]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24419_ (.A1(_15398_),
    .A2(net18732),
    .ZN(_15428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24420_ (.A1(_15426_),
    .A2(_15350_),
    .A3(_15428_),
    .ZN(_15429_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24421_ (.A1(_15425_),
    .A2(_15429_),
    .A3(net20009),
    .ZN(_15430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24422_ (.A1(net18708),
    .A2(_15207_),
    .Z(_15431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24423_ (.A1(net17215),
    .A2(net18704),
    .ZN(_15432_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24424_ (.A1(net18707),
    .A2(net17309),
    .A3(net18732),
    .ZN(_15433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24425_ (.A1(_15432_),
    .A2(_15433_),
    .A3(net19754),
    .ZN(_15434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24426_ (.A1(_15386_),
    .A2(net17831),
    .B(net19747),
    .ZN(_15435_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24427_ (.A1(_15320_),
    .A2(_15225_),
    .A3(net18708),
    .ZN(_15436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24428_ (.A1(_15435_),
    .A2(_15436_),
    .ZN(_15437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24429_ (.A1(_15434_),
    .A2(_15437_),
    .A3(net19745),
    .ZN(_15438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24430_ (.A1(_15438_),
    .A2(net20429),
    .A3(_15430_),
    .ZN(_15439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24431_ (.A1(_15423_),
    .A2(net20427),
    .A3(_15439_),
    .ZN(_15440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24432_ (.A1(_15403_),
    .A2(_15440_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24433_ (.A1(net17835),
    .A2(net18724),
    .A3(net17519),
    .ZN(_15441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24434_ (.A1(net20236),
    .A2(net20014),
    .A3(net17600),
    .ZN(_15442_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24435_ (.A1(_15219_),
    .A2(_15442_),
    .A3(net18723),
    .ZN(_15443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24436_ (.A1(_15441_),
    .A2(net19748),
    .A3(_15443_),
    .ZN(_15444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24437_ (.A1(_15333_),
    .A2(net18708),
    .A3(net17300),
    .ZN(_15445_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24438_ (.A1(net17306),
    .A2(net18724),
    .A3(net17512),
    .ZN(_15446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24439_ (.A1(_15445_),
    .A2(_15446_),
    .ZN(_15447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24440_ (.A1(_15447_),
    .A2(net19757),
    .ZN(_15448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24441_ (.A1(_15444_),
    .A2(net19742),
    .A3(_15448_),
    .ZN(_15449_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24442_ (.A1(net18204),
    .A2(net19769),
    .ZN(_15450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24443_ (.A1(net18724),
    .A2(_15243_),
    .ZN(_15451_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24444_ (.A1(_15450_),
    .A2(_15451_),
    .ZN(_15452_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24445_ (.A1(_15452_),
    .A2(_15153_),
    .B(net19757),
    .ZN(_15453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24446_ (.A1(_15333_),
    .A2(net18724),
    .A3(_15243_),
    .ZN(_15454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24447_ (.A1(_15442_),
    .A2(net454),
    .ZN(_15455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24448_ (.A1(_15455_),
    .A2(net18723),
    .ZN(_15456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24449_ (.A1(_15454_),
    .A2(_15456_),
    .ZN(_15457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24450_ (.A1(_15457_),
    .A2(net19748),
    .ZN(_15458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24451_ (.A1(_15453_),
    .A2(_15458_),
    .A3(net20009),
    .ZN(_15459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24452_ (.A1(_15449_),
    .A2(_15459_),
    .ZN(_15460_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24453_ (.A1(_15460_),
    .A2(net20231),
    .B(_15288_),
    .ZN(_15461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24454_ (.A1(_15322_),
    .A2(_15225_),
    .A3(net18734),
    .ZN(_15462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24455_ (.A1(net413),
    .A2(_15431_),
    .ZN(_15463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24456_ (.A1(_15463_),
    .A2(_15462_),
    .ZN(_15464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24457_ (.A1(net19754),
    .A2(_15464_),
    .ZN(_15465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24458_ (.A1(_15333_),
    .A2(_15243_),
    .ZN(_15466_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24459_ (.A1(_15466_),
    .A2(net18727),
    .A3(_15350_),
    .ZN(_15467_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24460_ (.A1(_15467_),
    .A2(net19759),
    .A3(_15228_),
    .ZN(_15468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24461_ (.A1(_15468_),
    .A2(_15465_),
    .ZN(_15469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24462_ (.A1(net20011),
    .A2(_15469_),
    .ZN(_15470_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24463_ (.A1(net17834),
    .A2(net18727),
    .A3(net17295),
    .ZN(_15471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24464_ (.A1(_15330_),
    .A2(net18714),
    .ZN(_15472_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24465_ (.A1(_15471_),
    .A2(net19762),
    .A3(_15472_),
    .ZN(_15473_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24466_ (.A1(_15220_),
    .A2(net17509),
    .B(net18733),
    .ZN(_15474_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24467_ (.A1(_15398_),
    .A2(net18712),
    .A3(net17309),
    .ZN(_15475_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24468_ (.A1(_15474_),
    .A2(_15475_),
    .A3(net19753),
    .ZN(_15476_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24469_ (.A1(_15473_),
    .A2(net19744),
    .A3(_15476_),
    .ZN(_15477_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24470_ (.A1(net20429),
    .A2(_15477_),
    .A3(_15470_),
    .ZN(_15478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24471_ (.A1(_15478_),
    .A2(_15461_),
    .ZN(_15479_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24472_ (.A1(net17838),
    .A2(net18707),
    .ZN(_15480_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24473_ (.A1(_15192_),
    .A2(_15372_),
    .Z(_15481_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24474_ (.A1(net19770),
    .A2(_15481_),
    .Z(_15482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24475_ (.I(_15482_),
    .ZN(_15483_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24476_ (.A1(_15480_),
    .A2(_15483_),
    .B(net18727),
    .ZN(_15484_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24477_ (.A1(_15484_),
    .A2(net19747),
    .A3(_15389_),
    .ZN(_15485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24478_ (.A1(_15302_),
    .A2(net19759),
    .Z(_15486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24479_ (.A1(_15177_),
    .A2(net17303),
    .ZN(_15487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24480_ (.A1(_15486_),
    .A2(_15487_),
    .B(net20009),
    .ZN(_15488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24481_ (.A1(_15485_),
    .A2(_15488_),
    .ZN(_15489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24482_ (.A1(_15895_[0]),
    .A2(net18714),
    .B(net19766),
    .ZN(_15490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24483_ (.A1(_15462_),
    .A2(_15490_),
    .B(net19742),
    .ZN(_15491_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _24484_ (.A1(net18714),
    .A2(_15886_[0]),
    .Z(_15492_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24485_ (.A1(_15472_),
    .A2(net19766),
    .A3(_15492_),
    .ZN(_15493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24486_ (.A1(_15491_),
    .A2(_15493_),
    .ZN(_15494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24487_ (.A1(_15489_),
    .A2(_15494_),
    .A3(net20430),
    .ZN(_15495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24488_ (.A1(_15225_),
    .A2(net18714),
    .ZN(_15496_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24489_ (.A1(_15496_),
    .A2(_15211_),
    .ZN(_15497_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24490_ (.A1(_15311_),
    .A2(net18734),
    .A3(net17511),
    .Z(_15498_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24491_ (.A1(_15497_),
    .A2(_15498_),
    .B(net19754),
    .ZN(_15499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24492_ (.A1(_15320_),
    .A2(_15225_),
    .A3(net18734),
    .ZN(_15500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24493_ (.A1(net18714),
    .A2(_15392_),
    .ZN(_15501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24494_ (.A1(_15500_),
    .A2(net19766),
    .A3(_15501_),
    .ZN(_15502_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24495_ (.A1(_15499_),
    .A2(net20009),
    .A3(_15502_),
    .ZN(_15503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24496_ (.A1(net17840),
    .A2(_15291_),
    .ZN(_15504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24497_ (.A1(_15888_[0]),
    .A2(net18713),
    .B(net19747),
    .ZN(_15505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24498_ (.A1(_15504_),
    .A2(_15505_),
    .B(net20009),
    .ZN(_15506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24499_ (.A1(net17836),
    .A2(net18727),
    .A3(_15333_),
    .ZN(_15507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24500_ (.A1(_15228_),
    .A2(_15507_),
    .A3(net19747),
    .ZN(_15508_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24501_ (.A1(_15506_),
    .A2(_15508_),
    .B(net20429),
    .ZN(_15509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24502_ (.A1(_15503_),
    .A2(_15509_),
    .ZN(_15510_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24503_ (.A1(_15495_),
    .A2(net20427),
    .A3(_15510_),
    .ZN(_15511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24504_ (.A1(_15511_),
    .A2(_15479_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24505_ (.A1(_15382_),
    .A2(net17518),
    .B(net19765),
    .ZN(_15512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24506_ (.A1(_15245_),
    .A2(_15311_),
    .Z(_15513_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24507_ (.A1(_15513_),
    .A2(net18726),
    .Z(_15514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24508_ (.I(_15290_),
    .ZN(_15515_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24509_ (.A1(_15515_),
    .A2(net18724),
    .Z(_15516_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24510_ (.I(_15516_),
    .ZN(_15517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24511_ (.A1(_15512_),
    .A2(_15514_),
    .A3(_15517_),
    .ZN(_15518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24512_ (.A1(_15295_),
    .A2(net18708),
    .ZN(_15519_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24513_ (.A1(_15519_),
    .A2(_15375_),
    .Z(_15520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24514_ (.A1(_15346_),
    .A2(net17303),
    .ZN(_15521_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24515_ (.A1(_15520_),
    .A2(net19765),
    .A3(_15521_),
    .ZN(_15522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24516_ (.A1(net19746),
    .A2(_15522_),
    .A3(_15518_),
    .ZN(_15523_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24517_ (.A1(net17836),
    .A2(net18715),
    .A3(net18702),
    .ZN(_15524_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24518_ (.A1(_15292_),
    .A2(_15524_),
    .B(net19742),
    .ZN(_15525_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24519_ (.A1(_15319_),
    .A2(net17831),
    .ZN(_15526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24520_ (.A1(_15177_),
    .A2(net17836),
    .ZN(_15527_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24521_ (.A1(_15526_),
    .A2(_15527_),
    .A3(net19759),
    .ZN(_15528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24522_ (.A1(_15525_),
    .A2(_15528_),
    .B(net20233),
    .ZN(_15529_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24523_ (.A1(_15529_),
    .A2(_15523_),
    .B(net20631),
    .ZN(_15530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24524_ (.A1(_15295_),
    .A2(net18731),
    .Z(_15531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24525_ (.A1(_15531_),
    .A2(_15513_),
    .ZN(_15532_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24526_ (.A1(_15416_),
    .A2(_15350_),
    .A3(_15333_),
    .ZN(_15533_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24527_ (.A1(_15532_),
    .A2(net19765),
    .A3(_15533_),
    .Z(_15534_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _24528_ (.A1(_15299_),
    .A2(_15150_),
    .A3(_15221_),
    .Z(_15535_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24529_ (.A1(_15535_),
    .A2(net19747),
    .A3(_15323_),
    .Z(_15536_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24530_ (.A1(_15534_),
    .A2(_15536_),
    .B(net19743),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _24531_ (.A1(_15320_),
    .A2(net18705),
    .A3(net19757),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24532_ (.I(_15382_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24533_ (.A1(_00550_),
    .A2(_00551_),
    .B(net19742),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24534_ (.A1(net18708),
    .A2(net17300),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24535_ (.A1(net17214),
    .A2(net17294),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24536_ (.A1(_15407_),
    .A2(_00554_),
    .A3(net19755),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24537_ (.A1(_00552_),
    .A2(_00555_),
    .B(net20429),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24538_ (.A1(_00556_),
    .A2(_00549_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24539_ (.A1(_15530_),
    .A2(_00557_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24540_ (.I(_15124_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24541_ (.A1(net18724),
    .A2(net17289),
    .B(net20009),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24542_ (.A1(_00560_),
    .A2(_15445_),
    .B(net19749),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24543_ (.A1(_15367_),
    .A2(net17308),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24544_ (.A1(net19768),
    .A2(_15481_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24545_ (.A1(_00563_),
    .A2(net18727),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _24546_ (.I(net412),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _24547_ (.A1(_00564_),
    .A2(_00565_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24548_ (.A1(_00562_),
    .A2(net20009),
    .A3(_00566_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24549_ (.A1(_00561_),
    .A2(_00567_),
    .B(net20233),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24550_ (.A1(_15275_),
    .A2(_15225_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24551_ (.A1(_00569_),
    .A2(_15516_),
    .B(net20009),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24552_ (.I(_15300_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _24553_ (.A1(_00571_),
    .A2(net19742),
    .B1(net18728),
    .B2(net17517),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24554_ (.A1(_00570_),
    .A2(_00572_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24555_ (.A1(_00573_),
    .A2(net19747),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24556_ (.A1(_00574_),
    .A2(_00568_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24557_ (.A1(net17201),
    .A2(net17213),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24558_ (.A1(_15389_),
    .A2(_00576_),
    .A3(net19759),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24559_ (.I(_15443_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24560_ (.A1(_00578_),
    .A2(net19747),
    .B(net19742),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24561_ (.A1(_00577_),
    .A2(_00579_),
    .B(net20429),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24562_ (.I(_15201_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24563_ (.A1(_00581_),
    .A2(_00559_),
    .B(net18730),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24564_ (.A1(_15316_),
    .A2(net17296),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24565_ (.A1(_00582_),
    .A2(_00583_),
    .A3(net19747),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24566_ (.A1(_15253_),
    .A2(_15436_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24567_ (.A1(_00584_),
    .A2(_00585_),
    .A3(net19742),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24568_ (.A1(_00580_),
    .A2(_00586_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24569_ (.A1(_00587_),
    .A2(_00575_),
    .A3(net20631),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24570_ (.A1(_00588_),
    .A2(_00558_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24571_ (.A1(_15268_),
    .A2(_15350_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24572_ (.A1(_15450_),
    .A2(net18722),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24573_ (.A1(_15220_),
    .A2(net18719),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _24574_ (.A1(net19747),
    .A2(_00589_),
    .A3(_00590_),
    .A4(_00591_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24575_ (.I(_15879_[0]),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24576_ (.A1(_00593_),
    .A2(net18722),
    .B(net19747),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24577_ (.A1(net18724),
    .A2(net17513),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24578_ (.A1(_00595_),
    .A2(_00594_),
    .B(net20009),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24579_ (.A1(_00596_),
    .A2(_00592_),
    .B(net20231),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24580_ (.A1(_15322_),
    .A2(_15295_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _24581_ (.A1(_00598_),
    .A2(net18727),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24582_ (.A1(net17200),
    .A2(net18706),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24583_ (.A1(_00599_),
    .A2(_00600_),
    .A3(net19752),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24584_ (.A1(_15216_),
    .A2(_15323_),
    .A3(net19759),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24585_ (.A1(_00601_),
    .A2(_00602_),
    .A3(net20012),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24586_ (.A1(_00603_),
    .A2(_00597_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24587_ (.A1(_15302_),
    .A2(net19747),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24588_ (.A1(_00605_),
    .A2(_15298_),
    .A3(_15357_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24589_ (.A1(_15319_),
    .A2(net17296),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24590_ (.A1(net18198),
    .A2(net19747),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24591_ (.A1(_00607_),
    .A2(_00608_),
    .B(net19742),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24592_ (.A1(_00606_),
    .A2(_00609_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24593_ (.A1(_15373_),
    .A2(net18708),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24594_ (.A1(_00611_),
    .A2(net19766),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24595_ (.A1(_15315_),
    .A2(net18735),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24596_ (.A1(_00612_),
    .A2(_00613_),
    .B(net20009),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24597_ (.A1(net17215),
    .A2(net17511),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24598_ (.A1(_15204_),
    .A2(_00615_),
    .A3(net19767),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24599_ (.A1(_00614_),
    .A2(_00616_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24600_ (.A1(_00617_),
    .A2(_00610_),
    .A3(net20232),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24601_ (.A1(_00604_),
    .A2(net20631),
    .A3(_00618_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24602_ (.A1(_15531_),
    .A2(net17839),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24603_ (.A1(_00620_),
    .A2(net19754),
    .A3(_15463_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24604_ (.A1(_15398_),
    .A2(net17302),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24605_ (.A1(_00622_),
    .A2(net18737),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24606_ (.A1(_15244_),
    .A2(net19767),
    .A3(_00623_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24607_ (.A1(_00621_),
    .A2(_00624_),
    .A3(net20009),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24608_ (.A1(_15257_),
    .A2(net18734),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24609_ (.A1(_00626_),
    .A2(net17291),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24610_ (.A1(_00627_),
    .A2(_15426_),
    .B(net20009),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24611_ (.A1(_15371_),
    .A2(net17298),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24612_ (.A1(_15269_),
    .A2(_00629_),
    .A3(net19760),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24613_ (.A1(_00628_),
    .A2(_00630_),
    .B(net20232),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24614_ (.A1(_00625_),
    .A2(_00631_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24615_ (.A1(_15295_),
    .A2(_15219_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24616_ (.A1(_00633_),
    .A2(net18728),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24617_ (.A1(_00634_),
    .A2(_15381_),
    .A3(net19760),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24618_ (.A1(net17516),
    .A2(net19759),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24619_ (.A1(_00636_),
    .A2(net17217),
    .B(net20009),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24620_ (.A1(_00635_),
    .A2(_00637_),
    .B(net20429),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24621_ (.A1(net17504),
    .A2(net18721),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24622_ (.A1(net17829),
    .A2(net18727),
    .A3(_15305_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24623_ (.A1(_00639_),
    .A2(net19752),
    .A3(_00640_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24624_ (.A1(_15500_),
    .A2(_15399_),
    .A3(net19761),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24625_ (.A1(_00641_),
    .A2(_00642_),
    .A3(net20012),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24626_ (.A1(_00638_),
    .A2(_00643_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24627_ (.A1(_00632_),
    .A2(_00644_),
    .A3(net20428),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24628_ (.A1(_00619_),
    .A2(_00645_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24629_ (.A1(net18203),
    .A2(net18732),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24630_ (.A1(_00599_),
    .A2(net19759),
    .A3(_00646_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24631_ (.A1(_15203_),
    .A2(net17508),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24632_ (.A1(_15367_),
    .A2(_15383_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24633_ (.A1(_00649_),
    .A2(net19747),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24634_ (.A1(_00648_),
    .A2(net18731),
    .B(_00650_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24635_ (.A1(_00647_),
    .A2(_00651_),
    .B(net19742),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24636_ (.A1(_00611_),
    .A2(_15225_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24637_ (.A1(_00653_),
    .A2(_00626_),
    .B(net19756),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24638_ (.A1(net18708),
    .A2(_15442_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _24639_ (.A1(net17218),
    .A2(_15211_),
    .B(_00655_),
    .C(net19765),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24640_ (.A1(_00654_),
    .A2(_00656_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24641_ (.A1(_00657_),
    .A2(net20009),
    .B(net20232),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24642_ (.A1(_00652_),
    .A2(_00658_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24643_ (.A1(_15316_),
    .A2(net19747),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24644_ (.A1(_00660_),
    .A2(_00582_),
    .B(net19742),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24645_ (.A1(_15388_),
    .A2(net650),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24646_ (.A1(_00661_),
    .A2(_00662_),
    .B(net20429),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24647_ (.A1(_15406_),
    .A2(net17304),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24648_ (.A1(_15343_),
    .A2(_00664_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24649_ (.A1(net17841),
    .A2(_00553_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24650_ (.A1(net18728),
    .A2(net17602),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24651_ (.A1(_15273_),
    .A2(_00666_),
    .A3(_00667_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24652_ (.A1(_00665_),
    .A2(_00668_),
    .A3(net19744),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24653_ (.A1(_00663_),
    .A2(_00669_),
    .B(net20631),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24654_ (.A1(_00659_),
    .A2(_00670_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24655_ (.A1(net19209),
    .A2(net18728),
    .B(net19747),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24656_ (.A1(_15321_),
    .A2(_00672_),
    .B(net20009),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24657_ (.A1(net17830),
    .A2(_15177_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24658_ (.A1(_00553_),
    .A2(_15350_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24659_ (.A1(_00674_),
    .A2(_00675_),
    .A3(net19752),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24660_ (.A1(_00676_),
    .A2(_00673_),
    .B(net20429),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24661_ (.A1(_15200_),
    .A2(_15204_),
    .A3(_00591_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24662_ (.A1(_15203_),
    .A2(net18711),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24663_ (.A1(net17514),
    .A2(net18733),
    .B(net19759),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24664_ (.A1(_00679_),
    .A2(net17212),
    .B(_00680_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24665_ (.A1(_00678_),
    .A2(_00681_),
    .A3(net20011),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24666_ (.A1(_00682_),
    .A2(_00677_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24667_ (.I(_15406_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24668_ (.A1(_15426_),
    .A2(_00684_),
    .B(net20009),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24669_ (.I(_15203_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24670_ (.A1(_00564_),
    .A2(net19765),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24671_ (.A1(_15472_),
    .A2(_00686_),
    .B(_00687_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24672_ (.A1(_00685_),
    .A2(_00688_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24673_ (.A1(net17507),
    .A2(net18734),
    .B(net19747),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24674_ (.A1(_00679_),
    .A2(_00690_),
    .B(net19742),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24675_ (.A1(net17293),
    .A2(net17296),
    .A3(net18716),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24676_ (.A1(_15177_),
    .A2(net17508),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24677_ (.A1(_00692_),
    .A2(_00693_),
    .A3(net19747),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24678_ (.A1(_00694_),
    .A2(_00691_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24679_ (.A1(_00695_),
    .A2(_00689_),
    .A3(net20430),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24680_ (.A1(_00683_),
    .A2(_00696_),
    .A3(net20631),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24681_ (.A1(_00671_),
    .A2(_00697_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24682_ (.A1(_15123_),
    .A2(net454),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _24683_ (.A1(_00698_),
    .A2(net18708),
    .A3(_15254_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24684_ (.A1(_00699_),
    .A2(_15258_),
    .A3(_00591_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24685_ (.A1(_15386_),
    .A2(_15383_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24686_ (.A1(_15345_),
    .A2(net18708),
    .A3(net17300),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24687_ (.A1(_00701_),
    .A2(_00702_),
    .A3(_15272_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24688_ (.A1(_00703_),
    .A2(net19764),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24689_ (.A1(_00700_),
    .A2(_00704_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24690_ (.A1(_00705_),
    .A2(net20010),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24691_ (.A1(net17510),
    .A2(net17289),
    .B(net18725),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24692_ (.A1(_00605_),
    .A2(_00707_),
    .B(net20009),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24693_ (.A1(_15531_),
    .A2(net17831),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24694_ (.A1(_15884_[0]),
    .A2(_15893_[0]),
    .B(net18723),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24695_ (.A1(_00709_),
    .A2(net19758),
    .A3(_00710_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24696_ (.A1(_00708_),
    .A2(_00711_),
    .B(net20429),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24697_ (.A1(_00706_),
    .A2(_00712_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24698_ (.A1(_15330_),
    .A2(net18712),
    .A3(net17309),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24699_ (.A1(_00714_),
    .A2(net19754),
    .A3(_15492_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24700_ (.A1(_15330_),
    .A2(net18735),
    .A3(_15350_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24701_ (.A1(_00611_),
    .A2(net17293),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24702_ (.A1(_00716_),
    .A2(_00717_),
    .A3(net19767),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24703_ (.A1(_00715_),
    .A2(_00718_),
    .A3(net19742),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24704_ (.A1(net17833),
    .A2(_15398_),
    .A3(net18736),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24705_ (.A1(_15303_),
    .A2(net19747),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24706_ (.A1(_00720_),
    .A2(_00721_),
    .B(net19742),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24707_ (.A1(_15416_),
    .A2(_00563_),
    .B(net19747),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24708_ (.A1(net17840),
    .A2(net18731),
    .A3(net18704),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24709_ (.A1(_00723_),
    .A2(_00724_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24710_ (.A1(_00722_),
    .A2(_00725_),
    .B(net20233),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24711_ (.A1(_00719_),
    .A2(_00726_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24712_ (.A1(_00713_),
    .A2(net20427),
    .A3(_00727_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24713_ (.I(_15275_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24714_ (.A1(_00589_),
    .A2(_00729_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24715_ (.A1(_00730_),
    .A2(net19751),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24716_ (.A1(_15467_),
    .A2(net19760),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24717_ (.A1(_00731_),
    .A2(_00732_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24718_ (.A1(_00733_),
    .A2(net20010),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24719_ (.A1(_15406_),
    .A2(net17293),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24720_ (.A1(_00735_),
    .A2(net19747),
    .A3(_15362_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24721_ (.I(_15885_[0]),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24722_ (.A1(_00737_),
    .A2(net18724),
    .B(net19747),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24723_ (.A1(_00738_),
    .A2(_00675_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24724_ (.A1(_00736_),
    .A2(_00739_),
    .A3(net19743),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24725_ (.A1(_00734_),
    .A2(net20429),
    .A3(_00740_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24726_ (.A1(net19768),
    .A2(net17600),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24727_ (.A1(net18195),
    .A2(_00742_),
    .B(net18708),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24728_ (.A1(_15320_),
    .A2(net18726),
    .A3(net18705),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24729_ (.A1(_00743_),
    .A2(_00744_),
    .A3(net19755),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24730_ (.A1(net18201),
    .A2(net18708),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24731_ (.A1(_00550_),
    .A2(_00746_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24732_ (.A1(_00745_),
    .A2(_00747_),
    .A3(net19742),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24733_ (.A1(_15398_),
    .A2(net18727),
    .B(net19759),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24734_ (.A1(_00749_),
    .A2(_15335_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24735_ (.A1(net17506),
    .A2(net18715),
    .B(net19747),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24736_ (.A1(_00582_),
    .A2(_00751_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24737_ (.A1(_00750_),
    .A2(_00752_),
    .A3(net20010),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24738_ (.A1(_00748_),
    .A2(net20231),
    .A3(_00753_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24739_ (.A1(_00741_),
    .A2(_00754_),
    .A3(net20631),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24740_ (.A1(_00728_),
    .A2(_00755_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24741_ (.A1(_15255_),
    .A2(net19759),
    .A3(net17301),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24742_ (.A1(net18197),
    .A2(net18202),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24743_ (.A1(_00756_),
    .A2(_00757_),
    .B(net19742),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24744_ (.A1(net18723),
    .A2(net17602),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24745_ (.A1(_00709_),
    .A2(net19747),
    .A3(_00759_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24746_ (.A1(_00758_),
    .A2(_00760_),
    .B(net20429),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _24747_ (.A1(_15299_),
    .A2(net17515),
    .A3(net18716),
    .B1(net17505),
    .B2(net18196),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24748_ (.A1(_00762_),
    .A2(_15486_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _24749_ (.A1(net17201),
    .A2(net17213),
    .B1(net18715),
    .B2(net18196),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24750_ (.A1(_00746_),
    .A2(net19747),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24751_ (.A1(_00764_),
    .A2(_00765_),
    .B(net20009),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24752_ (.A1(_00763_),
    .A2(_00766_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24753_ (.A1(_00761_),
    .A2(_00767_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24754_ (.A1(_15291_),
    .A2(net17294),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24755_ (.A1(net18199),
    .A2(_15450_),
    .B(net19749),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24756_ (.A1(_15515_),
    .A2(net17290),
    .B(net18723),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24757_ (.A1(_15893_[0]),
    .A2(net18724),
    .B(net19747),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24758_ (.A1(_00771_),
    .A2(_00772_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _24759_ (.A1(_00769_),
    .A2(_00770_),
    .B(_00773_),
    .C(net20009),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24760_ (.A1(_00593_),
    .A2(net18725),
    .B(net19747),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24761_ (.A1(_00775_),
    .A2(_15255_),
    .B(net20009),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24762_ (.A1(_15357_),
    .A2(_00765_),
    .A3(_00591_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24763_ (.A1(_00776_),
    .A2(_00777_),
    .B(net20231),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24764_ (.A1(_00774_),
    .A2(_00778_),
    .B(net20631),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24765_ (.A1(_00768_),
    .A2(_00779_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24766_ (.A1(_15367_),
    .A2(net17841),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24767_ (.A1(_15512_),
    .A2(_00781_),
    .A3(_00701_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24768_ (.A1(_15371_),
    .A2(net19747),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24769_ (.A1(_00783_),
    .A2(_00589_),
    .B(net20429),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24770_ (.A1(_00782_),
    .A2(_00784_),
    .B(net20010),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24771_ (.A1(_15315_),
    .A2(net18721),
    .A3(net17829),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24772_ (.A1(_00786_),
    .A2(net19761),
    .A3(_15500_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24773_ (.A1(net18722),
    .A2(net19209),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _24774_ (.A1(_00633_),
    .A2(net18722),
    .B(net19750),
    .C(_00788_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24775_ (.A1(_00787_),
    .A2(_00789_),
    .A3(net20429),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24776_ (.A1(_00785_),
    .A2(_00790_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24777_ (.A1(_15291_),
    .A2(net17295),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24778_ (.A1(_00562_),
    .A2(_00792_),
    .A3(net19750),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24779_ (.A1(_15507_),
    .A2(net19764),
    .A3(_00702_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24780_ (.A1(_00793_),
    .A2(_00794_),
    .A3(net20231),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24781_ (.A1(_15300_),
    .A2(net19759),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24782_ (.A1(_00796_),
    .A2(_15384_),
    .B(_15239_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24783_ (.A1(net17841),
    .A2(net18728),
    .B(net19759),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24784_ (.A1(_15315_),
    .A2(net18715),
    .A3(net17294),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24785_ (.A1(_00798_),
    .A2(_00799_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24786_ (.A1(_00797_),
    .A2(_00800_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24787_ (.A1(_00795_),
    .A2(_00801_),
    .A3(net20010),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24788_ (.A1(_00791_),
    .A2(_00802_),
    .A3(net20631),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24789_ (.A1(_00780_),
    .A2(_00803_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24790_ (.I(\sa21_sub[7] ),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24791_ (.A1(_00804_),
    .A2(_12815_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24792_ (.A1(net21330),
    .A2(net21314),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24793_ (.A1(_00806_),
    .A2(_00805_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24794_ (.A1(_00807_),
    .A2(_12770_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24795_ (.A1(_00804_),
    .A2(\sa21_sub[0] ),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24796_ (.A1(_12815_),
    .A2(net21314),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24797_ (.A1(_00810_),
    .A2(_00809_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24798_ (.A1(net20878),
    .A2(_12777_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24799_ (.A1(_00812_),
    .A2(_00808_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24800_ (.A1(_12785_),
    .A2(\sa03_sr[1] ),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24801_ (.A1(_12789_),
    .A2(_12830_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24802_ (.A1(_00814_),
    .A2(_00815_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24803_ (.A1(_00816_),
    .A2(_00813_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24804_ (.A1(_12777_),
    .A2(net20878),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24805_ (.A1(_12770_),
    .A2(net20880),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24806_ (.A1(_00819_),
    .A2(_00818_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24807_ (.A1(_12785_),
    .A2(_12830_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24808_ (.A1(_12789_),
    .A2(\sa03_sr[1] ),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24809_ (.A1(_00821_),
    .A2(_00822_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24810_ (.A1(_00820_),
    .A2(_00823_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24811_ (.A1(_00824_),
    .A2(_00817_),
    .A3(_10378_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24812_ (.A1(net21486),
    .A2(\text_in_r[17] ),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24813_ (.A1(_00825_),
    .A2(_00826_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24814_ (.I(net21150),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24815_ (.A1(_00828_),
    .A2(net20008),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24816_ (.A1(net20230),
    .A2(net21150),
    .A3(net20973),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24817_ (.A1(_00829_),
    .A2(_00830_),
    .ZN(_15903_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24818_ (.A1(net21005),
    .A2(net21272),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24819_ (.A1(net21002),
    .A2(net21375),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24820_ (.A1(_00831_),
    .A2(_00832_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24821_ (.A1(_00833_),
    .A2(net21443),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24822_ (.A1(_00831_),
    .A2(_00832_),
    .A3(net21010),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24823_ (.A1(_00834_),
    .A2(_00835_),
    .A3(net20879),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24824_ (.A1(net21443),
    .A2(net21375),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24825_ (.I(_00837_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24826_ (.A1(net21443),
    .A2(net21375),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24827_ (.A1(_00838_),
    .A2(_00839_),
    .B(net21272),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24828_ (.A1(net21010),
    .A2(net21005),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24829_ (.A1(_00841_),
    .A2(net21002),
    .A3(_00837_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24830_ (.A1(_00840_),
    .A2(net20881),
    .A3(_00842_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _24831_ (.A1(_00836_),
    .A2(_00843_),
    .B(net21486),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24832_ (.I(\text_in_r[16] ),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24833_ (.A1(_00845_),
    .A2(net21486),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24834_ (.A1(net20426),
    .A2(_00846_),
    .B(net21151),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24835_ (.A1(_00836_),
    .A2(_00843_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24836_ (.A1(_00848_),
    .A2(net21089),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24837_ (.I(net21151),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24838_ (.I(_00846_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24839_ (.A1(net20229),
    .A2(_00850_),
    .A3(_00851_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24840_ (.A1(_00852_),
    .A2(_00847_),
    .ZN(_15906_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24841_ (.A1(net21325),
    .A2(net21268),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24842_ (.A1(net21325),
    .A2(net21268),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24843_ (.A1(_00853_),
    .A2(_00854_),
    .B(net21440),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24844_ (.A1(_12834_),
    .A2(net20998),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24845_ (.A1(net21325),
    .A2(net21268),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24846_ (.A1(_00856_),
    .A2(net20994),
    .A3(_00857_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24847_ (.A1(_00855_),
    .A2(_00858_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24848_ (.A1(net21382),
    .A2(net21328),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24849_ (.I(_00860_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24850_ (.A1(_00859_),
    .A2(_00861_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24851_ (.A1(_00855_),
    .A2(_00858_),
    .A3(_00860_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24852_ (.A1(_00862_),
    .A2(_00863_),
    .B(net21486),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24853_ (.I(\text_in_r[18] ),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24854_ (.A1(_00865_),
    .A2(net21486),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24855_ (.I(net21149),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24856_ (.A1(_00864_),
    .A2(_00866_),
    .B(_00867_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24857_ (.A1(_00862_),
    .A2(_00863_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24858_ (.A1(_00869_),
    .A2(net21089),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24859_ (.I(_00866_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24860_ (.A1(_00870_),
    .A2(net21149),
    .A3(_00871_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24861_ (.A1(_00868_),
    .A2(_00872_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output358 (.I(net358),
    .Z(text_out[73]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24863_ (.A1(_00844_),
    .A2(_00846_),
    .B(_00850_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24864_ (.A1(_00849_),
    .A2(net21151),
    .A3(_00851_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24865_ (.A1(_00875_),
    .A2(_00874_),
    .ZN(_15897_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24866_ (.A1(_00864_),
    .A2(_00866_),
    .B(net21149),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24867_ (.A1(_00870_),
    .A2(_00867_),
    .A3(_00871_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24868_ (.A1(_00876_),
    .A2(_00877_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output357 (.I(net357),
    .Z(text_out[72]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24870_ (.A1(_12834_),
    .A2(net20974),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24871_ (.A1(net21325),
    .A2(net21315),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24872_ (.A1(_00879_),
    .A2(_00880_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24873_ (.A1(_12872_),
    .A2(_00881_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24874_ (.A1(net20974),
    .A2(net21325),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24875_ (.A1(_12834_),
    .A2(net21315),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24876_ (.A1(_00883_),
    .A2(_00884_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24877_ (.A1(_12879_),
    .A2(_00885_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24878_ (.A1(_00882_),
    .A2(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24879_ (.I(_00887_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24880_ (.A1(_12898_),
    .A2(net21439),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24881_ (.I(\sa03_sr[3] ),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24882_ (.A1(_12896_),
    .A2(net20972),
    .A3(_12897_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24883_ (.A1(_00889_),
    .A2(_00891_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24884_ (.I(_00892_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24885_ (.A1(_00888_),
    .A2(_00893_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24886_ (.A1(_00887_),
    .A2(_00892_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24887_ (.A1(_00894_),
    .A2(net21094),
    .A3(_00895_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24888_ (.A1(net21486),
    .A2(\text_in_r[19] ),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24889_ (.A1(_00896_),
    .A2(_00897_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24890_ (.A1(_00898_),
    .A2(net21148),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24891_ (.I(net21148),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24892_ (.A1(_00896_),
    .A2(_00900_),
    .A3(_00897_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24893_ (.A1(_00899_),
    .A2(_00901_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output356 (.I(net356),
    .Z(text_out[71]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output355 (.I(net355),
    .Z(text_out[70]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24896_ (.I(_15900_[0]),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24897_ (.A1(net20228),
    .A2(_00905_),
    .A3(net20007),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24898_ (.I(_00906_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24899_ (.A1(net19739),
    .A2(net18394),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output354 (.I(net354),
    .Z(text_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24901_ (.A1(net19731),
    .A2(net18393),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24902_ (.A1(_00908_),
    .A2(_00910_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output353 (.I(net353),
    .Z(text_out[69]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24904_ (.A1(_00911_),
    .A2(net18689),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24905_ (.A1(_12870_),
    .A2(net20974),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24906_ (.A1(net21322),
    .A2(net21315),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24907_ (.A1(_00914_),
    .A2(_00915_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24908_ (.I(_00916_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24909_ (.I(\sa32_sub[4] ),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24910_ (.A1(_12928_),
    .A2(_00918_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24911_ (.A1(\sa21_sub[4] ),
    .A2(\sa32_sub[4] ),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24912_ (.A1(_00919_),
    .A2(_00920_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24913_ (.A1(_00917_),
    .A2(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24914_ (.I(_00921_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24915_ (.A1(_00923_),
    .A2(_00916_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24916_ (.A1(_00922_),
    .A2(_00924_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24917_ (.I(_00925_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24918_ (.A1(net21437),
    .A2(_12889_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24919_ (.A1(_00926_),
    .A2(_00927_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24920_ (.A1(_12889_),
    .A2(net21437),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24921_ (.A1(_12889_),
    .A2(net21437),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24922_ (.A1(_00929_),
    .A2(_00930_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24923_ (.A1(_00925_),
    .A2(_00931_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24924_ (.A1(_00928_),
    .A2(_00932_),
    .A3(net21094),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24925_ (.A1(net21486),
    .A2(\text_in_r[20] ),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24926_ (.A1(_00933_),
    .A2(_00934_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24927_ (.A1(_00935_),
    .A2(net21146),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24928_ (.I(net21146),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24929_ (.A1(_00933_),
    .A2(_00937_),
    .A3(_00934_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24930_ (.A1(_00936_),
    .A2(_00938_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _24931_ (.I(_00939_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output352 (.I(net352),
    .Z(text_out[68]));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _24933_ (.A1(net18691),
    .A2(net17503),
    .B(_00913_),
    .C(net17819),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24934_ (.A1(net19205),
    .A2(net19741),
    .A3(net19731),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24935_ (.A1(_00898_),
    .A2(_00900_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24936_ (.A1(_00896_),
    .A2(net21148),
    .A3(_00897_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24937_ (.A1(_00944_),
    .A2(_00945_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output351 (.I(net351),
    .Z(text_out[67]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24939_ (.A1(net19739),
    .A2(net19736),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24940_ (.A1(net18682),
    .A2(net18675),
    .A3(net19203),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24941_ (.I(_00908_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output350 (.I(net350),
    .Z(text_out[66]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output349 (.I(net349),
    .Z(text_out[65]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output348 (.I(net348),
    .Z(text_out[64]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24945_ (.A1(net17813),
    .A2(net18691),
    .B(net17819),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24946_ (.A1(_00949_),
    .A2(_00954_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24947_ (.I(\sa03_sr[5] ),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24948_ (.A1(_00956_),
    .A2(_12958_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24949_ (.A1(net21378),
    .A2(net21320),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24950_ (.I(_00958_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24951_ (.A1(_00957_),
    .A2(_00959_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24952_ (.A1(_00957_),
    .A2(_00959_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24953_ (.A1(_00960_),
    .A2(_00961_),
    .A3(net21092),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24954_ (.A1(net21489),
    .A2(\text_in_r[21] ),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24955_ (.A1(_00962_),
    .A2(_00963_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24956_ (.A1(_00964_),
    .A2(\u0.tmp_w[21] ),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24957_ (.I(\u0.tmp_w[21] ),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24958_ (.A1(_00962_),
    .A2(_00966_),
    .A3(_00963_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24959_ (.A1(_00965_),
    .A2(_00967_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output347 (.I(net347),
    .Z(text_out[63]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24961_ (.A1(_00955_),
    .A2(_00942_),
    .A3(net20000),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24962_ (.A1(net19731),
    .A2(net18395),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _24963_ (.I(_00971_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24964_ (.I(_15899_[0]),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24965_ (.A1(net19739),
    .A2(net18180),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24966_ (.A1(_00972_),
    .A2(_00974_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output346 (.I(net346),
    .Z(text_out[62]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24968_ (.A1(_00975_),
    .A2(net18693),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24969_ (.I(_15904_[0]),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24970_ (.A1(net19731),
    .A2(_00978_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output345 (.I(net345),
    .Z(text_out[61]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24972_ (.A1(_00979_),
    .A2(net18670),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output344 (.I(net344),
    .Z(text_out[60]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output343 (.I(net343),
    .Z(text_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _24975_ (.A1(net17501),
    .A2(net18188),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output342 (.I(net342),
    .Z(text_out[59]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24977_ (.A1(_00984_),
    .A2(_00977_),
    .B(net20002),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24978_ (.A1(net19731),
    .A2(net19741),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _24979_ (.I(_00987_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _24980_ (.I(_15907_[0]),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _24981_ (.A1(net19739),
    .A2(_00989_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output341 (.I(net341),
    .Z(text_out[58]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output340 (.I(net340),
    .Z(text_out[57]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _24984_ (.A1(net18669),
    .A2(net17811),
    .B(net18673),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24985_ (.A1(net19204),
    .A2(net19731),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24986_ (.A1(net18397),
    .A2(net20006),
    .A3(net20227),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _24987_ (.A1(_00994_),
    .A2(net18178),
    .A3(net18701),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output339 (.I(net339),
    .Z(text_out[56]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _24989_ (.A1(_00993_),
    .A2(_00996_),
    .A3(net18188),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24990_ (.A1(net21377),
    .A2(net21318),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24991_ (.I(\sa03_sr[6] ),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _24992_ (.A1(_01000_),
    .A2(_13007_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _24993_ (.A1(_00999_),
    .A2(_01001_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _24994_ (.A1(net21489),
    .A2(\text_in_r[22] ),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _24995_ (.A1(_01002_),
    .A2(net21092),
    .B(_01003_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _24996_ (.I(\u0.tmp_w[22] ),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _24997_ (.A1(_01004_),
    .A2(_01005_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _24998_ (.A1(_01004_),
    .A2(_01005_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _24999_ (.A1(_01006_),
    .A2(_01007_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output338 (.I(net338),
    .Z(text_out[55]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25001_ (.A1(_00986_),
    .A2(_00998_),
    .B(net20222),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25002_ (.A1(_01010_),
    .A2(_00970_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25003_ (.A1(net21435),
    .A2(net21376),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25004_ (.A1(net21316),
    .A2(_01012_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _25005_ (.A1(net21315),
    .A2(net21258),
    .A3(_01013_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _25006_ (.I0(_01014_),
    .I1(\text_in_r[23] ),
    .S(net21489),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _25007_ (.A1(\u0.tmp_w[23] ),
    .A2(_01015_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output337 (.I(net337),
    .Z(text_out[54]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _25009_ (.I(_01016_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25010_ (.A1(net19739),
    .A2(net19741),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25011_ (.A1(net19731),
    .A2(_00973_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25012_ (.A1(_01019_),
    .A2(_01020_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output336 (.I(net336),
    .Z(text_out[53]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25014_ (.A1(_01021_),
    .A2(net18673),
    .B(net17820),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25015_ (.A1(net19205),
    .A2(net19737),
    .A3(net19731),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25016_ (.A1(net20227),
    .A2(net20006),
    .A3(_00978_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25017_ (.A1(_01024_),
    .A2(net18694),
    .A3(_01025_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25018_ (.A1(net20227),
    .A2(net20006),
    .A3(net18395),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25019_ (.I(_01027_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25020_ (.A1(net18685),
    .A2(_01028_),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25021_ (.A1(_01023_),
    .A2(_01026_),
    .A3(net17499),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25022_ (.I(_00995_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25023_ (.A1(_01031_),
    .A2(net18694),
    .B(net18189),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25024_ (.A1(net18679),
    .A2(_15920_[0]),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25025_ (.I(_00968_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output335 (.I(net335),
    .Z(text_out[52]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25027_ (.A1(_01032_),
    .A2(_01033_),
    .B(net19725),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25028_ (.A1(_01030_),
    .A2(_01036_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25029_ (.A1(_00971_),
    .A2(net18693),
    .B(net17819),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25030_ (.I(_15909_[0]),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25031_ (.A1(_01039_),
    .A2(net20006),
    .A3(net20227),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25032_ (.A1(_01040_),
    .A2(net18670),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25033_ (.A1(_01041_),
    .A2(net18668),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output334 (.I(net334),
    .Z(text_out[51]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25035_ (.A1(_01038_),
    .A2(_01042_),
    .B(net20002),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25036_ (.A1(net19739),
    .A2(_15907_[0]),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25037_ (.A1(_01045_),
    .A2(net18684),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25038_ (.A1(net17803),
    .A2(net18667),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output333 (.I(net333),
    .Z(text_out[50]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25040_ (.A1(_00971_),
    .A2(net18672),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25041_ (.A1(_01047_),
    .A2(net17819),
    .A3(_01049_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25042_ (.A1(_01044_),
    .A2(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output332 (.I(net332),
    .Z(text_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25044_ (.A1(_01037_),
    .A2(_01051_),
    .A3(net20225),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25045_ (.A1(net20424),
    .A2(_01011_),
    .A3(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25046_ (.A1(_00948_),
    .A2(net18684),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25047_ (.A1(net18175),
    .A2(net18193),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25048_ (.A1(net19205),
    .A2(net19738),
    .A3(net19739),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25049_ (.A1(net17501),
    .A2(net18665),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25050_ (.A1(_01056_),
    .A2(_01058_),
    .B(net20002),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25051_ (.A1(net19731),
    .A2(net19736),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25052_ (.A1(net18665),
    .A2(net18691),
    .A3(_01060_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25053_ (.A1(net18670),
    .A2(_00906_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _25054_ (.I(_15913_[0]),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25055_ (.A1(_01063_),
    .A2(net19739),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25056_ (.A1(net17497),
    .A2(net17802),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output331 (.I(net331),
    .Z(text_out[49]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25058_ (.A1(_01061_),
    .A2(_01065_),
    .A3(net17819),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25059_ (.A1(_01059_),
    .A2(_01067_),
    .B(net20222),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25060_ (.A1(_01057_),
    .A2(net18691),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25061_ (.A1(net21150),
    .A2(_00827_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25062_ (.A1(_00825_),
    .A2(_00828_),
    .A3(_00826_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25063_ (.A1(_01070_),
    .A2(_01071_),
    .ZN(_15898_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25064_ (.A1(net19198),
    .A2(net19731),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25065_ (.I(_01072_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25066_ (.A1(_01069_),
    .A2(_01073_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25067_ (.A1(_00948_),
    .A2(net18676),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25068_ (.A1(net19731),
    .A2(_01063_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output330 (.I(net330),
    .Z(text_out[48]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25070_ (.A1(_01075_),
    .A2(net17800),
    .B(net18189),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25071_ (.A1(_01074_),
    .A2(_01078_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25072_ (.A1(net19206),
    .A2(net19732),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25073_ (.A1(_01080_),
    .A2(net18183),
    .B(net18691),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output329 (.I(net329),
    .Z(text_out[47]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25075_ (.A1(_00949_),
    .A2(_01081_),
    .A3(net18188),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output328 (.I(net328),
    .Z(text_out[46]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25077_ (.A1(_01079_),
    .A2(_01083_),
    .A3(net20002),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25078_ (.A1(_01085_),
    .A2(_01068_),
    .B(_01018_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _25079_ (.I(_01020_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output327 (.I(net327),
    .Z(text_out[45]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25081_ (.A1(_00990_),
    .A2(net17494),
    .B(net18695),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25082_ (.A1(net19740),
    .A2(net18398),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25083_ (.A1(net17496),
    .A2(net18172),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25084_ (.A1(_01089_),
    .A2(_01091_),
    .B(net17823),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25085_ (.A1(net19739),
    .A2(net453),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25086_ (.A1(net18670),
    .A2(_01093_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25087_ (.A1(_01094_),
    .A2(net18189),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25088_ (.A1(net18396),
    .A2(net20007),
    .A3(net20228),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25089_ (.A1(_01096_),
    .A2(net18684),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25090_ (.I(_01097_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25091_ (.A1(net19205),
    .A2(net19739),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25092_ (.A1(_01098_),
    .A2(net18659),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25093_ (.A1(_01095_),
    .A2(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25094_ (.A1(_01092_),
    .A2(_01101_),
    .B(net20002),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25095_ (.A1(_00987_),
    .A2(net18684),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25096_ (.A1(net19199),
    .A2(net19736),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25097_ (.A1(_01103_),
    .A2(net18658),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25098_ (.A1(net19738),
    .A2(net427),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25099_ (.A1(_01106_),
    .A2(net18680),
    .A3(net19200),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25100_ (.A1(_01105_),
    .A2(net17819),
    .A3(_01107_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25101_ (.A1(net17827),
    .A2(net18691),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25102_ (.A1(net19205),
    .A2(net19741),
    .A3(net19739),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25103_ (.A1(_01109_),
    .A2(net18656),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25104_ (.A1(net19734),
    .A2(_00989_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25105_ (.A1(_00974_),
    .A2(net17798),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25106_ (.A1(_01113_),
    .A2(net18673),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25107_ (.A1(_01111_),
    .A2(_01114_),
    .A3(net18188),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output326 (.I(net326),
    .Z(text_out[44]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25109_ (.A1(_01108_),
    .A2(_01115_),
    .A3(net19729),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25110_ (.A1(_01102_),
    .A2(net20225),
    .A3(_01117_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25111_ (.A1(_01118_),
    .A2(_01086_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25112_ (.A1(_01054_),
    .A2(_01119_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25113_ (.A1(net19199),
    .A2(net19739),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25114_ (.A1(_00981_),
    .A2(_01120_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25115_ (.A1(net19201),
    .A2(_01090_),
    .A3(net18694),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25116_ (.A1(_01121_),
    .A2(net18194),
    .A3(_01122_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25117_ (.A1(net390),
    .A2(net18694),
    .B(net18189),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25118_ (.I(_01019_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25119_ (.A1(_01125_),
    .A2(net18699),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25120_ (.A1(_01020_),
    .A2(net18178),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output325 (.I(net325),
    .Z(text_out[43]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25122_ (.A1(_01127_),
    .A2(net18680),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25123_ (.A1(_01129_),
    .A2(_01126_),
    .A3(_01124_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25124_ (.A1(_01123_),
    .A2(_01130_),
    .A3(net19728),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25125_ (.A1(_01110_),
    .A2(net18676),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _25126_ (.I(_01096_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _25127_ (.A1(_01132_),
    .A2(_01133_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25128_ (.A1(net18684),
    .A2(_01076_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25129_ (.I(_15901_[0]),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25130_ (.A1(net19739),
    .A2(net18168),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25131_ (.A1(_01135_),
    .A2(_01137_),
    .B(net18189),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25132_ (.A1(_01134_),
    .A2(_01138_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _25133_ (.I(_01055_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25134_ (.A1(_01140_),
    .A2(net18682),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25135_ (.A1(_01062_),
    .A2(net17820),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25136_ (.A1(_01142_),
    .A2(_01141_),
    .B(net19725),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25137_ (.A1(_01139_),
    .A2(_01143_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25138_ (.A1(_01131_),
    .A2(_01144_),
    .B(net20222),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25139_ (.A1(_01103_),
    .A2(net18659),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25140_ (.A1(_01146_),
    .A2(_01121_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25141_ (.A1(_01147_),
    .A2(net20002),
    .B(net18194),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25142_ (.A1(net18682),
    .A2(net18665),
    .A3(net18673),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25143_ (.A1(_01060_),
    .A2(_01090_),
    .A3(net18694),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25144_ (.A1(_01149_),
    .A2(_01150_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25145_ (.A1(_01151_),
    .A2(net19728),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25146_ (.I(_15923_[0]),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25147_ (.A1(net18676),
    .A2(_01153_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25148_ (.A1(_01154_),
    .A2(net20000),
    .B(_00940_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25149_ (.A1(_01046_),
    .A2(_00943_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25150_ (.A1(_01155_),
    .A2(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25151_ (.A1(_01157_),
    .A2(net20222),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25152_ (.A1(_01148_),
    .A2(_01152_),
    .B(_01158_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25153_ (.A1(_01159_),
    .A2(_01145_),
    .B(net20630),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25154_ (.A1(net19731),
    .A2(net18394),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output324 (.I(net324),
    .Z(text_out[42]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25156_ (.A1(_01161_),
    .A2(net18701),
    .B(net17820),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25157_ (.A1(_01134_),
    .A2(_01163_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25158_ (.A1(_01064_),
    .A2(net18670),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _25159_ (.A1(_01165_),
    .A2(_01073_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25160_ (.A1(net426),
    .A2(net19741),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25161_ (.A1(_01167_),
    .A2(net19731),
    .A3(net18699),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25162_ (.A1(_01166_),
    .A2(_01168_),
    .A3(net17820),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25163_ (.A1(_01164_),
    .A2(_01169_),
    .A3(net19727),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25164_ (.A1(net17813),
    .A2(net17502),
    .B(net18672),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25165_ (.A1(_01021_),
    .A2(net18694),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25166_ (.A1(_01171_),
    .A2(_01172_),
    .A3(net17820),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25167_ (.A1(_01167_),
    .A2(_01060_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25168_ (.A1(_01174_),
    .A2(net18674),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25169_ (.A1(_00995_),
    .A2(net18694),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25170_ (.A1(_01176_),
    .A2(_01060_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25171_ (.A1(_01175_),
    .A2(_01177_),
    .A3(net18192),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25172_ (.A1(_01173_),
    .A2(_01178_),
    .A3(net20002),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _25173_ (.I(_01008_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output323 (.I(net323),
    .Z(text_out[41]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25175_ (.A1(_01170_),
    .A2(_01179_),
    .A3(_01180_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25176_ (.A1(_01094_),
    .A2(net17800),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25177_ (.A1(_01026_),
    .A2(_01183_),
    .A3(net18188),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _25178_ (.A1(_00950_),
    .A2(net18688),
    .B(net18186),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25179_ (.A1(_01099_),
    .A2(net18670),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25180_ (.A1(_01185_),
    .A2(net18663),
    .A3(net18166),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25181_ (.A1(_01184_),
    .A2(net20002),
    .A3(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25182_ (.A1(_00979_),
    .A2(net18684),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25183_ (.A1(_01189_),
    .A2(_01125_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25184_ (.A1(_01062_),
    .A2(net19203),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25185_ (.A1(_01191_),
    .A2(net17820),
    .A3(_01190_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25186_ (.A1(_00994_),
    .A2(_01104_),
    .A3(net18701),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25187_ (.A1(net18670),
    .A2(net19740),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25188_ (.A1(_01194_),
    .A2(_01106_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25189_ (.A1(_01193_),
    .A2(_01195_),
    .A3(net18192),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25190_ (.A1(net19725),
    .A2(_01196_),
    .A3(_01192_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25191_ (.A1(_01188_),
    .A2(net20222),
    .A3(_01197_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25192_ (.A1(_01182_),
    .A2(_01198_),
    .A3(_01018_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25193_ (.A1(_01160_),
    .A2(_01199_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25194_ (.A1(_01060_),
    .A2(net17806),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25195_ (.A1(_01200_),
    .A2(net18672),
    .A3(net18661),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25196_ (.A1(_01201_),
    .A2(_00996_),
    .A3(net18188),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25197_ (.A1(_00994_),
    .A2(net428),
    .A3(net18674),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25198_ (.A1(net17812),
    .A2(_01064_),
    .A3(net18690),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25199_ (.A1(_01203_),
    .A2(_01204_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25200_ (.A1(_01205_),
    .A2(net17819),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25201_ (.A1(_01202_),
    .A2(_01206_),
    .A3(net20001),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25202_ (.A1(net18664),
    .A2(net18697),
    .B(net17817),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25203_ (.A1(net18655),
    .A2(net18679),
    .A3(net17800),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25204_ (.A1(_01208_),
    .A2(_01209_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25205_ (.A1(_01097_),
    .A2(_01080_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25206_ (.A1(_01027_),
    .A2(net18670),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25207_ (.A1(_01212_),
    .A2(_00988_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25208_ (.A1(_01211_),
    .A2(_01213_),
    .B(net17819),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25209_ (.A1(_01210_),
    .A2(_01214_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25210_ (.A1(_01215_),
    .A2(net19726),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25211_ (.A1(_01207_),
    .A2(_01216_),
    .A3(net20223),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25212_ (.A1(net20227),
    .A2(net20006),
    .A3(net18392),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25213_ (.A1(_00987_),
    .A2(_01218_),
    .A3(net18684),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25214_ (.A1(_01219_),
    .A2(net17814),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25215_ (.A1(_00910_),
    .A2(net18671),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25216_ (.A1(_01221_),
    .A2(_01080_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25217_ (.A1(_01220_),
    .A2(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25218_ (.A1(_01060_),
    .A2(net17804),
    .A3(net18686),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25219_ (.A1(_00906_),
    .A2(net18177),
    .A3(net18671),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25220_ (.A1(_01225_),
    .A2(_01224_),
    .B(net17814),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25221_ (.A1(_01223_),
    .A2(_01226_),
    .B(net19725),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25222_ (.A1(net18661),
    .A2(net18672),
    .A3(net17806),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25223_ (.A1(_00913_),
    .A2(_01228_),
    .A3(net18187),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25224_ (.I(_01218_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25225_ (.A1(_01230_),
    .A2(net18687),
    .B(net18184),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25226_ (.I(_00910_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25227_ (.A1(_01232_),
    .A2(net18686),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25228_ (.A1(_01060_),
    .A2(_01025_),
    .A3(net18670),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25229_ (.A1(_01231_),
    .A2(_01233_),
    .A3(_01234_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25230_ (.A1(_01229_),
    .A2(_01235_),
    .A3(net20000),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25231_ (.A1(_01227_),
    .A2(_01236_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25232_ (.A1(_01237_),
    .A2(_01180_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25233_ (.A1(_01217_),
    .A2(_01238_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25234_ (.A1(_01239_),
    .A2(net20630),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output322 (.I(net322),
    .Z(text_out[40]));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _25236_ (.A1(net18684),
    .A2(_15918_[0]),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25237_ (.A1(_01069_),
    .A2(_01242_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25238_ (.A1(_15927_[0]),
    .A2(net18697),
    .B(net18189),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25239_ (.A1(_01203_),
    .A2(_01244_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25240_ (.A1(net17819),
    .A2(net17792),
    .B(_01245_),
    .C(net20001),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25241_ (.A1(_01087_),
    .A2(net18698),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25242_ (.A1(_01247_),
    .A2(net18191),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25243_ (.A1(net17807),
    .A2(net17495),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25244_ (.A1(_01249_),
    .A2(_01248_),
    .B(net20004),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25245_ (.A1(net18676),
    .A2(net19731),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25246_ (.I(_01251_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25247_ (.A1(_01136_),
    .A2(_00978_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25248_ (.I(net17790),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25249_ (.A1(net17791),
    .A2(_01254_),
    .B(net18189),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25250_ (.A1(_01120_),
    .A2(_00948_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25251_ (.A1(_01256_),
    .A2(net18674),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25252_ (.A1(_01255_),
    .A2(net17491),
    .A3(_01257_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25253_ (.A1(_01250_),
    .A2(_01258_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25254_ (.A1(_01246_),
    .A2(net20222),
    .A3(_01259_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25255_ (.A1(_15920_[0]),
    .A2(net18697),
    .B(net17817),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25256_ (.A1(net17493),
    .A2(net18666),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25257_ (.A1(_01261_),
    .A2(_01262_),
    .B(net20003),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25258_ (.A1(_01120_),
    .A2(net18676),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25259_ (.A1(_01264_),
    .A2(_01060_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25260_ (.A1(_01265_),
    .A2(net17820),
    .A3(_00996_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25261_ (.A1(_01263_),
    .A2(_01266_),
    .B(net20224),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25262_ (.A1(_01104_),
    .A2(net18676),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25263_ (.A1(_01268_),
    .A2(_00994_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25264_ (.A1(net18697),
    .A2(net18167),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25265_ (.A1(net17789),
    .A2(net18190),
    .A3(_01270_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25266_ (.A1(_00994_),
    .A2(_00974_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25267_ (.A1(_01272_),
    .A2(net18680),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25268_ (.A1(_01112_),
    .A2(net18680),
    .A3(net18178),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25269_ (.A1(_01273_),
    .A2(_01274_),
    .B(net17820),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25270_ (.A1(_01271_),
    .A2(_01275_),
    .A3(net20000),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25271_ (.A1(_01267_),
    .A2(_01276_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25272_ (.A1(_01018_),
    .A2(_01277_),
    .A3(_01260_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25273_ (.A1(_01278_),
    .A2(_01240_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25274_ (.A1(_01046_),
    .A2(_00994_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25275_ (.I(_01093_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25276_ (.A1(_01280_),
    .A2(net18677),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25277_ (.A1(_01279_),
    .A2(_01281_),
    .B(net20003),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25278_ (.A1(_00907_),
    .A2(net18686),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _25279_ (.A1(net17288),
    .A2(net19725),
    .B1(net18670),
    .B2(net18182),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25280_ (.A1(_01282_),
    .A2(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25281_ (.A1(_01285_),
    .A2(net17815),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25282_ (.A1(net17793),
    .A2(net18671),
    .B(net20000),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25283_ (.A1(_01287_),
    .A2(_01224_),
    .B(net17814),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25284_ (.A1(_01140_),
    .A2(net17827),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25285_ (.A1(_01253_),
    .A2(net19731),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25286_ (.A1(_01290_),
    .A2(net18670),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25287_ (.A1(net17287),
    .A2(net17801),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25288_ (.A1(_01289_),
    .A2(_01292_),
    .A3(net20000),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25289_ (.A1(_01288_),
    .A2(_01293_),
    .B(_01180_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25290_ (.A1(_01294_),
    .A2(_01286_),
    .B(_01018_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25291_ (.A1(_01291_),
    .A2(net492),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25292_ (.A1(_01296_),
    .A2(net17491),
    .B(net17816),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25293_ (.I(_01220_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25294_ (.A1(_01297_),
    .A2(_01298_),
    .B(net20001),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25295_ (.A1(_01023_),
    .A2(net18165),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25296_ (.A1(_01109_),
    .A2(net17802),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25297_ (.A1(net19203),
    .A2(_00910_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25298_ (.A1(_01302_),
    .A2(net18673),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25299_ (.A1(_01301_),
    .A2(_01303_),
    .A3(net17819),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25300_ (.A1(_01300_),
    .A2(_01304_),
    .A3(net19729),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25301_ (.A1(_01299_),
    .A2(_01305_),
    .A3(net19999),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25302_ (.A1(_01295_),
    .A2(_01306_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25303_ (.A1(net428),
    .A2(_00987_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25304_ (.A1(_01308_),
    .A2(net18189),
    .A3(_01251_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25305_ (.A1(_01309_),
    .A2(net20222),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25306_ (.A1(_01098_),
    .A2(_01040_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25307_ (.A1(_01166_),
    .A2(_01311_),
    .A3(net17820),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25308_ (.A1(_01310_),
    .A2(_01312_),
    .B(net19725),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _25309_ (.A1(_01103_),
    .A2(net18657),
    .B1(net18654),
    .B2(_01062_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25310_ (.A1(net18193),
    .A2(_01314_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25311_ (.A1(net18654),
    .A2(net18694),
    .A3(_01060_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25312_ (.A1(_01095_),
    .A2(_01316_),
    .B(_01180_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25313_ (.A1(_01315_),
    .A2(_01317_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25314_ (.A1(_01313_),
    .A2(_01318_),
    .B(net20630),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25315_ (.A1(_01025_),
    .A2(net18670),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25316_ (.A1(_01320_),
    .A2(net17800),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _25317_ (.A1(_01321_),
    .A2(net17820),
    .A3(_01211_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25318_ (.A1(_01019_),
    .A2(_01112_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25319_ (.A1(_01323_),
    .A2(net18674),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25320_ (.A1(_01252_),
    .A2(net18181),
    .B(net18189),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25321_ (.I(_01281_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25322_ (.A1(_01324_),
    .A2(net17486),
    .A3(_01326_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25323_ (.A1(_01322_),
    .A2(_01327_),
    .A3(net20222),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25324_ (.A1(_01264_),
    .A2(_01323_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25325_ (.A1(_01167_),
    .A2(net19733),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25326_ (.A1(_01330_),
    .A2(_01176_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25327_ (.A1(_01329_),
    .A2(net18192),
    .A3(_01331_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25328_ (.I(_00990_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25329_ (.A1(_01109_),
    .A2(_01333_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25330_ (.A1(_01334_),
    .A2(_01107_),
    .A3(net17819),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25331_ (.A1(_01332_),
    .A2(_01335_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25332_ (.A1(_01336_),
    .A2(net19999),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25333_ (.A1(_01328_),
    .A2(_01337_),
    .A3(net19730),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25334_ (.A1(_01319_),
    .A2(_01338_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25335_ (.A1(_01307_),
    .A2(_01339_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25336_ (.A1(_01269_),
    .A2(net18190),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25337_ (.A1(_01340_),
    .A2(net17796),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25338_ (.A1(_01106_),
    .A2(_01120_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25339_ (.A1(net18163),
    .A2(net18684),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25340_ (.A1(_01272_),
    .A2(net18680),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25341_ (.A1(_01343_),
    .A2(_01344_),
    .A3(net17824),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25342_ (.A1(_01341_),
    .A2(net20002),
    .A3(_01345_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25343_ (.I(_01186_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25344_ (.A1(_01347_),
    .A2(_01060_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25345_ (.A1(net17485),
    .A2(net18194),
    .A3(_01150_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25346_ (.A1(_00972_),
    .A2(net17819),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25347_ (.I(net17498),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25348_ (.A1(_01350_),
    .A2(_01351_),
    .B(net20002),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25349_ (.A1(_01349_),
    .A2(_01352_),
    .B(net20226),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25350_ (.A1(_01346_),
    .A2(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25351_ (.A1(net18674),
    .A2(_01031_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25352_ (.A1(_01355_),
    .A2(_00910_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25353_ (.A1(_01356_),
    .A2(net17489),
    .B(net20002),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25354_ (.A1(_01135_),
    .A2(net17799),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25355_ (.A1(_01358_),
    .A2(_01042_),
    .A3(net18188),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25356_ (.A1(_01357_),
    .A2(_01359_),
    .B(net19999),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25357_ (.A1(_01264_),
    .A2(net18666),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25358_ (.A1(_01361_),
    .A2(net17820),
    .A3(_01204_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25359_ (.A1(net18659),
    .A2(net17809),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25360_ (.A1(_01363_),
    .A2(net18680),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25361_ (.A1(_01026_),
    .A2(net18194),
    .A3(_01364_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25362_ (.A1(_01362_),
    .A2(_01365_),
    .A3(net20002),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25363_ (.A1(_01360_),
    .A2(_01366_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25364_ (.A1(_01367_),
    .A2(_01354_),
    .A3(net20424),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25365_ (.A1(_01041_),
    .A2(net18662),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25366_ (.A1(net18173),
    .A2(net18691),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25367_ (.A1(_00988_),
    .A2(net18690),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _25368_ (.A1(net19725),
    .A2(_01369_),
    .A3(_01370_),
    .A4(_01371_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _25369_ (.A1(_01342_),
    .A2(net18680),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25370_ (.A1(net17498),
    .A2(net19202),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25371_ (.A1(_01373_),
    .A2(_01374_),
    .A3(net20002),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25372_ (.A1(_01372_),
    .A2(_01375_),
    .A3(net17819),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25373_ (.A1(_00977_),
    .A2(_01107_),
    .A3(net20002),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25374_ (.I(_15911_[0]),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25375_ (.A1(_01378_),
    .A2(net18701),
    .B(net20000),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25376_ (.A1(net18178),
    .A2(net18680),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25377_ (.A1(_01379_),
    .A2(_01380_),
    .B(net17825),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25378_ (.A1(_01377_),
    .A2(_01381_),
    .B(net19999),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25379_ (.A1(_01376_),
    .A2(_01382_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25380_ (.A1(_01247_),
    .A2(net17820),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25381_ (.A1(net18660),
    .A2(net18696),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25382_ (.A1(_01384_),
    .A2(_01385_),
    .A3(_01121_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25383_ (.A1(net18170),
    .A2(net17802),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25384_ (.A1(net18164),
    .A2(net17820),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25385_ (.A1(_01387_),
    .A2(_01388_),
    .B(net19725),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25386_ (.A1(_01386_),
    .A2(_01389_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25387_ (.A1(_01189_),
    .A2(_01031_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25388_ (.A1(_00949_),
    .A2(_01391_),
    .A3(net18192),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25389_ (.A1(_01137_),
    .A2(net18699),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25390_ (.A1(_01393_),
    .A2(net17820),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25391_ (.A1(_01394_),
    .A2(net18169),
    .B(net20004),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25392_ (.A1(_01395_),
    .A2(_01392_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25393_ (.A1(_01396_),
    .A2(_01390_),
    .A3(net19999),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25394_ (.A1(_01383_),
    .A2(_01397_),
    .A3(net20630),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25395_ (.A1(_01368_),
    .A2(_01398_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25396_ (.A1(_01330_),
    .A2(_01333_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25397_ (.A1(_01140_),
    .A2(_01167_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25398_ (.A1(net18700),
    .A2(_01399_),
    .B(_01400_),
    .C(net17821),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25399_ (.A1(net19199),
    .A2(net18678),
    .B(net17818),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25400_ (.A1(_01373_),
    .A2(_01402_),
    .B(net20004),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25401_ (.A1(_01401_),
    .A2(_01403_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25402_ (.A1(_00974_),
    .A2(net17827),
    .B(net18688),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25403_ (.A1(_01230_),
    .A2(net18688),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _25404_ (.A1(_01405_),
    .A2(net17814),
    .A3(_01406_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25405_ (.A1(_00994_),
    .A2(net18684),
    .A3(_01137_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25406_ (.A1(_01355_),
    .A2(net17816),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25407_ (.A1(_01408_),
    .A2(_01409_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25408_ (.A1(_01407_),
    .A2(_01410_),
    .B(net20003),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25409_ (.A1(_01404_),
    .A2(_01411_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25410_ (.A1(_01412_),
    .A2(net20222),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25411_ (.A1(_01189_),
    .A2(net17820),
    .Z(_01414_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25412_ (.A1(_01414_),
    .A2(_01195_),
    .B(net19725),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25413_ (.A1(_01109_),
    .A2(net17819),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25414_ (.A1(_01416_),
    .A2(_01303_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25415_ (.A1(_01415_),
    .A2(_01417_),
    .B(net20222),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25416_ (.A1(net17500),
    .A2(net17802),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25417_ (.A1(_01081_),
    .A2(_01419_),
    .A3(net18188),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25418_ (.A1(_01040_),
    .A2(net18684),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25419_ (.A1(_01421_),
    .A2(net18666),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25420_ (.A1(_01320_),
    .A2(_01254_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25421_ (.A1(_01422_),
    .A2(_01423_),
    .A3(net17820),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25422_ (.A1(_01420_),
    .A2(_01424_),
    .A3(net19730),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25423_ (.A1(_01418_),
    .A2(_01425_),
    .B(net20630),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25424_ (.A1(_01413_),
    .A2(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25425_ (.I(net18681),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25426_ (.I(net17287),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25427_ (.A1(net18174),
    .A2(_01428_),
    .B(_01429_),
    .C(net18187),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25428_ (.A1(net17489),
    .A2(net17490),
    .B(net20001),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25429_ (.A1(_01430_),
    .A2(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25430_ (.A1(net18179),
    .A2(net18678),
    .B(_00940_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25431_ (.A1(net18681),
    .A2(net18689),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25432_ (.A1(_01433_),
    .A2(_01434_),
    .B(net19725),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25433_ (.A1(net17495),
    .A2(net18176),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25434_ (.I(_01283_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25435_ (.A1(_01437_),
    .A2(net17488),
    .A3(_01436_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25436_ (.A1(_01435_),
    .A2(_01438_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25437_ (.A1(_01432_),
    .A2(net20223),
    .A3(_01439_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25438_ (.A1(net18683),
    .A2(net18692),
    .A3(net17802),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25439_ (.A1(net17811),
    .A2(net18673),
    .B(net18188),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25440_ (.A1(_01441_),
    .A2(_01442_),
    .B(net19725),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25441_ (.A1(_00949_),
    .A2(_00954_),
    .A3(_01371_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25442_ (.A1(_01443_),
    .A2(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25443_ (.A1(net19741),
    .A2(net18678),
    .B(net17817),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25444_ (.A1(_01446_),
    .A2(_01105_),
    .B(net20005),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25445_ (.A1(net17495),
    .A2(net18664),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25446_ (.A1(_01421_),
    .A2(net18661),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25447_ (.A1(_01448_),
    .A2(_01449_),
    .A3(_00940_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25448_ (.A1(_01447_),
    .A2(_01450_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25449_ (.A1(_01445_),
    .A2(_01451_),
    .A3(net19999),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25450_ (.A1(_01440_),
    .A2(_01452_),
    .A3(net20630),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25451_ (.A1(_01453_),
    .A2(_01427_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25452_ (.A1(net17797),
    .A2(net17490),
    .B(_01126_),
    .C(net17820),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25453_ (.A1(net18684),
    .A2(_15917_[0]),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25454_ (.A1(_01449_),
    .A2(net18191),
    .A3(_01455_),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25455_ (.A1(_01454_),
    .A2(net19726),
    .A3(_01456_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25456_ (.A1(_01201_),
    .A2(net18188),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25457_ (.I(net17803),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25458_ (.A1(_01369_),
    .A2(_01459_),
    .B(net18188),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25459_ (.A1(_01458_),
    .A2(_01460_),
    .B(net20001),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25460_ (.A1(_01457_),
    .A2(_01461_),
    .A3(net20222),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25461_ (.A1(net18684),
    .A2(net19199),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25462_ (.A1(_01308_),
    .A2(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25463_ (.A1(_01464_),
    .A2(net18190),
    .B(net20000),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25464_ (.A1(_01268_),
    .A2(net17492),
    .B(net19200),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25465_ (.A1(_01466_),
    .A2(net17822),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25466_ (.A1(_01465_),
    .A2(_01467_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25467_ (.A1(net18166),
    .A2(net17819),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25468_ (.A1(_01469_),
    .A2(_01061_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25469_ (.A1(net17797),
    .A2(net18692),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25470_ (.A1(_01303_),
    .A2(net18188),
    .A3(_01471_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25471_ (.A1(_01470_),
    .A2(_01472_),
    .A3(net20002),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25472_ (.A1(_01468_),
    .A2(_01473_),
    .A3(net19999),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25473_ (.A1(_01462_),
    .A2(_01474_),
    .A3(net20630),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25474_ (.A1(net17788),
    .A2(net18657),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25475_ (.A1(net17810),
    .A2(net18694),
    .B(net18189),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25476_ (.A1(_01476_),
    .A2(_01477_),
    .B(net19725),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25477_ (.A1(_01024_),
    .A2(net18675),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25478_ (.A1(_01479_),
    .A2(_01125_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25479_ (.A1(_01176_),
    .A2(net17487),
    .B(net17820),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25480_ (.A1(_01480_),
    .A2(_01481_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25481_ (.A1(_01478_),
    .A2(_01482_),
    .B(net19998),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25482_ (.A1(_01393_),
    .A2(_01133_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25483_ (.A1(_01484_),
    .A2(net17818),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25484_ (.A1(net18664),
    .A2(net18678),
    .A3(net18661),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25485_ (.A1(_01485_),
    .A2(_01486_),
    .B(net20005),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25486_ (.A1(_01437_),
    .A2(_01243_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25487_ (.A1(net17819),
    .A2(_01488_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25488_ (.A1(_01489_),
    .A2(_01487_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25489_ (.A1(_01490_),
    .A2(_01483_),
    .B(net20630),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25490_ (.A1(net17826),
    .A2(net17795),
    .B(_01032_),
    .C(_01371_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25491_ (.A1(_01421_),
    .A2(net17800),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25492_ (.A1(_01493_),
    .A2(_01049_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25493_ (.I(_01257_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25494_ (.A1(_01494_),
    .A2(_01495_),
    .B(net18189),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25495_ (.A1(_01492_),
    .A2(_01496_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25496_ (.A1(_01497_),
    .A2(net20001),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25497_ (.A1(_01264_),
    .A2(net428),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25498_ (.A1(_15916_[0]),
    .A2(_15925_[0]),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25499_ (.A1(net18697),
    .A2(_01500_),
    .B(net17817),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25500_ (.A1(_01499_),
    .A2(_01501_),
    .B(net20005),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25501_ (.A1(net17794),
    .A2(net17805),
    .B(net18670),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25502_ (.A1(_01384_),
    .A2(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25503_ (.A1(_01502_),
    .A2(_01504_),
    .B(net20224),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25504_ (.A1(_01498_),
    .A2(_01505_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25505_ (.A1(_01506_),
    .A2(_01491_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25506_ (.A1(_01507_),
    .A2(_01475_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25507_ (.A1(net18656),
    .A2(net18692),
    .A3(net18663),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25508_ (.A1(_01340_),
    .A2(_01508_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25509_ (.A1(net18684),
    .A2(net19737),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25510_ (.A1(_01348_),
    .A2(net18162),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25511_ (.A1(_01511_),
    .A2(net17819),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25512_ (.A1(_01509_),
    .A2(net19729),
    .A3(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25513_ (.A1(net18691),
    .A2(_01330_),
    .B(_01437_),
    .C(net18188),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25514_ (.A1(_01098_),
    .A2(net18656),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25515_ (.A1(_01515_),
    .A2(_01479_),
    .A3(net17820),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25516_ (.A1(_01514_),
    .A2(net20002),
    .A3(_01516_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25517_ (.A1(_01513_),
    .A2(_01517_),
    .A3(net20222),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25518_ (.A1(_01140_),
    .A2(_01024_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25519_ (.A1(_01325_),
    .A2(_01257_),
    .A3(_01519_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25520_ (.A1(_01135_),
    .A2(net17819),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25521_ (.A1(_01521_),
    .A2(_01369_),
    .B(net20000),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25522_ (.A1(_01520_),
    .A2(_01522_),
    .B(net20222),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25523_ (.A1(_01265_),
    .A2(_01493_),
    .A3(net18189),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25524_ (.A1(_01289_),
    .A2(_01183_),
    .A3(net17819),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25525_ (.A1(_01524_),
    .A2(_01525_),
    .A3(net20001),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25526_ (.A1(_01523_),
    .A2(_01526_),
    .B(_01018_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25527_ (.A1(_01518_),
    .A2(_01527_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25528_ (.A1(net18697),
    .A2(net18394),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25529_ (.A1(_01499_),
    .A2(_01529_),
    .A3(net17818),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25530_ (.A1(_01080_),
    .A2(net18672),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _25531_ (.A1(net18191),
    .A2(_01531_),
    .A3(net451),
    .A4(net17808),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25532_ (.A1(_01530_),
    .A2(_01532_),
    .A3(net20004),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25533_ (.A1(_01256_),
    .A2(_01087_),
    .B(net18698),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25534_ (.A1(net18176),
    .A2(net18171),
    .A3(net18670),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25535_ (.A1(_01534_),
    .A2(net18185),
    .A3(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25536_ (.A1(_01510_),
    .A2(net19731),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25537_ (.A1(_01463_),
    .A2(_00940_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25538_ (.A1(_01537_),
    .A2(_01538_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25539_ (.A1(_01296_),
    .A2(_01539_),
    .B(net20000),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25540_ (.A1(_01536_),
    .A2(_01540_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25541_ (.A1(_01533_),
    .A2(_01180_),
    .A3(_01541_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25542_ (.A1(_01378_),
    .A2(net18678),
    .B(net17817),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25543_ (.A1(_01543_),
    .A2(net452),
    .B(net20000),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25544_ (.I(_01538_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25545_ (.A1(_01121_),
    .A2(_01371_),
    .A3(_01545_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25546_ (.A1(_01544_),
    .A2(_01546_),
    .B(_01180_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25547_ (.A1(_01280_),
    .A2(net18685),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25548_ (.A1(net18677),
    .A2(_15925_[0]),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _25549_ (.A1(net18185),
    .A2(_01233_),
    .A3(_01548_),
    .A4(_01549_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25550_ (.A1(_01140_),
    .A2(net18661),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25551_ (.A1(_01094_),
    .A2(net18171),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25552_ (.A1(_01551_),
    .A2(_01552_),
    .A3(net17816),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25553_ (.A1(_01550_),
    .A2(_01553_),
    .A3(net20003),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25554_ (.A1(_01547_),
    .A2(_01554_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25555_ (.A1(_01542_),
    .A2(net20425),
    .A3(_01555_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25556_ (.A1(_01556_),
    .A2(_01528_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _25557_ (.I(\sa30_sr[7] ),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25558_ (.A1(_01557_),
    .A2(net21313),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25559_ (.A1(_10391_),
    .A2(net21299),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25560_ (.A1(_01558_),
    .A2(_01559_),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25561_ (.A1(net21311),
    .A2(_01560_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25562_ (.A1(_10415_),
    .A2(_10416_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25563_ (.A1(_01562_),
    .A2(_13583_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25564_ (.A1(_10419_),
    .A2(_10420_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25565_ (.A1(_01564_),
    .A2(_13587_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25566_ (.A1(_01563_),
    .A2(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25567_ (.I(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25568_ (.A1(_01561_),
    .A2(_01567_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25569_ (.A1(net21100),
    .A2(_01560_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25570_ (.A1(_01569_),
    .A2(_01566_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _25571_ (.A1(net469),
    .A2(_01570_),
    .B(net21501),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25572_ (.I(\text_in_r[105] ),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25573_ (.A1(_01572_),
    .A2(net21501),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25574_ (.A1(net20934),
    .A2(_01571_),
    .B(net21209),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25575_ (.A1(_01568_),
    .A2(_01570_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25576_ (.A1(_01575_),
    .A2(_10378_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25577_ (.I(net21209),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25578_ (.I(_01573_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25579_ (.A1(_01577_),
    .A2(net20876),
    .A3(net19724),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25580_ (.A1(_01574_),
    .A2(_01579_),
    .ZN(_15935_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25581_ (.A1(net21481),
    .A2(net21432),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25582_ (.A1(_01580_),
    .A2(net21362),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25583_ (.A1(_10339_),
    .A2(_10357_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25584_ (.A1(net21481),
    .A2(net21432),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25585_ (.A1(_01582_),
    .A2(_01583_),
    .B(net20987),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25586_ (.A1(_01581_),
    .A2(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25587_ (.A1(_10391_),
    .A2(_01557_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25588_ (.A1(net21313),
    .A2(net21299),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25589_ (.A1(_01587_),
    .A2(_01586_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25590_ (.A1(_01585_),
    .A2(net20875),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25591_ (.A1(_01581_),
    .A2(_01584_),
    .A3(net20877),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25592_ (.A1(_01589_),
    .A2(_01590_),
    .B(net21501),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25593_ (.I(\text_in_r[104] ),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25594_ (.A1(_01592_),
    .A2(net21501),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25595_ (.A1(_01591_),
    .A2(net20933),
    .B(net21210),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25596_ (.A1(_01589_),
    .A2(_01590_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25597_ (.A1(_01595_),
    .A2(net21076),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25598_ (.I(net21210),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25599_ (.I(_01593_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25600_ (.A1(net20221),
    .A2(_01597_),
    .A3(net20874),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25601_ (.A1(_01599_),
    .A2(_01594_),
    .ZN(_15940_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25602_ (.A1(_10427_),
    .A2(net21054),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25603_ (.A1(_10424_),
    .A2(_10426_),
    .A3(net21475),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25604_ (.A1(_01600_),
    .A2(_01601_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25605_ (.A1(_01602_),
    .A2(net20920),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25606_ (.A1(_01600_),
    .A2(_01601_),
    .A3(net503),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25607_ (.A1(_01603_),
    .A2(_01604_),
    .B(net21502),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25608_ (.I(\text_in_r[106] ),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25609_ (.A1(_01606_),
    .A2(net21502),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25610_ (.I(net21235),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25611_ (.A1(_01605_),
    .A2(_01607_),
    .B(_01608_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25612_ (.A1(_01603_),
    .A2(_01604_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25613_ (.A1(_01610_),
    .A2(net21075),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25614_ (.I(_01607_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25615_ (.A1(_01611_),
    .A2(net21235),
    .A3(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25616_ (.A1(_01609_),
    .A2(_01613_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output321 (.I(net321),
    .Z(text_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _25618_ (.A1(_01571_),
    .A2(_01573_),
    .B(_01577_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25619_ (.A1(_01578_),
    .A2(net21209),
    .A3(_01576_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25620_ (.A1(_01616_),
    .A2(_01615_),
    .ZN(_15930_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25621_ (.A1(_01605_),
    .A2(_01607_),
    .B(net21235),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25622_ (.A1(_01611_),
    .A2(_01608_),
    .A3(_01612_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25623_ (.A1(_01617_),
    .A2(_01618_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output320 (.I(net320),
    .Z(text_out[39]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output319 (.I(net319),
    .Z(text_out[38]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25626_ (.A1(_01591_),
    .A2(_01593_),
    .B(_01597_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25627_ (.A1(_01596_),
    .A2(net21210),
    .A3(_01598_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25628_ (.A1(_01621_),
    .A2(_01622_),
    .ZN(_15929_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25629_ (.A1(net19720),
    .A2(net19192),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25630_ (.A1(_10466_),
    .A2(_13689_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25631_ (.A1(net21420),
    .A2(\sa00_sr[3] ),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25632_ (.A1(_01624_),
    .A2(_01625_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25633_ (.I(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25634_ (.A1(_10423_),
    .A2(net20970),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25635_ (.A1(net21309),
    .A2(net21298),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25636_ (.A1(_01628_),
    .A2(_01629_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25637_ (.A1(_01627_),
    .A2(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25638_ (.I(_01630_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25639_ (.A1(_01632_),
    .A2(_01626_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25640_ (.A1(_01631_),
    .A2(_01633_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25641_ (.A1(net21305),
    .A2(_13679_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25642_ (.A1(_01634_),
    .A2(_01635_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25643_ (.A1(_10459_),
    .A2(_13679_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25644_ (.A1(_01631_),
    .A2(_01633_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25645_ (.A1(_01637_),
    .A2(_01638_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25646_ (.A1(_01636_),
    .A2(_01639_),
    .A3(net21075),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25647_ (.A1(net21501),
    .A2(\text_in_r[107] ),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25648_ (.A1(_01640_),
    .A2(_01641_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25649_ (.A1(_01642_),
    .A2(net21234),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25650_ (.I(net21234),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25651_ (.A1(_01640_),
    .A2(_01644_),
    .A3(_01641_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25652_ (.A1(_01643_),
    .A2(_01645_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25653_ (.A1(_01623_),
    .A2(net18636),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25654_ (.A1(net20985),
    .A2(_13655_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25655_ (.I(_10542_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25656_ (.A1(\sa30_sr[3] ),
    .A2(net21298),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25657_ (.A1(_01649_),
    .A2(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _25658_ (.A1(\sa30_sr[3] ),
    .A2(net21298),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25659_ (.A1(_01652_),
    .A2(_10542_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25660_ (.A1(_01651_),
    .A2(_01653_),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25661_ (.A1(_01648_),
    .A2(_01654_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25662_ (.A1(_01648_),
    .A2(_01654_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25663_ (.A1(_01655_),
    .A2(_01656_),
    .A3(net21075),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25664_ (.A1(net21501),
    .A2(\text_in_r[108] ),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25665_ (.A1(_01657_),
    .A2(_01658_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25666_ (.A1(_01659_),
    .A2(net21233),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25667_ (.I(net21233),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25668_ (.A1(_01657_),
    .A2(_01661_),
    .A3(_01658_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25669_ (.A1(_01660_),
    .A2(_01662_),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output318 (.I(net318),
    .Z(text_out[37]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25671_ (.A1(_01647_),
    .A2(net19715),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output317 (.I(net317),
    .Z(text_out[36]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25673_ (.A1(net19192),
    .A2(_15936_[0]),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25674_ (.A1(_01642_),
    .A2(_01644_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25675_ (.A1(_01640_),
    .A2(net21234),
    .A3(_01641_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25676_ (.A1(_01668_),
    .A2(_01669_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output316 (.I(net316),
    .Z(text_out[35]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25678_ (.A1(_01667_),
    .A2(net18623),
    .Z(_01672_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25679_ (.I(_15938_[0]),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25680_ (.A1(_01673_),
    .A2(net19189),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25681_ (.A1(_01672_),
    .A2(net17483),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25682_ (.A1(\sa30_sr[5] ),
    .A2(_13651_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25683_ (.A1(_01676_),
    .A2(_10581_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25684_ (.A1(_01676_),
    .A2(_10581_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25685_ (.A1(_01677_),
    .A2(_01678_),
    .A3(net21065),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25686_ (.A1(net21491),
    .A2(\text_in_r[109] ),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25687_ (.A1(_01679_),
    .A2(_01680_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25688_ (.A1(_01681_),
    .A2(net21232),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25689_ (.A1(_01681_),
    .A2(net21232),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25690_ (.A1(_01682_),
    .A2(_01683_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output315 (.I(net315),
    .Z(text_out[34]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output314 (.I(net314),
    .Z(text_out[33]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25693_ (.A1(_01665_),
    .A2(_01675_),
    .B(net19711),
    .ZN(_01687_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output313 (.I(net313),
    .Z(text_out[32]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25695_ (.A1(_01667_),
    .A2(net18636),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25696_ (.I(_01689_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25697_ (.A1(net19720),
    .A2(net19189),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25698_ (.A1(_01690_),
    .A2(net18621),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25699_ (.A1(_01659_),
    .A2(_01661_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25700_ (.A1(_01657_),
    .A2(net21233),
    .A3(_01658_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25701_ (.A1(_01693_),
    .A2(_01694_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output312 (.I(net312),
    .Z(text_out[31]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output311 (.I(net311),
    .Z(text_out[30]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25704_ (.A1(net19189),
    .A2(net17991),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25705_ (.A1(net17983),
    .A2(net19192),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25706_ (.A1(_01698_),
    .A2(_01699_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output310 (.I(net310),
    .Z(text_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25708_ (.A1(_01700_),
    .A2(net18632),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25709_ (.A1(_01692_),
    .A2(net19706),
    .A3(_01702_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25710_ (.A1(\sa10_sr[6] ),
    .A2(\sa30_sr[6] ),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25711_ (.A1(_13742_),
    .A2(_01704_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25712_ (.A1(_01705_),
    .A2(net20955),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25713_ (.A1(_01705_),
    .A2(net20955),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25714_ (.A1(net21492),
    .A2(\text_in_r[110] ),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _25715_ (.A1(_01706_),
    .A2(net21492),
    .A3(_01707_),
    .B(_01708_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25716_ (.A1(_01709_),
    .A2(net21231),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25717_ (.A1(_01709_),
    .A2(net21231),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25718_ (.A1(_01710_),
    .A2(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output309 (.I(net309),
    .Z(text_out[29]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25720_ (.A1(_01687_),
    .A2(_01703_),
    .B(net20422),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25721_ (.A1(net18648),
    .A2(net19192),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25722_ (.I(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output308 (.I(net308),
    .Z(text_out[28]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25724_ (.A1(_01716_),
    .A2(net18637),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25725_ (.A1(net19189),
    .A2(net17989),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25726_ (.A1(_01719_),
    .A2(net18634),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25727_ (.A1(_01720_),
    .A2(net19702),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25728_ (.A1(_15945_[0]),
    .A2(net19189),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25729_ (.A1(net18646),
    .A2(net17778),
    .A3(net18626),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25730_ (.A1(_01718_),
    .A2(_01721_),
    .A3(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25731_ (.A1(net18650),
    .A2(net19189),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output307 (.I(net307),
    .Z(text_out[27]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25733_ (.A1(_01690_),
    .A2(net18158),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output306 (.I(net306),
    .Z(text_out[26]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25735_ (.I(_15947_[0]),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25736_ (.A1(_01729_),
    .A2(net19190),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25737_ (.A1(net18647),
    .A2(net18632),
    .A3(net466),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output305 (.I(net305),
    .Z(text_out[25]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25739_ (.A1(_01727_),
    .A2(_01731_),
    .A3(net19706),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output304 (.I(net304),
    .Z(text_out[24]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25741_ (.A1(_01724_),
    .A2(_01733_),
    .A3(net19711),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _25742_ (.A1(net21298),
    .A2(net20915),
    .A3(net21050),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25743_ (.A1(net21500),
    .A2(\text_in_r[111] ),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25744_ (.A1(_01736_),
    .A2(net21065),
    .B(_01737_),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _25745_ (.A1(\u0.w[0][15] ),
    .A2(_01738_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _25746_ (.I(_01739_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output303 (.I(net303),
    .Z(text_out[23]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25748_ (.A1(_01714_),
    .A2(_01735_),
    .B(_01740_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25749_ (.I(_15932_[0]),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25750_ (.A1(net19189),
    .A2(_01743_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _25751_ (.I(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25752_ (.A1(_01745_),
    .A2(net18636),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25753_ (.I(_01746_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output302 (.I(net302),
    .Z(text_out[22]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output301 (.I(net301),
    .Z(text_out[21]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25756_ (.A1(net19192),
    .A2(_01743_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25757_ (.A1(net18634),
    .A2(_01750_),
    .B(_01663_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25758_ (.A1(_01718_),
    .A2(_01747_),
    .A3(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25759_ (.I(_15941_[0]),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25760_ (.A1(net19192),
    .A2(_01753_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25761_ (.I(_01754_),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25762_ (.I(_15931_[0]),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25763_ (.A1(net19189),
    .A2(_01756_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25764_ (.I(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output300 (.I(net300),
    .Z(text_out[20]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25766_ (.A1(_01755_),
    .A2(_01758_),
    .B(net18638),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25767_ (.A1(net18623),
    .A2(_01744_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _25768_ (.I(_01761_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25769_ (.A1(net19192),
    .A2(net17992),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25770_ (.A1(_01762_),
    .A2(_01763_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output299 (.I(net299),
    .Z(text_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25772_ (.A1(_01764_),
    .A2(_01760_),
    .B(net19703),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25773_ (.A1(_01752_),
    .A2(_01766_),
    .B(net19711),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25774_ (.A1(net19723),
    .A2(net19189),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25775_ (.A1(_01768_),
    .A2(net18636),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25776_ (.A1(net18650),
    .A2(net19720),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25777_ (.A1(_01769_),
    .A2(net18156),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25778_ (.A1(net18653),
    .A2(net19720),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output298 (.I(net298),
    .Z(text_out[19]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25780_ (.A1(net19723),
    .A2(net19192),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25781_ (.A1(_01772_),
    .A2(net18623),
    .A3(_01774_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25782_ (.A1(_01771_),
    .A2(_01775_),
    .A3(net19704),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _25783_ (.I(_01684_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output297 (.I(net297),
    .Z(text_out[18]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25785_ (.A1(_01744_),
    .A2(net18640),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25786_ (.A1(net19192),
    .A2(_15945_[0]),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25787_ (.A1(_01779_),
    .A2(net17774),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output296 (.I(net296),
    .Z(text_out[17]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25789_ (.A1(net19189),
    .A2(net17985),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output295 (.I(net295),
    .Z(text_out[16]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25791_ (.A1(_01763_),
    .A2(_01783_),
    .A3(net18623),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25792_ (.A1(_01781_),
    .A2(net19712),
    .A3(_01785_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25793_ (.A1(_01776_),
    .A2(net19183),
    .A3(_01786_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25794_ (.A1(_01767_),
    .A2(net20422),
    .A3(_01787_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25795_ (.A1(_01742_),
    .A2(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25796_ (.A1(net19192),
    .A2(net17991),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25797_ (.A1(_01790_),
    .A2(net18636),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output294 (.I(net294),
    .Z(text_out[15]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25799_ (.A1(net18636),
    .A2(_15954_[0]),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25800_ (.A1(_01791_),
    .A2(_01793_),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output293 (.I(net293),
    .Z(text_out[14]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25802_ (.A1(_01794_),
    .A2(net19710),
    .B(_01777_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25803_ (.I(_15936_[0]),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25804_ (.A1(net19189),
    .A2(_01797_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25805_ (.A1(net19192),
    .A2(net17986),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25806_ (.A1(_01798_),
    .A2(_01799_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output292 (.I(net292),
    .Z(text_out[13]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _25808_ (.A1(_01800_),
    .A2(net18643),
    .B(net19702),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25809_ (.A1(_01774_),
    .A2(_01757_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25810_ (.A1(_01803_),
    .A2(net18633),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25811_ (.A1(net19192),
    .A2(net17990),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25812_ (.I(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output291 (.I(net291),
    .Z(text_out[12]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25814_ (.A1(_01806_),
    .A2(net18642),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25815_ (.A1(_01802_),
    .A2(_01804_),
    .A3(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25816_ (.A1(_01796_),
    .A2(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25817_ (.A1(_01755_),
    .A2(net18638),
    .B(net19715),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25818_ (.I(_01719_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25819_ (.A1(_01812_),
    .A2(net18634),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25820_ (.I(_01798_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25821_ (.A1(_01814_),
    .A2(net18638),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25822_ (.A1(_01811_),
    .A2(net17281),
    .A3(_01815_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25823_ (.I(_15943_[0]),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25824_ (.A1(net19192),
    .A2(_01817_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25825_ (.A1(_01818_),
    .A2(net18623),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25826_ (.A1(net19189),
    .A2(net17988),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25827_ (.A1(_01819_),
    .A2(net470),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25828_ (.A1(_01821_),
    .A2(_01721_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25829_ (.A1(_01816_),
    .A2(_01822_),
    .A3(net19186),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25830_ (.A1(_01810_),
    .A2(_01823_),
    .A3(net20422),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25831_ (.A1(net19192),
    .A2(_01756_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25832_ (.A1(_01825_),
    .A2(net18636),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25833_ (.A1(_01674_),
    .A2(net18623),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25834_ (.A1(_01826_),
    .A2(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25835_ (.A1(net17480),
    .A2(net19715),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25836_ (.A1(_01828_),
    .A2(_01829_),
    .B(net19711),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25837_ (.A1(net19192),
    .A2(_15941_[0]),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25838_ (.A1(net19722),
    .A2(net19193),
    .B(net17766),
    .C(net18627),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25839_ (.A1(net19189),
    .A2(net18652),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25840_ (.A1(_01833_),
    .A2(net18642),
    .A3(net17772),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25841_ (.A1(_01832_),
    .A2(net19712),
    .A3(_01834_),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25842_ (.A1(_01830_),
    .A2(_01835_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25843_ (.A1(net19189),
    .A2(net17984),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25844_ (.I(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25845_ (.A1(_01838_),
    .A2(net18636),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25846_ (.A1(_01839_),
    .A2(_01761_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25847_ (.I(_01799_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25848_ (.A1(_01841_),
    .A2(net18636),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25849_ (.A1(_01842_),
    .A2(net19702),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25850_ (.A1(_01840_),
    .A2(_01843_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output290 (.I(net290),
    .Z(text_out[127]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25852_ (.A1(_01723_),
    .A2(net19712),
    .A3(net17276),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25853_ (.A1(_01844_),
    .A2(_01846_),
    .A3(net19711),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _25854_ (.I(_01712_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output289 (.I(net289),
    .Z(text_out[126]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25856_ (.A1(_01836_),
    .A2(_01847_),
    .A3(_01848_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25857_ (.A1(_01824_),
    .A2(_01850_),
    .A3(net20218),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25858_ (.A1(_01789_),
    .A2(_01851_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _25859_ (.A1(net18641),
    .A2(_15961_[0]),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25860_ (.A1(_01725_),
    .A2(net18623),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25861_ (.A1(_01843_),
    .A2(_01852_),
    .A3(_01853_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25862_ (.A1(_01730_),
    .A2(_01750_),
    .A3(net18631),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25863_ (.A1(_01802_),
    .A2(_01855_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25864_ (.A1(_01854_),
    .A2(_01856_),
    .A3(net19711),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25865_ (.A1(net18647),
    .A2(_01762_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25866_ (.A1(_01674_),
    .A2(net18636),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25867_ (.I(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25868_ (.A1(_01860_),
    .A2(net18617),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25869_ (.A1(_01861_),
    .A2(_01858_),
    .A3(net19706),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25870_ (.A1(_01833_),
    .A2(_01770_),
    .A3(net18642),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25871_ (.A1(net19194),
    .A2(net17770),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25872_ (.I(_01864_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output288 (.I(net288),
    .Z(text_out[125]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25874_ (.A1(_01865_),
    .A2(net18632),
    .B(net19706),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25875_ (.A1(_01863_),
    .A2(_01867_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25876_ (.A1(_01868_),
    .A2(_01862_),
    .A3(net19186),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25877_ (.A1(_01869_),
    .A2(_01857_),
    .A3(net20422),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25878_ (.A1(_01780_),
    .A2(net18623),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25879_ (.A1(_01871_),
    .A2(net17784),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25880_ (.A1(net19189),
    .A2(net17986),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25881_ (.I(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25882_ (.A1(_01874_),
    .A2(net18643),
    .B(net19708),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25883_ (.A1(_01872_),
    .A2(_01875_),
    .B(net19711),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25884_ (.A1(_01729_),
    .A2(net19192),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25885_ (.A1(_01877_),
    .A2(net18623),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25886_ (.A1(_01878_),
    .A2(_01725_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _25887_ (.I(_15945_[0]),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25888_ (.A1(net19191),
    .A2(_01880_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25889_ (.A1(_01881_),
    .A2(net18643),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25890_ (.A1(_01879_),
    .A2(net19706),
    .A3(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25891_ (.A1(_01876_),
    .A2(_01883_),
    .B(net20422),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25892_ (.A1(net389),
    .A2(net19723),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25893_ (.A1(_01885_),
    .A2(_01691_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25894_ (.A1(_01886_),
    .A2(net18633),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25895_ (.A1(net17470),
    .A2(net18620),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25896_ (.A1(_01887_),
    .A2(_01888_),
    .A3(net19712),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25897_ (.A1(net17466),
    .A2(net17284),
    .B(net18633),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25898_ (.A1(_01803_),
    .A2(net18643),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25899_ (.A1(_01890_),
    .A2(_01891_),
    .A3(net19707),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output287 (.I(net287),
    .Z(text_out[124]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25901_ (.A1(_01889_),
    .A2(_01892_),
    .A3(net19711),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25902_ (.A1(_01884_),
    .A2(_01894_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25903_ (.A1(_01895_),
    .A2(net20219),
    .A3(_01870_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _25904_ (.A1(_01716_),
    .A2(_01827_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25905_ (.A1(net389),
    .A2(net19192),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25906_ (.A1(_01769_),
    .A2(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25907_ (.A1(_01897_),
    .A2(_01899_),
    .A3(net19711),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25908_ (.A1(_01691_),
    .A2(net18636),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25909_ (.A1(_01901_),
    .A2(_01763_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25910_ (.A1(_01672_),
    .A2(net17779),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25911_ (.A1(_01902_),
    .A2(_01903_),
    .A3(_01777_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25912_ (.A1(_01900_),
    .A2(_01904_),
    .A3(net19703),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25913_ (.A1(_01684_),
    .A2(net18634),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25914_ (.A1(_01722_),
    .A2(net18636),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25915_ (.I(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25916_ (.A1(_01908_),
    .A2(_01831_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25917_ (.A1(_15957_[0]),
    .A2(net18152),
    .B(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output286 (.I(net286),
    .Z(text_out[123]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25919_ (.A1(_01910_),
    .A2(net19715),
    .B(_01848_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25920_ (.A1(_01905_),
    .A2(_01912_),
    .B(_01740_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25921_ (.A1(net18635),
    .A2(_01758_),
    .B(net17480),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25922_ (.I(net18617),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25923_ (.A1(_01915_),
    .A2(net18638),
    .B(net19715),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _25924_ (.A1(net18636),
    .A2(_01790_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _25925_ (.I(_01917_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25926_ (.A1(_01914_),
    .A2(_01916_),
    .A3(_01918_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25927_ (.A1(_01769_),
    .A2(_01763_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25928_ (.A1(_01897_),
    .A2(_01920_),
    .A3(net19716),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25929_ (.A1(_01919_),
    .A2(_01921_),
    .A3(net19185),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _25930_ (.I(_01647_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25931_ (.A1(_01923_),
    .A2(net17779),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25932_ (.A1(_01924_),
    .A2(net19715),
    .A3(net17282),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _25933_ (.I(_15933_[0]),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25934_ (.A1(net19192),
    .A2(_01926_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25935_ (.A1(_01927_),
    .A2(net18636),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _25936_ (.I(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25937_ (.A1(_01929_),
    .A2(net17479),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25938_ (.A1(_01872_),
    .A2(_01930_),
    .A3(net19703),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25939_ (.A1(net19711),
    .A2(_01931_),
    .A3(_01925_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25940_ (.A1(_01932_),
    .A2(_01922_),
    .A3(_01848_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25941_ (.A1(_01933_),
    .A2(_01913_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25942_ (.A1(_01934_),
    .A2(_01896_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25943_ (.A1(_01689_),
    .A2(net19712),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25944_ (.A1(_01871_),
    .A2(net17478),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25945_ (.A1(_01935_),
    .A2(_01936_),
    .B(_01848_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25946_ (.A1(_01898_),
    .A2(net18640),
    .A3(net17476),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25947_ (.A1(_01768_),
    .A2(net17768),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25948_ (.A1(_01939_),
    .A2(net18626),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25949_ (.A1(_01938_),
    .A2(_01940_),
    .A3(net19710),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25950_ (.A1(_01937_),
    .A2(_01941_),
    .B(net19711),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25951_ (.A1(_01818_),
    .A2(net18636),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25952_ (.A1(_01943_),
    .A2(_01691_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25953_ (.A1(_01762_),
    .A2(net17772),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output285 (.I(net285),
    .Z(text_out[122]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25955_ (.A1(_01945_),
    .A2(_01944_),
    .B(net19705),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _25956_ (.A1(net18161),
    .A2(net18625),
    .A3(net17765),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25957_ (.A1(_01768_),
    .A2(_01699_),
    .A3(net18642),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25958_ (.A1(_01949_),
    .A2(net19702),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25959_ (.A1(_01948_),
    .A2(_01950_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25960_ (.A1(_01947_),
    .A2(_01951_),
    .B(_01848_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25961_ (.A1(_01952_),
    .A2(_01942_),
    .B(_01740_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _25962_ (.A1(_01798_),
    .A2(net18623),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _25963_ (.A1(net17769),
    .A2(_01954_),
    .B(net19708),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25964_ (.A1(_01955_),
    .A2(_01834_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25965_ (.A1(_01956_),
    .A2(net20422),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25966_ (.A1(_01672_),
    .A2(_01833_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25967_ (.A1(_01873_),
    .A2(_01699_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25968_ (.A1(_01959_),
    .A2(net18642),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25969_ (.A1(_01958_),
    .A2(_01960_),
    .B(net19712),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25970_ (.A1(_01957_),
    .A2(_01961_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _25971_ (.A1(net19192),
    .A2(net17786),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25972_ (.A1(net18620),
    .A2(net18633),
    .A3(net17460),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25973_ (.A1(_01699_),
    .A2(net18633),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25974_ (.A1(_01964_),
    .A2(net19707),
    .A3(_01965_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25975_ (.A1(net18154),
    .A2(net18642),
    .B(net19712),
    .C(_01799_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25976_ (.A1(_01848_),
    .A2(net17277),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25977_ (.A1(_01966_),
    .A2(_01967_),
    .B(_01968_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25978_ (.A1(_01969_),
    .A2(_01962_),
    .B(net19711),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25979_ (.A1(_01970_),
    .A2(_01953_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _25980_ (.A1(net18648),
    .A2(net19195),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _25981_ (.A1(_01972_),
    .A2(net18634),
    .A3(_01825_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25982_ (.A1(net19189),
    .A2(net17777),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _25983_ (.A1(net19718),
    .A2(net17771),
    .A3(net17459),
    .A4(net19188),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25984_ (.A1(_01973_),
    .A2(_01975_),
    .B(net19713),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _25985_ (.A1(net18155),
    .A2(net18156),
    .A3(net18627),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _25986_ (.A1(net18634),
    .A2(_15957_[0]),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25987_ (.A1(_01977_),
    .A2(net19713),
    .A3(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25988_ (.A1(_01979_),
    .A2(net19711),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25989_ (.A1(net18161),
    .A2(net18625),
    .A3(_01691_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _25990_ (.A1(_01981_),
    .A2(_01834_),
    .A3(net19710),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _25991_ (.A1(_01820_),
    .A2(net18623),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25992_ (.A1(_01983_),
    .A2(net17474),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25993_ (.A1(net17982),
    .A2(net18641),
    .B(net19710),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25994_ (.A1(_01984_),
    .A2(_01985_),
    .B(net19711),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25995_ (.A1(_01982_),
    .A2(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _25996_ (.A1(_01976_),
    .A2(_01980_),
    .B(_01987_),
    .C(_01848_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _25997_ (.A1(_01762_),
    .A2(net17461),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25998_ (.A1(_01758_),
    .A2(net18638),
    .B(net19703),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _25999_ (.A1(_01989_),
    .A2(_01990_),
    .B(net19711),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26000_ (.A1(_01673_),
    .A2(_01926_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26001_ (.A1(_01992_),
    .A2(net19191),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26002_ (.A1(_01871_),
    .A2(net17271),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26003_ (.A1(_01994_),
    .A2(net17209),
    .A3(net19703),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26004_ (.A1(_01995_),
    .A2(_01991_),
    .B(_01848_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26005_ (.A1(_15952_[0]),
    .A2(net18636),
    .B(_01689_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26006_ (.A1(_01997_),
    .A2(net19710),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26007_ (.A1(net18641),
    .A2(_15963_[0]),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26008_ (.A1(_01958_),
    .A2(net19710),
    .A3(_01999_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26009_ (.A1(_01998_),
    .A2(net19711),
    .A3(_02000_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26010_ (.A1(_01996_),
    .A2(_02001_),
    .B(net20421),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26011_ (.A1(_01988_),
    .A2(_02002_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26012_ (.A1(_01971_),
    .A2(_02003_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26013_ (.A1(net17473),
    .A2(net17477),
    .A3(net18636),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26014_ (.A1(_01775_),
    .A2(net19703),
    .A3(_02004_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26015_ (.A1(_01783_),
    .A2(net17787),
    .A3(net18624),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26016_ (.A1(net468),
    .A2(_01750_),
    .A3(net18639),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26017_ (.A1(_02006_),
    .A2(_02007_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26018_ (.A1(_02008_),
    .A2(net19712),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26019_ (.A1(_02005_),
    .A2(_02009_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26020_ (.A1(_02010_),
    .A2(_01848_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26021_ (.A1(net18161),
    .A2(net18644),
    .A3(net17783),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26022_ (.A1(net17478),
    .A2(net464),
    .A3(net18623),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26023_ (.A1(_02012_),
    .A2(net19712),
    .A3(_02013_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26024_ (.A1(net18616),
    .A2(net18636),
    .A3(_01974_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26025_ (.A1(net17471),
    .A2(net680),
    .A3(net18623),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26026_ (.A1(_02015_),
    .A2(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26027_ (.A1(_02017_),
    .A2(net19703),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26028_ (.A1(_02014_),
    .A2(_02018_),
    .A3(net20422),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26029_ (.A1(_02011_),
    .A2(_02019_),
    .A3(net19182),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26030_ (.A1(net18161),
    .A2(net18645),
    .A3(net18622),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26031_ (.A1(_02021_),
    .A2(_01751_),
    .B(_01848_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26032_ (.A1(_01772_),
    .A2(net18640),
    .A3(_01768_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26033_ (.A1(net18161),
    .A2(net18625),
    .A3(net17476),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26034_ (.A1(_02023_),
    .A2(_02024_),
    .A3(net19712),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26035_ (.A1(_02022_),
    .A2(_02025_),
    .B(net19182),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26036_ (.A1(_01943_),
    .A2(net17784),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26037_ (.A1(_01879_),
    .A2(_02027_),
    .A3(net19706),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26038_ (.I(_01672_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26039_ (.A1(_02023_),
    .A2(net19712),
    .A3(_02029_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26040_ (.A1(_02028_),
    .A2(_02030_),
    .A3(_01848_),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26041_ (.A1(_02026_),
    .A2(_02031_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26042_ (.A1(_02020_),
    .A2(_02032_),
    .A3(net20220),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26043_ (.A1(_01906_),
    .A2(_01750_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26044_ (.A1(_01813_),
    .A2(net19702),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26045_ (.A1(_02034_),
    .A2(_02035_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26046_ (.A1(_01831_),
    .A2(net18636),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _26047_ (.A1(_01972_),
    .A2(_01777_),
    .A3(_02037_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26048_ (.A1(_01746_),
    .A2(_01777_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26049_ (.A1(_02039_),
    .A2(_02038_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26050_ (.A1(_02036_),
    .A2(_02040_),
    .B(_01848_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26051_ (.A1(_01878_),
    .A2(net17271),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26052_ (.A1(net18647),
    .A2(net17476),
    .A3(net18636),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26053_ (.A1(_02043_),
    .A2(_02042_),
    .A3(net19711),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26054_ (.A1(_01838_),
    .A2(net18629),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26055_ (.A1(_01944_),
    .A2(_01777_),
    .A3(_02045_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26056_ (.A1(_02044_),
    .A2(_02046_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26057_ (.A1(_02047_),
    .A2(net19714),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26058_ (.A1(_02041_),
    .A2(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26059_ (.A1(_01863_),
    .A2(_01804_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26060_ (.A1(_02050_),
    .A2(net19712),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26061_ (.A1(_01700_),
    .A2(net18636),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26062_ (.A1(_01623_),
    .A2(_01837_),
    .B(net18636),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26063_ (.A1(_02052_),
    .A2(_02053_),
    .B(net19706),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26064_ (.A1(_02051_),
    .A2(net19184),
    .A3(_02054_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26065_ (.A1(net17468),
    .A2(_01993_),
    .A3(net18623),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26066_ (.A1(_01909_),
    .A2(_02056_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26067_ (.A1(_02057_),
    .A2(net19712),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26068_ (.A1(_01949_),
    .A2(net19706),
    .B(_01777_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26069_ (.A1(_02058_),
    .A2(_02059_),
    .B(net20422),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26070_ (.A1(_02055_),
    .A2(_02060_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26071_ (.A1(_02049_),
    .A2(_02061_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26072_ (.A1(net20421),
    .A2(_02062_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26073_ (.A1(_02033_),
    .A2(_02063_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26074_ (.A1(_01918_),
    .A2(net17765),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26075_ (.A1(_02064_),
    .A2(_01843_),
    .B(net19711),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26076_ (.A1(_01730_),
    .A2(net18636),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26077_ (.A1(net17270),
    .A2(net17475),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26078_ (.A1(_02067_),
    .A2(_01821_),
    .A3(net19717),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26079_ (.A1(_02065_),
    .A2(_02068_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26080_ (.A1(_01983_),
    .A2(net18161),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26081_ (.A1(_02070_),
    .A2(net19709),
    .A3(_01960_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26082_ (.A1(_01898_),
    .A2(net17472),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26083_ (.A1(_02072_),
    .A2(net18633),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26084_ (.A1(net17211),
    .A2(_02073_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26085_ (.A1(_02071_),
    .A2(_02074_),
    .A3(net19711),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26086_ (.A1(_02069_),
    .A2(_02075_),
    .A3(net20422),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26087_ (.A1(net18161),
    .A2(net18619),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26088_ (.A1(_02077_),
    .A2(net18627),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26089_ (.A1(_02078_),
    .A2(_01902_),
    .A3(net19716),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26090_ (.I(net17280),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26091_ (.A1(net19703),
    .A2(net17780),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26092_ (.A1(_02080_),
    .A2(_02081_),
    .B(net19711),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26093_ (.A1(_02079_),
    .A2(_02082_),
    .B(net20422),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26094_ (.A1(_01899_),
    .A2(_01977_),
    .A3(net19716),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26095_ (.A1(_01725_),
    .A2(net18153),
    .A3(net18645),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26096_ (.A1(net18159),
    .A2(net18627),
    .A3(net17776),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26097_ (.A1(_02085_),
    .A2(_02086_),
    .A3(net19703),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26098_ (.A1(_02084_),
    .A2(_02087_),
    .A3(net19711),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26099_ (.A1(_02083_),
    .A2(_02088_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26100_ (.A1(_02076_),
    .A2(_02089_),
    .A3(net20219),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26101_ (.A1(net17771),
    .A2(net18623),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26102_ (.A1(net18639),
    .A2(net17764),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _26103_ (.A1(_02091_),
    .A2(net19712),
    .A3(_02092_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26104_ (.A1(_02093_),
    .A2(_01848_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26105_ (.A1(_01815_),
    .A2(net19703),
    .Z(_02095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26106_ (.A1(_01819_),
    .A2(_01725_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26107_ (.A1(_02095_),
    .A2(_02096_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26108_ (.A1(_02094_),
    .A2(_02097_),
    .B(net19711),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26109_ (.A1(_01723_),
    .A2(net19712),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26110_ (.A1(net17210),
    .A2(net17772),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26111_ (.A1(_02099_),
    .A2(_02100_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26112_ (.A1(_01871_),
    .A2(_01929_),
    .A3(net19717),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26113_ (.A1(_02101_),
    .A2(_02102_),
    .A3(_01848_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26114_ (.A1(_02098_),
    .A2(_02103_),
    .B(_01740_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26115_ (.A1(net18157),
    .A2(net17464),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26116_ (.A1(net18628),
    .A2(net19193),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26117_ (.A1(_02106_),
    .A2(net19704),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26118_ (.A1(_02105_),
    .A2(_02107_),
    .B(net20422),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26119_ (.A1(_01758_),
    .A2(net18638),
    .B(net19715),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26120_ (.A1(_01897_),
    .A2(_02109_),
    .A3(net17481),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26121_ (.A1(_02108_),
    .A2(_02110_),
    .B(net19183),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26122_ (.A1(_01772_),
    .A2(net18161),
    .A3(net18639),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26123_ (.A1(net17279),
    .A2(net18619),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26124_ (.A1(_02112_),
    .A2(_02113_),
    .A3(net19704),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26125_ (.A1(net17775),
    .A2(net17285),
    .A3(net17278),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26126_ (.A1(_02114_),
    .A2(_02115_),
    .A3(net20422),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26127_ (.A1(_02111_),
    .A2(_02116_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26128_ (.A1(_02104_),
    .A2(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26129_ (.A1(_02090_),
    .A2(_02118_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26130_ (.A1(_01943_),
    .A2(net17767),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26131_ (.I(_01992_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26132_ (.A1(_01963_),
    .A2(net18625),
    .A3(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26133_ (.A1(_02121_),
    .A2(net19710),
    .A3(_02119_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26134_ (.A1(_01959_),
    .A2(net18633),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26135_ (.A1(_01718_),
    .A2(_01721_),
    .A3(_02123_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26136_ (.A1(_02124_),
    .A2(_02122_),
    .B(net19182),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26137_ (.A1(_02053_),
    .A2(_01779_),
    .B(net19712),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26138_ (.A1(net17275),
    .A2(net17465),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26139_ (.A1(_02127_),
    .A2(net19710),
    .B(_01777_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26140_ (.A1(_02128_),
    .A2(_02126_),
    .B(net20422),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26141_ (.A1(_02129_),
    .A2(_02125_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26142_ (.A1(net18648),
    .A2(net18627),
    .B(net19704),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26143_ (.A1(_02112_),
    .A2(_02131_),
    .B(net19711),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26144_ (.A1(_01923_),
    .A2(_01885_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26145_ (.A1(_01722_),
    .A2(_01831_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26146_ (.A1(_02134_),
    .A2(net18627),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26147_ (.A1(_02133_),
    .A2(net19704),
    .A3(_02135_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26148_ (.A1(_02132_),
    .A2(_02136_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _26149_ (.A1(_01825_),
    .A2(_01761_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26150_ (.A1(net17782),
    .A2(net18636),
    .B(net19705),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26151_ (.A1(_02138_),
    .A2(_02139_),
    .B(_01777_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26152_ (.A1(_01972_),
    .A2(net17272),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26153_ (.A1(_02141_),
    .A2(net17462),
    .B(net19703),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26154_ (.A1(_02140_),
    .A2(_02142_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26155_ (.A1(_02143_),
    .A2(net20422),
    .A3(_02137_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26156_ (.A1(_02144_),
    .A2(_02130_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26157_ (.A1(_01740_),
    .A2(_02145_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26158_ (.A1(_01901_),
    .A2(net17461),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26159_ (.A1(_02099_),
    .A2(_02147_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26160_ (.A1(net17273),
    .A2(net17464),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26161_ (.A1(net17283),
    .A2(net18635),
    .B(net19715),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26162_ (.A1(_02149_),
    .A2(_02150_),
    .B(net19185),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26163_ (.A1(_02148_),
    .A2(_02151_),
    .B(net20422),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26164_ (.A1(net18627),
    .A2(net19722),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26165_ (.A1(_01771_),
    .A2(net19714),
    .A3(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26166_ (.A1(_01943_),
    .A2(_01725_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26167_ (.A1(_01762_),
    .A2(net17787),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26168_ (.A1(_02155_),
    .A2(_02156_),
    .A3(net19704),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26169_ (.A1(_02154_),
    .A2(_02157_),
    .A3(net19184),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26170_ (.A1(_02158_),
    .A2(_02152_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26171_ (.I(net17274),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26172_ (.A1(_01843_),
    .A2(_02160_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26173_ (.A1(net17286),
    .A2(net17779),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26174_ (.A1(net18630),
    .A2(net17271),
    .B(net19705),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26175_ (.A1(_02163_),
    .A2(_02162_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26176_ (.A1(_02161_),
    .A2(net19184),
    .A3(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26177_ (.A1(net18634),
    .A2(net17777),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26178_ (.A1(net17463),
    .A2(_02166_),
    .A3(net19712),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26179_ (.A1(_02167_),
    .A2(net19711),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26180_ (.I(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26181_ (.A1(_01762_),
    .A2(net17766),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26182_ (.A1(net17783),
    .A2(net17464),
    .A3(net18644),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26183_ (.A1(_02170_),
    .A2(net19704),
    .A3(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26184_ (.A1(_02169_),
    .A2(_02172_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26185_ (.A1(_02173_),
    .A2(_02165_),
    .A3(net20422),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26186_ (.A1(_02159_),
    .A2(net20421),
    .A3(_02174_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26187_ (.A1(_02146_),
    .A2(_02175_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26188_ (.A1(_01770_),
    .A2(net18632),
    .A3(net18617),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26189_ (.A1(net18158),
    .A2(net18643),
    .A3(_01864_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26190_ (.A1(_02176_),
    .A2(_02177_),
    .A3(net19715),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26191_ (.A1(_02066_),
    .A2(net18618),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26192_ (.A1(_02176_),
    .A2(_02179_),
    .B(net19715),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26193_ (.A1(_02178_),
    .A2(_02180_),
    .B(net19187),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26194_ (.A1(net17784),
    .A2(net18632),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26195_ (.A1(_02053_),
    .A2(net19706),
    .A3(_02182_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26196_ (.A1(_01692_),
    .A2(net19706),
    .A3(_01852_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26197_ (.A1(_02183_),
    .A2(net19711),
    .A3(_02184_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26198_ (.A1(_02181_),
    .A2(_02185_),
    .A3(_01848_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26199_ (.I(_15951_[0]),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26200_ (.A1(_02187_),
    .A2(net18627),
    .B(net19704),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26201_ (.A1(_02155_),
    .A2(_02188_),
    .B(net19711),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26202_ (.A1(net17274),
    .A2(net17784),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26203_ (.A1(_01916_),
    .A2(_02190_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26204_ (.A1(_02189_),
    .A2(_02191_),
    .B(_01848_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26205_ (.A1(_02096_),
    .A2(net17458),
    .B(net19716),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26206_ (.A1(_02193_),
    .A2(net17208),
    .B(net19711),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26207_ (.A1(_02192_),
    .A2(_02194_),
    .B(_01740_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26208_ (.A1(_02186_),
    .A2(_02195_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26209_ (.A1(_01772_),
    .A2(net18161),
    .A3(net18623),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26210_ (.A1(_15950_[0]),
    .A2(net17981),
    .B(net18639),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26211_ (.A1(_02197_),
    .A2(net19712),
    .A3(_02198_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26212_ (.A1(_01806_),
    .A2(net17467),
    .B(net18627),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26213_ (.A1(_02200_),
    .A2(_02109_),
    .B(net19711),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26214_ (.A1(_02199_),
    .A2(_02201_),
    .B(net20422),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26215_ (.A1(_02045_),
    .A2(net19705),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26216_ (.A1(net17469),
    .A2(net18619),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26217_ (.A1(_02106_),
    .A2(_02120_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26218_ (.A1(_02203_),
    .A2(_02204_),
    .A3(_02205_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26219_ (.A1(_01943_),
    .A2(net465),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26220_ (.A1(net19193),
    .A2(_01880_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26221_ (.A1(net17780),
    .A2(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26222_ (.A1(_02209_),
    .A2(net18628),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26223_ (.A1(_02207_),
    .A2(net19712),
    .A3(_02210_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26224_ (.A1(_02206_),
    .A2(_02211_),
    .A3(net19711),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26225_ (.A1(_02212_),
    .A2(_02202_),
    .B(net20421),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26226_ (.A1(_01997_),
    .A2(net17199),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26227_ (.A1(_02214_),
    .A2(net19703),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26228_ (.A1(net17484),
    .A2(net18160),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26229_ (.A1(_01929_),
    .A2(net17785),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26230_ (.A1(_02216_),
    .A2(_02217_),
    .A3(net19717),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26231_ (.A1(_02215_),
    .A2(net19187),
    .A3(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26232_ (.A1(net17469),
    .A2(net17271),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26233_ (.A1(_01983_),
    .A2(net18618),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26234_ (.A1(_02220_),
    .A2(_02221_),
    .A3(net19717),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26235_ (.A1(_01983_),
    .A2(_01898_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26236_ (.A1(_02223_),
    .A2(_01811_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26237_ (.A1(_02222_),
    .A2(net19711),
    .A3(_02224_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26238_ (.A1(_02219_),
    .A2(_02225_),
    .A3(net20422),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26239_ (.A1(_02213_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26240_ (.A1(_02196_),
    .A2(_02227_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26241_ (.A1(_01897_),
    .A2(_02095_),
    .A3(net17482),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26242_ (.A1(_01806_),
    .A2(net18639),
    .B(net19702),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26243_ (.A1(net18623),
    .A2(net17764),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26244_ (.A1(_02229_),
    .A2(_02230_),
    .B(net19711),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26245_ (.A1(_02228_),
    .A2(_02231_),
    .B(net20421),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26246_ (.A1(net17765),
    .A2(_01750_),
    .B(net18628),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26247_ (.A1(net18623),
    .A2(_15959_[0]),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _26248_ (.A1(_02233_),
    .A2(net19704),
    .A3(_02234_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26249_ (.A1(_01923_),
    .A2(net18160),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26250_ (.A1(net17475),
    .A2(net17784),
    .A3(net18627),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26251_ (.A1(_02236_),
    .A2(_02237_),
    .A3(net19703),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26252_ (.A1(_02235_),
    .A2(_02238_),
    .A3(net19711),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26253_ (.A1(_02239_),
    .A2(_02232_),
    .B(_01848_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26254_ (.A1(net17773),
    .A2(net18636),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26255_ (.A1(_01983_),
    .A2(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26256_ (.A1(_02242_),
    .A2(_02182_),
    .B(net19705),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26257_ (.A1(_01881_),
    .A2(net18623),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _26258_ (.A1(_01746_),
    .A2(_02244_),
    .A3(net19705),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26259_ (.A1(_02245_),
    .A2(net19711),
    .A3(_02243_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26260_ (.A1(net18645),
    .A2(net19722),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26261_ (.A1(_02077_),
    .A2(net18645),
    .B(net19703),
    .C(_02247_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26262_ (.A1(_02241_),
    .A2(_01725_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26263_ (.A1(_01977_),
    .A2(net19716),
    .A3(_02249_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26264_ (.A1(_02248_),
    .A2(_02250_),
    .A3(net19184),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26265_ (.A1(net20421),
    .A2(_02251_),
    .A3(_02246_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26266_ (.A1(_02240_),
    .A2(_02252_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26267_ (.A1(net17781),
    .A2(net18623),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26268_ (.A1(_02229_),
    .A2(_02254_),
    .A3(net17471),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26269_ (.A1(net17987),
    .A2(net18639),
    .B(net19712),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26270_ (.A1(_02197_),
    .A2(_02256_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26271_ (.A1(_02255_),
    .A2(net19711),
    .A3(_02257_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26272_ (.A1(_02241_),
    .A2(net18155),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26273_ (.A1(_02259_),
    .A2(net19704),
    .A3(_02056_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26274_ (.A1(_01757_),
    .A2(_02208_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26275_ (.A1(_02261_),
    .A2(net18645),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26276_ (.A1(net17766),
    .A2(net17783),
    .A3(net18628),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26277_ (.A1(_02262_),
    .A2(_02263_),
    .A3(net19712),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26278_ (.A1(_02260_),
    .A2(_02264_),
    .A3(net19184),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26279_ (.A1(_02258_),
    .A2(_02265_),
    .A3(_01740_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26280_ (.A1(_01923_),
    .A2(net470),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26281_ (.A1(_02261_),
    .A2(net18627),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26282_ (.A1(_02267_),
    .A2(_02268_),
    .A3(net19703),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26283_ (.A1(_02066_),
    .A2(net19703),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26284_ (.A1(_02270_),
    .A2(_02096_),
    .B(net19711),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26285_ (.A1(_02269_),
    .A2(_02271_),
    .B(_01740_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26286_ (.A1(_01981_),
    .A2(_02207_),
    .A3(net19712),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26287_ (.A1(_02043_),
    .A2(_01855_),
    .A3(net19705),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26288_ (.A1(_02273_),
    .A2(net19711),
    .A3(_02274_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26289_ (.A1(_02272_),
    .A2(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26290_ (.A1(_02266_),
    .A2(_02276_),
    .A3(_01848_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26291_ (.A1(_02277_),
    .A2(_02253_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _26292_ (.I(\sa30_sub[7] ),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26293_ (.A1(_02278_),
    .A2(\sa30_sub[0] ),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26294_ (.A1(_11190_),
    .A2(net21286),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26295_ (.A1(_02279_),
    .A2(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26296_ (.A1(_02281_),
    .A2(net21045),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26297_ (.A1(_11190_),
    .A2(_02278_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26298_ (.A1(\sa30_sub[0] ),
    .A2(\sa30_sub[7] ),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26299_ (.A1(_02283_),
    .A2(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26300_ (.A1(_02285_),
    .A2(net21295),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26301_ (.A1(_02282_),
    .A2(_02286_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26302_ (.A1(\sa11_sr[1] ),
    .A2(\sa01_sr[1] ),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26303_ (.A1(_02288_),
    .A2(_14317_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26304_ (.A1(_11215_),
    .A2(_14327_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26305_ (.A1(_02289_),
    .A2(_02290_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26306_ (.A1(_02291_),
    .A2(_02287_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26307_ (.A1(_02288_),
    .A2(_14327_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26308_ (.A1(_11215_),
    .A2(_14317_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26309_ (.A1(_02293_),
    .A2(_02294_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26310_ (.A1(_02282_),
    .A2(_02286_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26311_ (.A1(_02295_),
    .A2(_02296_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26312_ (.A1(_02292_),
    .A2(_02297_),
    .B(net21493),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26313_ (.I(\text_in_r[73] ),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26314_ (.A1(_02299_),
    .A2(net21493),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26315_ (.A1(_02298_),
    .A2(_02300_),
    .B(net21182),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26316_ (.A1(_02292_),
    .A2(_02297_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26317_ (.A1(net21072),
    .A2(_02302_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26318_ (.I(_02300_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26319_ (.A1(_02303_),
    .A2(_07833_),
    .A3(_02304_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26320_ (.A1(_02301_),
    .A2(_02305_),
    .ZN(_15971_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26321_ (.A1(_11149_),
    .A2(_11166_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26322_ (.A1(net21468),
    .A2(net21410),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26323_ (.A1(_02306_),
    .A2(_02307_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26324_ (.A1(net20981),
    .A2(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26325_ (.A1(_02306_),
    .A2(net21347),
    .A3(_02307_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26326_ (.A1(_02309_),
    .A2(_02310_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26327_ (.A1(net20871),
    .A2(_02311_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26328_ (.A1(net690),
    .A2(_02310_),
    .A3(net20872),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26329_ (.A1(_02313_),
    .A2(_02312_),
    .B(net21493),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26330_ (.I(\text_in_r[72] ),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26331_ (.A1(_02315_),
    .A2(net21493),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26332_ (.A1(net20217),
    .A2(net20932),
    .B(net21183),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26333_ (.A1(_02312_),
    .A2(_02313_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26334_ (.A1(_10378_),
    .A2(_02318_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26335_ (.I(_02316_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26336_ (.A1(net21108),
    .A2(net19997),
    .A3(net20870),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26337_ (.A1(_02317_),
    .A2(_02321_),
    .ZN(_15976_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26338_ (.A1(_11222_),
    .A2(_11224_),
    .A3(net21463),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26339_ (.A1(_11223_),
    .A2(_11221_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26340_ (.A1(\sa11_sr[2] ),
    .A2(\sa30_sub[2] ),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26341_ (.A1(_02323_),
    .A2(_11250_),
    .A3(_02324_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26342_ (.A1(_02322_),
    .A2(_02325_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26343_ (.A1(_02326_),
    .A2(net21049),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26344_ (.A1(_02322_),
    .A2(net20869),
    .A3(net20909),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26345_ (.A1(_02327_),
    .A2(_02328_),
    .B(net21493),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26346_ (.I(\text_in_r[74] ),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26347_ (.A1(_02330_),
    .A2(net21496),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26348_ (.A1(_02329_),
    .A2(_02331_),
    .B(_07839_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26349_ (.A1(_02327_),
    .A2(_02328_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26350_ (.A1(_02333_),
    .A2(net21071),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26351_ (.I(_02331_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26352_ (.A1(_02334_),
    .A2(net21207),
    .A3(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26353_ (.A1(_02332_),
    .A2(_02336_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output284 (.I(net284),
    .Z(text_out[121]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26355_ (.A1(_02298_),
    .A2(_02300_),
    .B(_07833_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26356_ (.A1(_02303_),
    .A2(net21182),
    .A3(_02304_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26357_ (.A1(_02338_),
    .A2(_02339_),
    .ZN(_15966_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26358_ (.A1(_02329_),
    .A2(_02331_),
    .B(net21207),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26359_ (.A1(_02334_),
    .A2(_07839_),
    .A3(_02335_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26360_ (.A1(_02340_),
    .A2(_02341_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output283 (.I(net283),
    .Z(text_out[120]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output282 (.I(net282),
    .Z(text_out[11]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26363_ (.A1(net19696),
    .A2(_15969_[0]),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _26364_ (.I(_02344_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26365_ (.A1(_11266_),
    .A2(_14400_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26366_ (.A1(\sa11_sr[3] ),
    .A2(\sa01_sr[3] ),
    .ZN(_02347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26367_ (.A1(_02346_),
    .A2(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26368_ (.I(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26369_ (.A1(_11221_),
    .A2(net20968),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26370_ (.A1(net21293),
    .A2(net21285),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26371_ (.A1(_02351_),
    .A2(_02350_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26372_ (.A1(_02349_),
    .A2(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26373_ (.I(_02352_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26374_ (.A1(_02348_),
    .A2(_02354_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26375_ (.A1(_02355_),
    .A2(_02353_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26376_ (.A1(net21291),
    .A2(_14393_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26377_ (.A1(_02357_),
    .A2(_02356_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26378_ (.A1(_11259_),
    .A2(_14393_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26379_ (.A1(_02353_),
    .A2(_02355_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26380_ (.A1(_02360_),
    .A2(_02359_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26381_ (.A1(_02358_),
    .A2(_02361_),
    .A3(net21068),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26382_ (.A1(net21497),
    .A2(\text_in_r[75] ),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26383_ (.A1(_02363_),
    .A2(_02362_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26384_ (.A1(_02364_),
    .A2(net21206),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26385_ (.A1(_02362_),
    .A2(_07843_),
    .A3(_02363_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26386_ (.A1(_02365_),
    .A2(_02366_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output281 (.I(net281),
    .Z(text_out[119]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output280 (.I(net280),
    .Z(text_out[118]));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26389_ (.A1(\sa30_sub[3] ),
    .A2(net21285),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26390_ (.A1(_11342_),
    .A2(_02370_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26391_ (.I(_02370_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26392_ (.A1(_02372_),
    .A2(_11341_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26393_ (.A1(_02371_),
    .A2(_02373_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26394_ (.I(net21290),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26395_ (.A1(_02375_),
    .A2(_14419_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26396_ (.A1(_02374_),
    .A2(_02376_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26397_ (.A1(_02374_),
    .A2(_02376_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26398_ (.A1(_02377_),
    .A2(net21071),
    .A3(_02378_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26399_ (.A1(net21497),
    .A2(\text_in_r[76] ),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26400_ (.A1(_02379_),
    .A2(_02380_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26401_ (.A1(_02381_),
    .A2(_07849_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26402_ (.A1(_02379_),
    .A2(net21205),
    .A3(_02380_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26403_ (.A1(_02382_),
    .A2(_02383_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output279 (.I(net279),
    .Z(text_out[117]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26405_ (.A1(net17763),
    .A2(net18614),
    .B(net19686),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output278 (.I(net278),
    .Z(text_out[116]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26407_ (.A1(net19175),
    .A2(net19699),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26408_ (.A1(_02364_),
    .A2(_07843_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26409_ (.A1(_02362_),
    .A2(net21206),
    .A3(_02363_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26410_ (.A1(_02390_),
    .A2(_02389_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output277 (.I(net277),
    .Z(text_out[115]));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _26412_ (.A1(_02388_),
    .A2(net691),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26413_ (.A1(_02314_),
    .A2(_02316_),
    .B(_07828_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _26414_ (.A1(_02319_),
    .A2(net21183),
    .A3(_02320_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26415_ (.A1(_02395_),
    .A2(_02394_),
    .ZN(_15965_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26416_ (.A1(net19172),
    .A2(net19699),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26417_ (.A1(_15981_[0]),
    .A2(net19696),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output276 (.I(net276),
    .Z(text_out[114]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26419_ (.A1(net18584),
    .A2(_02397_),
    .A3(net18598),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26420_ (.A1(_02386_),
    .A2(_02393_),
    .A3(_02399_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26421_ (.A1(net19175),
    .A2(net19696),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output275 (.I(net275),
    .Z(text_out[113]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output274 (.I(net274),
    .Z(text_out[112]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output273 (.I(net273),
    .Z(text_out[111]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output272 (.I(net272),
    .Z(text_out[110]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26426_ (.A1(net19699),
    .A2(_15972_[0]),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26427_ (.A1(_02401_),
    .A2(net18614),
    .A3(net18148),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output271 (.I(net271),
    .Z(text_out[10]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _26429_ (.I(_15983_[0]),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26430_ (.A1(_02409_),
    .A2(net19698),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output270 (.I(net270),
    .Z(text_out[109]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26432_ (.A1(net18584),
    .A2(net444),
    .A3(net18593),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26433_ (.A1(_02407_),
    .A2(net19692),
    .A3(_02412_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26434_ (.A1(\sa11_sr[6] ),
    .A2(\sa30_sub[6] ),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26435_ (.A1(_14478_),
    .A2(_02414_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26436_ (.A1(_02415_),
    .A2(net20950),
    .Z(_02416_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26437_ (.A1(_02415_),
    .A2(net20950),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26438_ (.A1(net21496),
    .A2(\text_in_r[78] ),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _26439_ (.A1(_02416_),
    .A2(net21495),
    .A3(_02417_),
    .B(_02418_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26440_ (.A1(_02419_),
    .A2(\u0.w[1][14] ),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26441_ (.A1(_02419_),
    .A2(\u0.w[1][14] ),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26442_ (.A1(_02420_),
    .A2(_02421_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26443_ (.A1(_02400_),
    .A2(_02413_),
    .B(net20418),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _26444_ (.I(_15968_[0]),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26445_ (.A1(net19696),
    .A2(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output269 (.I(net269),
    .Z(text_out[108]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26447_ (.A1(_02425_),
    .A2(net691),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _26448_ (.I(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26449_ (.A1(net19699),
    .A2(net18391),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26450_ (.A1(net688),
    .A2(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26451_ (.A1(net19696),
    .A2(_15967_[0]),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26452_ (.A1(_02431_),
    .A2(net18606),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26453_ (.A1(net19699),
    .A2(_15977_[0]),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26454_ (.A1(_02432_),
    .A2(_02433_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output268 (.I(net268),
    .Z(text_out[107]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26456_ (.A1(_02430_),
    .A2(_02434_),
    .B(net19686),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26457_ (.A1(_02424_),
    .A2(net19699),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26458_ (.A1(_02381_),
    .A2(net21205),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26459_ (.A1(_02379_),
    .A2(_07849_),
    .A3(_02380_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26460_ (.A1(_02438_),
    .A2(_02439_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output267 (.I(net267),
    .Z(text_out[106]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26462_ (.A1(net18596),
    .A2(_02437_),
    .B(net19678),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26463_ (.A1(net19181),
    .A2(net19701),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output266 (.I(net266),
    .Z(text_out[105]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26465_ (.A1(net19696),
    .A2(net18390),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26466_ (.A1(_02443_),
    .A2(net18614),
    .A3(_02445_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26467_ (.A1(_02442_),
    .A2(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26468_ (.A1(_02447_),
    .A2(net20418),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26469_ (.A1(_02436_),
    .A2(_02448_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26470_ (.A1(net21289),
    .A2(_11304_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26471_ (.A1(_02450_),
    .A2(_11379_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26472_ (.A1(_02450_),
    .A2(_11379_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26473_ (.A1(_02451_),
    .A2(_02452_),
    .A3(net21071),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26474_ (.A1(net21496),
    .A2(\text_in_r[77] ),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26475_ (.A1(_02453_),
    .A2(_02454_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _26476_ (.A1(_02455_),
    .A2(net21204),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26477_ (.A1(_02455_),
    .A2(net21204),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26478_ (.A1(_02456_),
    .A2(_02457_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output265 (.I(net265),
    .Z(text_out[104]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output264 (.I(net264),
    .Z(text_out[103]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26481_ (.A1(_02423_),
    .A2(_02449_),
    .B(net19994),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26482_ (.A1(net19175),
    .A2(net19173),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26483_ (.A1(net19178),
    .A2(net19696),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26484_ (.A1(_02462_),
    .A2(_02463_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26485_ (.A1(_02464_),
    .A2(net18589),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26486_ (.A1(_02463_),
    .A2(net18605),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _26487_ (.I(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26488_ (.A1(_02467_),
    .A2(net18576),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output263 (.I(net263),
    .Z(text_out[102]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26490_ (.A1(_02465_),
    .A2(_02468_),
    .A3(net19695),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26491_ (.A1(net19699),
    .A2(_15981_[0]),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26492_ (.A1(_02471_),
    .A2(net450),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26493_ (.A1(net17755),
    .A2(net17757),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output262 (.I(net262),
    .Z(text_out[101]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26495_ (.A1(net19696),
    .A2(_15977_[0]),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26496_ (.A1(_02429_),
    .A2(_02475_),
    .A3(net18589),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26497_ (.A1(_02473_),
    .A2(net19678),
    .A3(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output261 (.I(net261),
    .Z(text_out[100]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26499_ (.A1(_02470_),
    .A2(_02477_),
    .A3(net20417),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26500_ (.A1(net19172),
    .A2(net19696),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26501_ (.A1(net18574),
    .A2(net18149),
    .A3(net18614),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26502_ (.A1(net19700),
    .A2(_02409_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output260 (.I(net260),
    .Z(text_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26504_ (.A1(net17758),
    .A2(net17753),
    .A3(net18598),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output259 (.I(net259),
    .Z(done));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26506_ (.A1(_02481_),
    .A2(_02484_),
    .B(net19683),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _26507_ (.I(_15974_[0]),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26508_ (.A1(_02487_),
    .A2(net19696),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26509_ (.A1(net17752),
    .A2(net18148),
    .A3(net18594),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26510_ (.A1(_02396_),
    .A2(net18605),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input258 (.I(text_in[9]),
    .Z(net258));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26512_ (.A1(_02489_),
    .A2(net18140),
    .B(net19686),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _26513_ (.I(_02422_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input257 (.I(text_in[99]),
    .Z(net257));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26515_ (.A1(_02486_),
    .A2(_02492_),
    .B(_02493_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _26516_ (.I(_02458_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input256 (.I(text_in[98]),
    .Z(net256));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input255 (.I(net563),
    .Z(net255));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26519_ (.A1(_02479_),
    .A2(_02495_),
    .A3(net19676),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _26520_ (.A1(net21285),
    .A2(net20908),
    .A3(net20948),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26521_ (.A1(net21496),
    .A2(\text_in_r[79] ),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26522_ (.A1(_02500_),
    .A2(net21067),
    .B(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _26523_ (.A1(\u0.w[1][15] ),
    .A2(_02502_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input254 (.I(net564),
    .Z(net254));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26525_ (.A1(_02461_),
    .A2(_02499_),
    .A3(net20415),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26526_ (.A1(net19181),
    .A2(net19696),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26527_ (.A1(_02506_),
    .A2(net450),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26528_ (.A1(net19699),
    .A2(net18390),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26529_ (.A1(_02507_),
    .A2(net18139),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26530_ (.A1(net18573),
    .A2(_02433_),
    .A3(net18597),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26531_ (.A1(_02509_),
    .A2(_02510_),
    .B(net19691),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26532_ (.I(_15967_[0]),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26533_ (.A1(net19699),
    .A2(_02512_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _26534_ (.A1(_02513_),
    .A2(_02345_),
    .B(net18609),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26535_ (.A1(_02488_),
    .A2(net18586),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26536_ (.I(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input253 (.I(net555),
    .Z(net253));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26538_ (.A1(_02514_),
    .A2(_02516_),
    .B(net19682),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26539_ (.A1(_02511_),
    .A2(_02518_),
    .B(_02493_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26540_ (.A1(_02345_),
    .A2(net18594),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26541_ (.A1(_02520_),
    .A2(net19686),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26542_ (.A1(net19696),
    .A2(_15972_[0]),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26543_ (.A1(_02433_),
    .A2(net18136),
    .A3(net18614),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26544_ (.A1(_02521_),
    .A2(_02523_),
    .B(_02493_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26545_ (.A1(_02522_),
    .A2(net692),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26546_ (.I(_15979_[0]),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26547_ (.A1(_02526_),
    .A2(net19699),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26548_ (.A1(_02525_),
    .A2(net17749),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26549_ (.A1(net17763),
    .A2(net18614),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26550_ (.A1(_02528_),
    .A2(net19682),
    .A3(_02529_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input252 (.I(net557),
    .Z(net252));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26552_ (.A1(_02524_),
    .A2(_02530_),
    .B(net19995),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26553_ (.A1(_02519_),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26554_ (.A1(net18387),
    .A2(net19699),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26555_ (.I(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26556_ (.A1(_02535_),
    .A2(net449),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26557_ (.A1(_02399_),
    .A2(net19678),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26558_ (.A1(net19696),
    .A2(_15979_[0]),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26559_ (.A1(_02534_),
    .A2(_02538_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26560_ (.A1(_02539_),
    .A2(net449),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26561_ (.A1(_02540_),
    .A2(net19686),
    .A3(net17457),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26562_ (.A1(net17455),
    .A2(_02537_),
    .B(_02541_),
    .C(_02493_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26563_ (.I(_02508_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26564_ (.A1(_02543_),
    .A2(net449),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26565_ (.A1(net18589),
    .A2(_15990_[0]),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26566_ (.A1(_02544_),
    .A2(_02545_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26567_ (.A1(_02546_),
    .A2(net19694),
    .B(_02493_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26568_ (.I(_15972_[0]),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26569_ (.A1(net19696),
    .A2(_02548_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _26570_ (.A1(_02549_),
    .A2(net691),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26571_ (.A1(_02550_),
    .A2(net19678),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26572_ (.A1(_02551_),
    .A2(_02536_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26573_ (.A1(net18583),
    .A2(_02431_),
    .A3(net18591),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26574_ (.A1(net19699),
    .A2(net18389),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26575_ (.A1(_02554_),
    .A2(net691),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26576_ (.A1(_02553_),
    .A2(_02555_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26577_ (.A1(_02552_),
    .A2(_02556_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input251 (.I(text_in[93]),
    .Z(net251));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26579_ (.A1(_02547_),
    .A2(_02557_),
    .B(net19676),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26580_ (.A1(_02542_),
    .A2(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26581_ (.I(_02503_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26582_ (.A1(_02533_),
    .A2(_02560_),
    .A3(net20211),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26583_ (.A1(_02505_),
    .A2(_02562_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26584_ (.A1(_02515_),
    .A2(_02388_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26585_ (.A1(net18575),
    .A2(net18147),
    .A3(net18608),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26586_ (.A1(net17268),
    .A2(net19679),
    .A3(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26587_ (.A1(net19179),
    .A2(net19699),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26588_ (.A1(net18569),
    .A2(net18151),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input250 (.I(text_in[92]),
    .Z(net250));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26590_ (.A1(_02567_),
    .A2(net18608),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26591_ (.A1(net18145),
    .A2(_02437_),
    .A3(net18600),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26592_ (.A1(_02569_),
    .A2(_02570_),
    .A3(net19687),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26593_ (.A1(_02565_),
    .A2(_02571_),
    .A3(_02496_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26594_ (.A1(_02471_),
    .A2(net18587),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26595_ (.A1(_02573_),
    .A2(_02445_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26596_ (.I(_15969_[0]),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26597_ (.A1(net19699),
    .A2(_02575_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26598_ (.A1(net17761),
    .A2(_02576_),
    .A3(net449),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26599_ (.A1(_02574_),
    .A2(net19686),
    .A3(_02577_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26600_ (.A1(net18583),
    .A2(net18150),
    .A3(net18614),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26601_ (.A1(_02579_),
    .A2(net19678),
    .A3(net17457),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26602_ (.A1(_02578_),
    .A2(net19992),
    .A3(_02580_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26603_ (.A1(_02581_),
    .A2(_02572_),
    .B(net20417),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26604_ (.A1(_02480_),
    .A2(net18608),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26605_ (.A1(_02583_),
    .A2(_02429_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26606_ (.A1(_02406_),
    .A2(net692),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26607_ (.I(_02585_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26608_ (.A1(net17454),
    .A2(net18150),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26609_ (.A1(_02584_),
    .A2(_02587_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input249 (.I(net561),
    .Z(net249));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input248 (.I(net596),
    .Z(net248));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26612_ (.A1(_02588_),
    .A2(net19675),
    .B(net19684),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26613_ (.A1(_02467_),
    .A2(net18578),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26614_ (.A1(_02592_),
    .A2(net17268),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26615_ (.A1(_02593_),
    .A2(net19996),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26616_ (.I(_15993_[0]),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26617_ (.A1(net19996),
    .A2(_02595_),
    .A3(net18589),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26618_ (.A1(_02397_),
    .A2(net450),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26619_ (.A1(_02597_),
    .A2(_02433_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26620_ (.A1(_02596_),
    .A2(_02598_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26621_ (.A1(_02599_),
    .A2(net19695),
    .B(net20417),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26622_ (.A1(_02591_),
    .A2(_02594_),
    .B(_02600_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26623_ (.A1(_02582_),
    .A2(_02601_),
    .B(net20413),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26624_ (.A1(_02507_),
    .A2(net18577),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input247 (.I(text_in[8]),
    .Z(net247));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26626_ (.A1(net18593),
    .A2(net19700),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26627_ (.A1(_02605_),
    .A2(net18133),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26628_ (.A1(_02603_),
    .A2(net19680),
    .A3(_02606_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26629_ (.A1(_02488_),
    .A2(net18605),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26630_ (.I(_02608_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26631_ (.A1(net17267),
    .A2(net18570),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26632_ (.A1(_02428_),
    .A2(net18585),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26633_ (.A1(_02610_),
    .A2(_02611_),
    .A3(net19689),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26634_ (.A1(_02607_),
    .A2(_02612_),
    .A3(net19674),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _26635_ (.A1(net17748),
    .A2(net18614),
    .B(net19678),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26636_ (.A1(_02401_),
    .A2(net18596),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _26637_ (.A1(net450),
    .A2(_15997_[0]),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26638_ (.A1(_02615_),
    .A2(_02614_),
    .A3(_02616_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26639_ (.A1(net18135),
    .A2(_02549_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26640_ (.A1(_02618_),
    .A2(net18611),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26641_ (.A1(_02437_),
    .A2(net444),
    .A3(net18593),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26642_ (.A1(_02619_),
    .A2(_02620_),
    .A3(net19681),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26643_ (.A1(_02617_),
    .A2(_02621_),
    .A3(net19991),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26644_ (.A1(_02613_),
    .A2(_02622_),
    .A3(net20417),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26645_ (.A1(net19181),
    .A2(net19178),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26646_ (.A1(net18568),
    .A2(net18572),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input246 (.I(net599),
    .Z(net246));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26648_ (.A1(_02625_),
    .A2(net18600),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26649_ (.A1(net18138),
    .A2(net18608),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26650_ (.A1(_02628_),
    .A2(net18572),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26651_ (.A1(_02627_),
    .A2(_02629_),
    .A3(net19679),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26652_ (.A1(net446),
    .A2(net17760),
    .A3(net18601),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26653_ (.A1(net19696),
    .A2(_02512_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26654_ (.A1(net18569),
    .A2(net17743),
    .A3(net18608),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26655_ (.A1(_02631_),
    .A2(_02633_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26656_ (.A1(_02634_),
    .A2(net19687),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26657_ (.A1(_02630_),
    .A2(_02635_),
    .A3(net19992),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input245 (.I(text_in[88]),
    .Z(net245));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26659_ (.A1(net19696),
    .A2(net18388),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26660_ (.A1(_02638_),
    .A2(net18607),
    .B(net19686),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26661_ (.A1(_02639_),
    .A2(_02574_),
    .B(net19991),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26662_ (.A1(net18595),
    .A2(_02482_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26663_ (.A1(_02641_),
    .A2(_02401_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _26664_ (.I(_15981_[0]),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26665_ (.A1(net19696),
    .A2(_02643_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26666_ (.I(_02644_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26667_ (.A1(_02645_),
    .A2(net18612),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26668_ (.A1(_02642_),
    .A2(net19695),
    .A3(_02646_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26669_ (.A1(_02640_),
    .A2(_02647_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26670_ (.A1(_02636_),
    .A2(_02493_),
    .A3(_02648_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26671_ (.A1(net20212),
    .A2(_02649_),
    .A3(_02623_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26672_ (.A1(_02650_),
    .A2(_02602_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26673_ (.A1(_02549_),
    .A2(net691),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26674_ (.A1(_02651_),
    .A2(net18135),
    .B(net19686),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26675_ (.A1(_02652_),
    .A2(_02509_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26676_ (.I(_02506_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26677_ (.A1(_02654_),
    .A2(_02585_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26678_ (.I(_02482_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26679_ (.A1(_02608_),
    .A2(_02656_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26680_ (.A1(_02655_),
    .A2(_02657_),
    .B(net19690),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26681_ (.A1(_02653_),
    .A2(_02658_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26682_ (.A1(_02659_),
    .A2(net19994),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26683_ (.A1(_02388_),
    .A2(net18614),
    .A3(_02445_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26684_ (.I(_02661_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26685_ (.A1(net18575),
    .A2(_02554_),
    .A3(net18591),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26686_ (.A1(_02662_),
    .A2(_02663_),
    .B(net19689),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26687_ (.A1(net18149),
    .A2(net18614),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26688_ (.A1(_02665_),
    .A2(net19678),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26689_ (.A1(_02573_),
    .A2(net17761),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26690_ (.A1(_02666_),
    .A2(_02667_),
    .B(net19993),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26691_ (.A1(_02664_),
    .A2(_02668_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26692_ (.A1(_02660_),
    .A2(net20417),
    .A3(_02669_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26693_ (.A1(net19699),
    .A2(_15983_[0]),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26694_ (.I(_02671_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26695_ (.A1(net18143),
    .A2(_02672_),
    .B(net19686),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26696_ (.A1(_02388_),
    .A2(net18590),
    .A3(net18134),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26697_ (.A1(_02673_),
    .A2(_02674_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26698_ (.A1(net17760),
    .A2(_02508_),
    .A3(net691),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26699_ (.A1(_02480_),
    .A2(net17749),
    .A3(net18608),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26700_ (.A1(_02676_),
    .A2(_02677_),
    .B(net19688),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26701_ (.A1(_02675_),
    .A2(_02678_),
    .B(net19672),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26702_ (.A1(net19700),
    .A2(net18141),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26703_ (.A1(_02680_),
    .A2(net18593),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26704_ (.A1(_02681_),
    .A2(net18581),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26705_ (.A1(_02682_),
    .A2(net19680),
    .A3(_02540_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26706_ (.A1(net445),
    .A2(net18600),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26707_ (.I(net18575),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26708_ (.A1(_02671_),
    .A2(net18608),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26709_ (.A1(_02684_),
    .A2(_02685_),
    .B(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26710_ (.I(_02538_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26711_ (.A1(_02688_),
    .A2(net18608),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26712_ (.A1(_02689_),
    .A2(net19679),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26713_ (.A1(_02687_),
    .A2(_02690_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26714_ (.A1(_02683_),
    .A2(_02691_),
    .A3(net19992),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26715_ (.A1(_02679_),
    .A2(_02692_),
    .A3(_02493_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26716_ (.A1(_02670_),
    .A2(_02693_),
    .A3(net20416),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26717_ (.A1(_02632_),
    .A2(net691),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26718_ (.A1(_02695_),
    .A2(net19678),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26719_ (.A1(_02428_),
    .A2(net17741),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26720_ (.A1(_02696_),
    .A2(_02697_),
    .B(net19992),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26721_ (.A1(_02575_),
    .A2(_02487_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26722_ (.A1(net19697),
    .A2(_02699_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26723_ (.A1(net17747),
    .A2(net17448),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26724_ (.A1(net17452),
    .A2(_02701_),
    .A3(net19693),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26725_ (.A1(_02698_),
    .A2(_02702_),
    .B(net20213),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26726_ (.A1(net449),
    .A2(_15999_[0]),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26727_ (.A1(_02655_),
    .A2(net19685),
    .A3(_02704_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26728_ (.A1(net450),
    .A2(_15988_[0]),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26729_ (.A1(_02706_),
    .A2(_02665_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26730_ (.I(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26731_ (.A1(_02708_),
    .A2(net19685),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26732_ (.A1(_02705_),
    .A2(net19996),
    .A3(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26733_ (.A1(_02703_),
    .A2(_02710_),
    .B(net20412),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26734_ (.A1(net18571),
    .A2(_02462_),
    .A3(net18589),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26735_ (.A1(_15993_[0]),
    .A2(net18589),
    .B(_02712_),
    .C(net19684),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26736_ (.I(_02513_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26737_ (.A1(_02507_),
    .A2(_02714_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26738_ (.A1(net18139),
    .A2(net18592),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _26739_ (.I(_15977_[0]),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26740_ (.A1(net19697),
    .A2(_02717_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26741_ (.A1(_02716_),
    .A2(_02718_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26742_ (.A1(_02715_),
    .A2(_02719_),
    .B(net19689),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26743_ (.A1(_02713_),
    .A2(_02720_),
    .A3(net19991),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26744_ (.A1(_02388_),
    .A2(net18595),
    .A3(_02480_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26745_ (.A1(_02509_),
    .A2(net19691),
    .A3(net18129),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26746_ (.A1(net18386),
    .A2(net18615),
    .B(net19695),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26747_ (.A1(net17751),
    .A2(net17756),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26748_ (.A1(_02724_),
    .A2(_02725_),
    .B(net19991),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26749_ (.A1(_02723_),
    .A2(_02726_),
    .B(net20417),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26750_ (.A1(_02721_),
    .A2(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26751_ (.A1(_02711_),
    .A2(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26752_ (.A1(_02694_),
    .A2(_02729_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26753_ (.A1(_02586_),
    .A2(_02475_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26754_ (.A1(_02597_),
    .A2(net17756),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26755_ (.A1(_02730_),
    .A2(_02731_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26756_ (.A1(_02732_),
    .A2(net19684),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26757_ (.A1(net17759),
    .A2(net18614),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26758_ (.A1(net19701),
    .A2(_02717_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26759_ (.A1(_02734_),
    .A2(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26760_ (.A1(_02465_),
    .A2(_02736_),
    .A3(net19693),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26761_ (.A1(_02733_),
    .A2(_02737_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26762_ (.A1(_02738_),
    .A2(net20213),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26763_ (.A1(_02681_),
    .A2(net17761),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26764_ (.A1(_02740_),
    .A2(_02661_),
    .A3(net19680),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26765_ (.I(_02566_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26766_ (.A1(net18128),
    .A2(_02718_),
    .B(net18610),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26767_ (.A1(net17743),
    .A2(_02437_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26768_ (.A1(_02744_),
    .A2(net18601),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26769_ (.A1(_02743_),
    .A2(net19689),
    .A3(_02745_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26770_ (.A1(_02741_),
    .A2(_02746_),
    .A3(net20417),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26771_ (.A1(_02739_),
    .A2(net19676),
    .A3(_02747_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26772_ (.A1(net18604),
    .A2(net18614),
    .A3(net18573),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26773_ (.A1(net17456),
    .A2(_02749_),
    .B(_02493_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26774_ (.A1(_02462_),
    .A2(_02566_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26775_ (.A1(_02751_),
    .A2(net18611),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26776_ (.A1(net18604),
    .A2(net18596),
    .A3(net17758),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26777_ (.A1(_02752_),
    .A2(_02753_),
    .A3(net19682),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26778_ (.A1(_02750_),
    .A2(_02754_),
    .B(net19676),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26779_ (.A1(_02527_),
    .A2(net450),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26780_ (.A1(net17445),
    .A2(net18144),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26781_ (.A1(_02642_),
    .A2(_02757_),
    .A3(net19692),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26782_ (.A1(_02752_),
    .A2(net19682),
    .A3(net17745),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26783_ (.A1(_02758_),
    .A2(_02759_),
    .A3(_02493_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26784_ (.A1(_02755_),
    .A2(_02760_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26785_ (.A1(_02748_),
    .A2(_02761_),
    .A3(net20211),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26786_ (.A1(_02553_),
    .A2(net19678),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26787_ (.A1(_02763_),
    .A2(_02603_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26788_ (.A1(_02734_),
    .A2(net17753),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26789_ (.A1(net18583),
    .A2(net18134),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26790_ (.A1(_02766_),
    .A2(net18589),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26791_ (.A1(_02765_),
    .A2(net19686),
    .A3(_02767_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26792_ (.A1(_02764_),
    .A2(_02768_),
    .B(net19673),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26793_ (.A1(_02673_),
    .A2(net19991),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26794_ (.A1(_02527_),
    .A2(net692),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26795_ (.A1(_02771_),
    .A2(_02700_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26796_ (.A1(_02598_),
    .A2(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26797_ (.A1(_02773_),
    .A2(net19684),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26798_ (.A1(_02770_),
    .A2(_02774_),
    .B(net20417),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26799_ (.A1(_02769_),
    .A2(_02775_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26800_ (.A1(_02433_),
    .A2(net18614),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _26801_ (.A1(_02496_),
    .A2(_02654_),
    .A3(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26802_ (.I(_02425_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26803_ (.A1(_02779_),
    .A2(net18614),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26804_ (.A1(_02780_),
    .A2(_02496_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26805_ (.A1(_02778_),
    .A2(_02781_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26806_ (.I(_02521_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26807_ (.I(_02437_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26808_ (.A1(_02458_),
    .A2(net18589),
    .A3(_02784_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26809_ (.A1(_02783_),
    .A2(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26810_ (.A1(_02782_),
    .A2(_02786_),
    .B(_02493_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26811_ (.I(_02490_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26812_ (.A1(_02788_),
    .A2(net17760),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26813_ (.A1(_02641_),
    .A2(_02700_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26814_ (.A1(_02789_),
    .A2(_02790_),
    .A3(net19991),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26815_ (.A1(net17740),
    .A2(net18602),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26816_ (.A1(_02677_),
    .A2(_02496_),
    .A3(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26817_ (.A1(_02791_),
    .A2(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26818_ (.A1(_02794_),
    .A2(net19685),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26819_ (.A1(_02787_),
    .A2(_02795_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26820_ (.A1(_02776_),
    .A2(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26821_ (.A1(_02797_),
    .A2(net20415),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26822_ (.A1(_02762_),
    .A2(_02798_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26823_ (.A1(_02388_),
    .A2(_02463_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26824_ (.A1(_02799_),
    .A2(net18589),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26825_ (.A1(_02800_),
    .A2(_02584_),
    .A3(net19684),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26826_ (.A1(net17443),
    .A2(net19683),
    .A3(_02345_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26827_ (.A1(_02801_),
    .A2(net19672),
    .A3(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26828_ (.A1(_02592_),
    .A2(_02712_),
    .A3(net19684),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26829_ (.A1(net18579),
    .A2(net18568),
    .A3(net18607),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26830_ (.A1(net18579),
    .A2(net18599),
    .A3(_02429_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26831_ (.A1(_02805_),
    .A2(_02806_),
    .A3(net19687),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26832_ (.A1(_02804_),
    .A2(_02807_),
    .A3(net19991),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26833_ (.A1(_02803_),
    .A2(_02808_),
    .A3(net20213),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26834_ (.A1(net18603),
    .A2(net691),
    .A3(net18145),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26835_ (.A1(_02552_),
    .A2(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26836_ (.I(_02657_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26837_ (.A1(net17750),
    .A2(net18603),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26838_ (.A1(_02812_),
    .A2(_02813_),
    .A3(net19690),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26839_ (.A1(_02811_),
    .A2(_02814_),
    .A3(net19994),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26840_ (.A1(_02688_),
    .A2(net18602),
    .B(net19678),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26841_ (.A1(_02543_),
    .A2(net18592),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26842_ (.I(_02817_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26843_ (.A1(_02816_),
    .A2(_02818_),
    .A3(_02540_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26844_ (.A1(_02437_),
    .A2(net17762),
    .A3(net449),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26845_ (.A1(_02528_),
    .A2(net19681),
    .A3(_02820_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26846_ (.A1(_02819_),
    .A2(_02821_),
    .A3(net19676),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26847_ (.A1(_02815_),
    .A2(_02822_),
    .A3(net20418),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26848_ (.A1(_02809_),
    .A2(_02823_),
    .A3(net20211),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26849_ (.A1(_02467_),
    .A2(net17753),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26850_ (.A1(_02825_),
    .A2(net447),
    .B(net19683),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26851_ (.A1(_02432_),
    .A2(_02443_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26852_ (.I(_02563_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26853_ (.A1(_02827_),
    .A2(_02828_),
    .B(net19686),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26854_ (.A1(_02826_),
    .A2(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26855_ (.A1(_02830_),
    .A2(net20214),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26856_ (.A1(_02401_),
    .A2(_02624_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26857_ (.A1(_02832_),
    .A2(net449),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26858_ (.A1(net17443),
    .A2(net18575),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26859_ (.A1(_02833_),
    .A2(_02834_),
    .B(net19683),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26860_ (.A1(_02465_),
    .A2(_02514_),
    .B(net19693),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26861_ (.A1(_02835_),
    .A2(_02836_),
    .B(net20417),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26862_ (.A1(_02831_),
    .A2(_02837_),
    .A3(net19991),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26863_ (.A1(net18614),
    .A2(net18131),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _26864_ (.A1(_02716_),
    .A2(_02839_),
    .A3(net19678),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26865_ (.A1(_02840_),
    .A2(_02493_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _26866_ (.A1(_02550_),
    .A2(net19686),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26867_ (.A1(_02771_),
    .A2(_02401_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26868_ (.A1(net17265),
    .A2(net17264),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26869_ (.A1(_02841_),
    .A2(_02844_),
    .B(net19994),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26870_ (.A1(_02609_),
    .A2(net18139),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26871_ (.A1(_02537_),
    .A2(_02846_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26872_ (.A1(_02576_),
    .A2(net450),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26873_ (.I(_02848_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _26874_ (.A1(_02849_),
    .A2(_02573_),
    .A3(net19683),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26875_ (.A1(_02847_),
    .A2(_02850_),
    .A3(_02493_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26876_ (.A1(_02845_),
    .A2(_02851_),
    .B(net20211),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26877_ (.A1(_02838_),
    .A2(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26878_ (.A1(_02824_),
    .A2(_02853_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _26879_ (.A1(net17760),
    .A2(_02671_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _26880_ (.A1(net17269),
    .A2(_02433_),
    .B1(_02854_),
    .B2(net18614),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26881_ (.A1(_02855_),
    .A2(net19694),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26882_ (.A1(net18589),
    .A2(_02717_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _26883_ (.A1(net17744),
    .A2(_02857_),
    .A3(net19694),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26884_ (.A1(_02858_),
    .A2(net19675),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26885_ (.A1(_02856_),
    .A2(_02859_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26886_ (.A1(net17744),
    .A2(net18149),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26887_ (.A1(net17448),
    .A2(net18589),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26888_ (.A1(_02861_),
    .A2(net19683),
    .A3(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26889_ (.I(net17450),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26890_ (.A1(_02864_),
    .A2(_02614_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26891_ (.A1(_02863_),
    .A2(net19676),
    .A3(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26892_ (.A1(_02860_),
    .A2(net20413),
    .A3(_02866_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26893_ (.A1(_02849_),
    .A2(_02506_),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26894_ (.A1(_02868_),
    .A2(_02817_),
    .B(net19689),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26895_ (.A1(_02686_),
    .A2(net19678),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26896_ (.A1(_02428_),
    .A2(_02714_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26897_ (.A1(_02870_),
    .A2(_02871_),
    .B(net19674),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26898_ (.A1(_02869_),
    .A2(_02872_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26899_ (.A1(net19176),
    .A2(net18589),
    .B(net19686),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26900_ (.A1(_02833_),
    .A2(_02874_),
    .B(net19991),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26901_ (.A1(net17737),
    .A2(net18568),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26902_ (.A1(net17742),
    .A2(_02735_),
    .A3(net18589),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26903_ (.A1(_02876_),
    .A2(_02877_),
    .A3(net19687),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26904_ (.A1(_02875_),
    .A2(_02878_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26905_ (.A1(_02873_),
    .A2(_02879_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26906_ (.A1(_02880_),
    .A2(net20211),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26907_ (.A1(_02867_),
    .A2(_02881_),
    .A3(net20418),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26908_ (.A1(net19699),
    .A2(net18133),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _26909_ (.A1(net17451),
    .A2(net19686),
    .A3(_02883_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _26910_ (.A1(_02884_),
    .A2(net19676),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26911_ (.A1(net17757),
    .A2(net18612),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26912_ (.A1(net17444),
    .A2(net19685),
    .A3(net17441),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26913_ (.A1(_02885_),
    .A2(_02887_),
    .B(net20412),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26914_ (.A1(net17446),
    .A2(net18136),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26915_ (.I(net17739),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26916_ (.A1(_02681_),
    .A2(_02890_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26917_ (.A1(_02889_),
    .A2(_02891_),
    .A3(net19686),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26918_ (.A1(_02641_),
    .A2(net17752),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26919_ (.A1(_02386_),
    .A2(_02893_),
    .A3(_02393_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26920_ (.A1(_02892_),
    .A2(_02894_),
    .A3(net19676),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26921_ (.A1(_02888_),
    .A2(_02895_),
    .B(net20418),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26922_ (.A1(net19173),
    .A2(net18613),
    .B(_02468_),
    .C(net19684),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26923_ (.A1(net17445),
    .A2(net18580),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26924_ (.A1(net17442),
    .A2(net17746),
    .B(_02898_),
    .C(net19694),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26925_ (.A1(_02897_),
    .A2(_02899_),
    .A3(net19677),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26926_ (.A1(net448),
    .A2(net18130),
    .B(net19678),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26927_ (.A1(net17744),
    .A2(net17754),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26928_ (.A1(_02902_),
    .A2(_02901_),
    .B(net19676),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26929_ (.A1(_02583_),
    .A2(net17741),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _26930_ (.A1(_02904_),
    .A2(_02537_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26931_ (.A1(_02903_),
    .A2(_02905_),
    .B(net20211),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26932_ (.A1(_02900_),
    .A2(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26933_ (.A1(_02896_),
    .A2(_02907_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26934_ (.A1(_02882_),
    .A2(_02908_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26935_ (.A1(_02520_),
    .A2(net19678),
    .Z(_02909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26936_ (.A1(_02756_),
    .A2(net444),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26937_ (.A1(_02605_),
    .A2(net18132),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26938_ (.A1(_02909_),
    .A2(net17262),
    .A3(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26939_ (.A1(_02628_),
    .A2(net18575),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26940_ (.A1(_02605_),
    .A2(_02890_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26941_ (.A1(_02816_),
    .A2(_02913_),
    .A3(_02914_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26942_ (.A1(_02912_),
    .A2(_02915_),
    .A3(net19993),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26943_ (.A1(_02832_),
    .A2(net18588),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26944_ (.A1(_15986_[0]),
    .A2(net18385),
    .B(net18607),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26945_ (.A1(_02917_),
    .A2(net19678),
    .A3(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26946_ (.A1(_02605_),
    .A2(net18389),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26947_ (.A1(_02816_),
    .A2(_02920_),
    .A3(net17449),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26948_ (.A1(_02919_),
    .A2(_02921_),
    .A3(net19673),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26949_ (.A1(_02916_),
    .A2(_02922_),
    .A3(net20214),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26950_ (.A1(net17263),
    .A2(net18144),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26951_ (.A1(net17453),
    .A2(net18580),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26952_ (.A1(_02924_),
    .A2(_02925_),
    .A3(net19677),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26953_ (.A1(_02628_),
    .A2(net17447),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26954_ (.A1(net17751),
    .A2(net18569),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26955_ (.A1(_02927_),
    .A2(_02928_),
    .A3(net19992),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26956_ (.A1(_02926_),
    .A2(_02929_),
    .A3(net19678),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26957_ (.A1(_02443_),
    .A2(net18589),
    .A3(net18137),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26958_ (.A1(_02735_),
    .A2(net18589),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26959_ (.A1(_02931_),
    .A2(net19996),
    .A3(_02932_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26960_ (.A1(_02708_),
    .A2(net19675),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26961_ (.A1(_02780_),
    .A2(net19675),
    .B(net19685),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26962_ (.A1(_02933_),
    .A2(_02934_),
    .A3(_02935_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26963_ (.A1(_02930_),
    .A2(_02936_),
    .A3(net20418),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26964_ (.A1(_02923_),
    .A2(_02937_),
    .A3(net20211),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26965_ (.I(_02445_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _26966_ (.A1(net17736),
    .A2(net449),
    .B1(net20216),
    .B2(net20215),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26967_ (.A1(_02940_),
    .A2(net17444),
    .B(net19693),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _26968_ (.A1(_02751_),
    .A2(net18609),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26969_ (.A1(net18581),
    .A2(net18609),
    .A3(_02883_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26970_ (.A1(_02942_),
    .A2(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26971_ (.A1(_02944_),
    .A2(net19674),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26972_ (.A1(_02941_),
    .A2(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _26973_ (.A1(_02616_),
    .A2(net19991),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26974_ (.A1(_02947_),
    .A2(_02481_),
    .B(net19678),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26975_ (.A1(_02410_),
    .A2(net18609),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26976_ (.A1(_02949_),
    .A2(_02742_),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26977_ (.A1(_02942_),
    .A2(net19674),
    .A3(_02950_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26978_ (.A1(_02948_),
    .A2(_02951_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26979_ (.A1(_02946_),
    .A2(_02952_),
    .A3(net20213),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _26980_ (.I(_15987_[0]),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26981_ (.A1(_02954_),
    .A2(net691),
    .B(net19686),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26982_ (.A1(_02955_),
    .A2(_02898_),
    .B(net19991),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26983_ (.A1(net18128),
    .A2(net18610),
    .B(net19680),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26984_ (.A1(_02854_),
    .A2(net18591),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26985_ (.A1(_02957_),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26986_ (.A1(_02956_),
    .A2(_02959_),
    .B(_02493_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26987_ (.A1(_02843_),
    .A2(net17738),
    .B(net19683),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _26988_ (.A1(_02961_),
    .A2(net17266),
    .B(net19994),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26989_ (.A1(_02960_),
    .A2(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26990_ (.A1(_02953_),
    .A2(_02963_),
    .A3(net20414),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26991_ (.A1(_02938_),
    .A2(_02964_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26992_ (.A1(net449),
    .A2(net19178),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26993_ (.A1(_02799_),
    .A2(net449),
    .B(net19686),
    .C(_02965_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _26994_ (.A1(_02472_),
    .A2(net18582),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26995_ (.A1(_02712_),
    .A2(_02967_),
    .A3(net19678),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _26996_ (.A1(_02966_),
    .A2(_02968_),
    .A3(_02496_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _26997_ (.A1(net18613),
    .A2(_02645_),
    .B(_02886_),
    .C(net19678),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _26998_ (.A1(_02525_),
    .A2(_02472_),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _26999_ (.A1(_02939_),
    .A2(net18612),
    .B(net19678),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27000_ (.A1(_02971_),
    .A2(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27001_ (.A1(_02970_),
    .A2(_02973_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27002_ (.A1(_02974_),
    .A2(_02458_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27003_ (.A1(_02969_),
    .A2(_02975_),
    .A3(net20417),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27004_ (.A1(_02789_),
    .A2(net19686),
    .A3(_02620_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27005_ (.A1(_02910_),
    .A2(_02722_),
    .A3(net19678),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27006_ (.A1(_02977_),
    .A2(_02978_),
    .A3(net19991),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27007_ (.A1(_02843_),
    .A2(net19678),
    .A3(_02949_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27008_ (.A1(net18584),
    .A2(net18136),
    .A3(net449),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27009_ (.A1(net18146),
    .A2(net18142),
    .A3(net18602),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27010_ (.A1(_02981_),
    .A2(_02982_),
    .A3(net19686),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27011_ (.A1(_02980_),
    .A2(_02983_),
    .A3(net19673),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27012_ (.A1(_02979_),
    .A2(_02493_),
    .A3(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27013_ (.A1(_02976_),
    .A2(_02985_),
    .A3(net20412),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27014_ (.A1(_02443_),
    .A2(net18590),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27015_ (.A1(_02987_),
    .A2(_02848_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27016_ (.A1(_02988_),
    .A2(net19991),
    .A3(net18146),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27017_ (.A1(_02432_),
    .A2(net18142),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27018_ (.A1(_02433_),
    .A2(_02445_),
    .A3(net18599),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27019_ (.A1(_02990_),
    .A2(_02991_),
    .B(net19991),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27020_ (.A1(_02989_),
    .A2(_02992_),
    .B(net19678),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27021_ (.A1(net18388),
    .A2(net18607),
    .B(_02496_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27022_ (.A1(_02994_),
    .A2(_02917_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27023_ (.A1(_02472_),
    .A2(net18571),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27024_ (.A1(_02772_),
    .A2(_02996_),
    .A3(_02496_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27025_ (.A1(_02995_),
    .A2(_02997_),
    .A3(net19686),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27026_ (.A1(_02993_),
    .A2(_02493_),
    .A3(_02998_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27027_ (.A1(_02842_),
    .A2(_02393_),
    .A3(_02563_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27028_ (.A1(net18131),
    .A2(net18590),
    .B(net19686),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27029_ (.A1(_03001_),
    .A2(_02555_),
    .B(net19991),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27030_ (.A1(_03000_),
    .A2(_03002_),
    .B(_02493_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27031_ (.A1(_02507_),
    .A2(_02566_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27032_ (.A1(_03004_),
    .A2(_02676_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27033_ (.A1(_03005_),
    .A2(net19687),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27034_ (.A1(net18587),
    .A2(_15995_[0]),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27035_ (.A1(_03007_),
    .A2(net19678),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27036_ (.A1(_03008_),
    .A2(_02689_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27037_ (.A1(_02784_),
    .A2(net18615),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27038_ (.A1(_03009_),
    .A2(_03010_),
    .B(_02496_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27039_ (.A1(_03006_),
    .A2(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27040_ (.A1(_03003_),
    .A2(_03012_),
    .B(net20412),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27041_ (.A1(_02999_),
    .A2(_03013_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27042_ (.A1(_02986_),
    .A2(_03014_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27043_ (.I(\sa31_sub[7] ),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27044_ (.A1(_03015_),
    .A2(\sa31_sub[0] ),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27045_ (.A1(_12002_),
    .A2(\sa31_sub[7] ),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27046_ (.A1(_03017_),
    .A2(_03016_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27047_ (.A1(_03018_),
    .A2(net21031),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27048_ (.A1(_12002_),
    .A2(_03015_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27049_ (.A1(\sa31_sub[0] ),
    .A2(\sa31_sub[7] ),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27050_ (.A1(_03020_),
    .A2(_03021_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27051_ (.A1(_03022_),
    .A2(net21283),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27052_ (.A1(_03019_),
    .A2(_03023_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27053_ (.I(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27054_ (.A1(\sa02_sr[1] ),
    .A2(\sa12_sr[1] ),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27055_ (.A1(_03026_),
    .A2(_15064_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27056_ (.A1(_12024_),
    .A2(_15062_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27057_ (.A1(_03027_),
    .A2(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27058_ (.A1(_03025_),
    .A2(_03029_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27059_ (.A1(_15064_),
    .A2(_12024_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27060_ (.A1(_03026_),
    .A2(_15062_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27061_ (.A1(_03031_),
    .A2(_03032_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27062_ (.A1(_03033_),
    .A2(_03024_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27063_ (.A1(_03030_),
    .A2(_03034_),
    .B(net21513),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27064_ (.I(\text_in_r[41] ),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27065_ (.A1(_03036_),
    .A2(net21513),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27066_ (.A1(_03035_),
    .A2(net20931),
    .B(net21156),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27067_ (.A1(_03030_),
    .A2(_03034_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27068_ (.A1(_03039_),
    .A2(net21087),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27069_ (.I(net21156),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27070_ (.I(_03037_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27071_ (.A1(_03040_),
    .A2(_03041_),
    .A3(_03042_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27072_ (.A1(_03043_),
    .A2(_03038_),
    .ZN(_16007_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27073_ (.A1(net649),
    .A2(\sa12_sr[0] ),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27074_ (.A1(net649),
    .A2(\sa12_sr[0] ),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27075_ (.A1(_03044_),
    .A2(_03045_),
    .B(_15059_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27076_ (.I(_03045_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27077_ (.A1(net21457),
    .A2(net21399),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27078_ (.A1(_03047_),
    .A2(net21333),
    .A3(_03048_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27079_ (.A1(_03046_),
    .A2(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27080_ (.A1(_03050_),
    .A2(net20867),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27081_ (.A1(_03046_),
    .A2(_03049_),
    .A3(net20868),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27082_ (.A1(_03051_),
    .A2(_03052_),
    .B(net21512),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27083_ (.I(\text_in_r[40] ),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27084_ (.A1(_03054_),
    .A2(net21512),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27085_ (.A1(_03053_),
    .A2(_03055_),
    .B(net21157),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27086_ (.A1(_03051_),
    .A2(_03052_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27087_ (.A1(_03057_),
    .A2(_10378_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27088_ (.I(net21157),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27089_ (.I(_03055_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27090_ (.A1(_03058_),
    .A2(_03059_),
    .A3(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27091_ (.A1(_03061_),
    .A2(_03056_),
    .ZN(_16012_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27092_ (.A1(_12031_),
    .A2(_12033_),
    .A3(net21452),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27093_ (.A1(_12032_),
    .A2(_12030_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27094_ (.A1(net21395),
    .A2(\sa31_sub[2] ),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27095_ (.A1(_03063_),
    .A2(_12057_),
    .A3(_03064_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27096_ (.A1(_03062_),
    .A2(_03065_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27097_ (.A1(_03066_),
    .A2(net20809),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27098_ (.A1(_03062_),
    .A2(_03065_),
    .A3(net20905),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27099_ (.A1(_03067_),
    .A2(_03068_),
    .B(net21513),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27100_ (.I(\text_in_r[42] ),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27101_ (.A1(_03070_),
    .A2(net21513),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27102_ (.I(net21180),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27103_ (.A1(_03069_),
    .A2(_03071_),
    .B(_03072_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27104_ (.A1(_03067_),
    .A2(_03068_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27105_ (.A1(_03074_),
    .A2(net21087),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27106_ (.I(_03071_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27107_ (.A1(_03075_),
    .A2(net21180),
    .A3(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27108_ (.A1(_03073_),
    .A2(_03077_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input244 (.I(net594),
    .Z(net244));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27110_ (.A1(_03035_),
    .A2(_03037_),
    .B(_03041_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27111_ (.A1(_03040_),
    .A2(net21156),
    .A3(_03042_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27112_ (.A1(_03080_),
    .A2(_03079_),
    .ZN(_16002_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27113_ (.A1(_03069_),
    .A2(_03071_),
    .B(net21180),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27114_ (.A1(_03075_),
    .A2(_03072_),
    .A3(_03076_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27115_ (.A1(_03081_),
    .A2(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input243 (.I(net591),
    .Z(net243));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input242 (.I(net593),
    .Z(net242));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27118_ (.I(_16003_[0]),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27119_ (.A1(net19660),
    .A2(_03085_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27120_ (.A1(\sa31_sub[2] ),
    .A2(net21273),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27121_ (.A1(_03087_),
    .A2(_15131_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27122_ (.A1(_12030_),
    .A2(net20967),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27123_ (.A1(net21282),
    .A2(net21273),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27124_ (.A1(_03089_),
    .A2(_03090_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27125_ (.A1(_15135_),
    .A2(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27126_ (.A1(_03088_),
    .A2(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27127_ (.A1(\sa12_sr[3] ),
    .A2(\sa02_sr[3] ),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27128_ (.A1(_03094_),
    .A2(net21014),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27129_ (.A1(\sa12_sr[3] ),
    .A2(\sa02_sr[3] ),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27130_ (.A1(net21392),
    .A2(\sa02_sr[3] ),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27131_ (.A1(_03096_),
    .A2(_03097_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27132_ (.A1(_03098_),
    .A2(net21280),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27133_ (.A1(_03095_),
    .A2(_03099_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27134_ (.A1(_03093_),
    .A2(_03100_),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27135_ (.A1(_03093_),
    .A2(_03100_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27136_ (.A1(_03101_),
    .A2(net21088),
    .A3(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27137_ (.A1(net21513),
    .A2(\text_in_r[43] ),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27138_ (.A1(_03103_),
    .A2(net21179),
    .A3(_03104_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27139_ (.A1(_03087_),
    .A2(_03098_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27140_ (.A1(_03094_),
    .A2(_03091_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27141_ (.A1(_03106_),
    .A2(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27142_ (.A1(_15135_),
    .A2(net21280),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27143_ (.A1(_15131_),
    .A2(net21014),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27144_ (.A1(_03109_),
    .A2(_03110_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27145_ (.I(_03111_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27146_ (.A1(_03108_),
    .A2(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27147_ (.A1(_03094_),
    .A2(_03091_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27148_ (.A1(_03087_),
    .A2(_03098_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27149_ (.A1(_03114_),
    .A2(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27150_ (.A1(_03116_),
    .A2(_03111_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27151_ (.A1(_03113_),
    .A2(_03117_),
    .A3(net21088),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27152_ (.I(net21179),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27153_ (.A1(net21088),
    .A2(\text_in_r[43] ),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27154_ (.A1(_03118_),
    .A2(_03119_),
    .A3(_03120_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27155_ (.A1(_03105_),
    .A2(_03121_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input241 (.I(net578),
    .Z(net241));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27157_ (.A1(_03086_),
    .A2(net19165),
    .Z(_03124_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _27158_ (.A1(\sa12_sr[4] ),
    .A2(\sa02_sr[4] ),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27159_ (.A1(net21279),
    .A2(net21275),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27160_ (.A1(_03125_),
    .A2(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _27161_ (.A1(net21279),
    .A2(net21275),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27162_ (.A1(_03128_),
    .A2(_12148_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27163_ (.A1(_03127_),
    .A2(_03129_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27164_ (.I(net21278),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27165_ (.A1(_03131_),
    .A2(_15156_),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27166_ (.A1(_03130_),
    .A2(_03132_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27167_ (.A1(net21278),
    .A2(_15156_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27168_ (.A1(_03127_),
    .A2(_03129_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27169_ (.A1(_03134_),
    .A2(_03135_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27170_ (.A1(_03133_),
    .A2(_03136_),
    .A3(net21081),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27171_ (.A1(net21513),
    .A2(\text_in_r[44] ),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27172_ (.A1(_03137_),
    .A2(_03138_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27173_ (.A1(_03139_),
    .A2(net21178),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27174_ (.I(net21178),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27175_ (.A1(_03137_),
    .A2(_03141_),
    .A3(_03138_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27176_ (.A1(_03140_),
    .A2(_03142_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input240 (.I(text_in[83]),
    .Z(net240));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27178_ (.A1(_03124_),
    .A2(net19985),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input239 (.I(net589),
    .Z(net239));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27180_ (.I(_16013_[0]),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27181_ (.A1(net19663),
    .A2(_03147_),
    .Z(_03148_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27182_ (.A1(_03103_),
    .A2(_03119_),
    .A3(_03104_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27183_ (.A1(_03118_),
    .A2(net21179),
    .A3(_03120_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27184_ (.A1(_03149_),
    .A2(_03150_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input238 (.I(net590),
    .Z(net238));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input237 (.I(text_in[80]),
    .Z(net237));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27187_ (.A1(_03148_),
    .A2(net19154),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27188_ (.I(_16004_[0]),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27189_ (.A1(_03155_),
    .A2(_03083_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27190_ (.A1(_03156_),
    .A2(net19160),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _27191_ (.I(_03157_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27192_ (.A1(net19668),
    .A2(net17980),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27193_ (.A1(_03158_),
    .A2(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27194_ (.A1(_03145_),
    .A2(net17261),
    .A3(_03160_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27195_ (.A1(net18564),
    .A2(net19668),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27196_ (.I(_03162_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input236 (.I(text_in[7]),
    .Z(net236));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27198_ (.A1(_03163_),
    .A2(net19151),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27199_ (.I(_03165_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input235 (.I(text_in[79]),
    .Z(net235));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27201_ (.A1(net17433),
    .A2(net19165),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27202_ (.A1(_03155_),
    .A2(net19668),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27203_ (.A1(net19160),
    .A2(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27204_ (.A1(_03168_),
    .A2(net17259),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27205_ (.A1(_03139_),
    .A2(_03141_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27206_ (.A1(_03137_),
    .A2(net21178),
    .A3(_03138_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27207_ (.A1(_03172_),
    .A2(_03173_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input234 (.I(net597),
    .Z(net234));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input233 (.I(text_in[77]),
    .Z(net233));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27210_ (.A1(_03166_),
    .A2(_03171_),
    .B(net19973),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27211_ (.A1(net21277),
    .A2(_15154_),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27212_ (.I(_12187_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27213_ (.A1(_03178_),
    .A2(_03179_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27214_ (.I(net21277),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27215_ (.A1(_03181_),
    .A2(_15154_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27216_ (.A1(_03182_),
    .A2(_12187_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27217_ (.A1(_03180_),
    .A2(_03183_),
    .A3(net21085),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27218_ (.A1(net21507),
    .A2(\text_in_r[45] ),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27219_ (.A1(_03184_),
    .A2(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27220_ (.A1(_03186_),
    .A2(net21177),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27221_ (.A1(_03186_),
    .A2(net21177),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27222_ (.A1(_03187_),
    .A2(_03188_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input232 (.I(net577),
    .Z(net232));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27224_ (.A1(_03161_),
    .A2(_03177_),
    .A3(net20210),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _27225_ (.I(_16012_[0]),
    .ZN(_16001_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27226_ (.A1(net18566),
    .A2(net19148),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27227_ (.A1(net19671),
    .A2(_03083_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27228_ (.A1(_03192_),
    .A2(net19143),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input231 (.I(text_in[75]),
    .Z(net231));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27230_ (.A1(_03194_),
    .A2(net19162),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27231_ (.A1(_03193_),
    .A2(_03151_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27232_ (.I(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27233_ (.A1(_03198_),
    .A2(_03192_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27234_ (.A1(_03196_),
    .A2(_03199_),
    .A3(net19974),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27235_ (.A1(net19663),
    .A2(_16017_[0]),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input230 (.I(net583),
    .Z(net230));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27237_ (.A1(_03201_),
    .A2(net19153),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27238_ (.A1(_03203_),
    .A2(net17434),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input229 (.I(net579),
    .Z(net229));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27240_ (.A1(net19661),
    .A2(net17975),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input228 (.I(net571),
    .Z(net228));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27242_ (.A1(_03159_),
    .A2(_03206_),
    .A3(net19165),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27243_ (.A1(_03204_),
    .A2(net19986),
    .A3(_03208_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _27244_ (.I(_03189_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input227 (.I(net575),
    .Z(net227));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input226 (.I(text_in[70]),
    .Z(net226));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27247_ (.A1(_03200_),
    .A2(_03209_),
    .A3(net19962),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27248_ (.A1(\sa12_sr[6] ),
    .A2(\sa31_sub[6] ),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27249_ (.A1(_15233_),
    .A2(_03214_),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27250_ (.A1(net20946),
    .A2(_03215_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _27251_ (.I0(_03216_),
    .I1(\text_in_r[46] ),
    .S(net21511),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27252_ (.A1(_03217_),
    .A2(\u0.w[2][14] ),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27253_ (.A1(_03217_),
    .A2(\u0.w[2][14] ),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27254_ (.A1(_03218_),
    .A2(_03219_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input225 (.I(text_in[6]),
    .Z(net225));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27256_ (.A1(_03191_),
    .A2(_03213_),
    .A3(net20411),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27257_ (.A1(_03083_),
    .A2(_16005_[0]),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27258_ (.I(_03223_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27259_ (.A1(_03224_),
    .A2(net19149),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27260_ (.A1(_03225_),
    .A2(net19985),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27261_ (.A1(net19148),
    .A2(net19663),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input224 (.I(text_in[69]),
    .Z(net224));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27263_ (.A1(net19660),
    .A2(_16017_[0]),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27264_ (.A1(_03227_),
    .A2(net19160),
    .A3(_03229_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27265_ (.A1(_03226_),
    .A2(_03165_),
    .A3(net17431),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27266_ (.A1(net19667),
    .A2(net17978),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27267_ (.A1(_03232_),
    .A2(net19155),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27268_ (.I(_03233_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27269_ (.A1(net18566),
    .A2(net19656),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input223 (.I(text_in[68]),
    .Z(net223));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27271_ (.A1(_03234_),
    .A2(net18125),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27272_ (.I(_16019_[0]),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27273_ (.A1(net19656),
    .A2(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27274_ (.A1(net18561),
    .A2(net19167),
    .A3(net17428),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27275_ (.A1(_03237_),
    .A2(_03240_),
    .A3(net19977),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27276_ (.A1(_03231_),
    .A2(_03241_),
    .A3(net20206),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27277_ (.A1(net19146),
    .A2(net19659),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27278_ (.A1(_03234_),
    .A2(net18560),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27279_ (.A1(_03078_),
    .A2(_03238_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27280_ (.A1(_03158_),
    .A2(net17427),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input222 (.I(net558),
    .Z(net222));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27282_ (.A1(_03244_),
    .A2(_03246_),
    .A3(net19977),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27283_ (.A1(_03232_),
    .A2(net19168),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _27284_ (.I(_03249_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27285_ (.I(_16010_[0]),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27286_ (.A1(_03083_),
    .A2(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27287_ (.A1(_03250_),
    .A2(net17424),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27288_ (.A1(_03227_),
    .A2(net19154),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27289_ (.A1(_03253_),
    .A2(net19985),
    .A3(net18122),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27290_ (.A1(_03248_),
    .A2(_03255_),
    .A3(net19962),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _27291_ (.I(_03220_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input221 (.I(text_in[66]),
    .Z(net221));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27293_ (.A1(_03242_),
    .A2(_03256_),
    .A3(_03257_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _27294_ (.A1(net21274),
    .A2(net20900),
    .A3(_12190_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27295_ (.A1(net21501),
    .A2(\text_in_r[47] ),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27296_ (.A1(_03260_),
    .A2(net21085),
    .B(_03261_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27297_ (.A1(\u0.w[2][15] ),
    .A2(_03262_),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input220 (.I(net559),
    .Z(net220));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27299_ (.A1(_03222_),
    .A2(_03259_),
    .A3(net20406),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27300_ (.I(_16008_[0]),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27301_ (.A1(_03083_),
    .A2(_03266_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27302_ (.A1(_03267_),
    .A2(net19168),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27303_ (.A1(_03268_),
    .A2(_03154_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27304_ (.A1(_03224_),
    .A2(net19162),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27305_ (.A1(_03270_),
    .A2(net19969),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27306_ (.A1(_03269_),
    .A2(_03271_),
    .B(_03257_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27307_ (.A1(net19657),
    .A2(_16008_[0]),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27308_ (.A1(_03273_),
    .A2(net19168),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27309_ (.I(_16015_[0]),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27310_ (.A1(net19667),
    .A2(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27311_ (.A1(_03274_),
    .A2(net17420),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input219 (.I(text_in[64]),
    .Z(net219));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27313_ (.A1(_03277_),
    .A2(net19986),
    .A3(_03225_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input218 (.I(text_in[63]),
    .Z(net218));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27315_ (.A1(_03272_),
    .A2(_03279_),
    .B(net20209),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27316_ (.A1(net19663),
    .A2(_16013_[0]),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27317_ (.I(_03282_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27318_ (.A1(net19671),
    .A2(net19667),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27319_ (.A1(_03283_),
    .A2(_03284_),
    .A3(net19155),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27320_ (.A1(net18567),
    .A2(net19660),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27321_ (.A1(net19667),
    .A2(net17979),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27322_ (.A1(_03286_),
    .A2(_03287_),
    .A3(net19155),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input217 (.I(text_in[62]),
    .Z(net217));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27324_ (.A1(_03285_),
    .A2(_03288_),
    .B(net19975),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27325_ (.A1(net19663),
    .A2(_03085_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input216 (.I(text_in[61]),
    .Z(net216));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27327_ (.A1(_03291_),
    .A2(_03224_),
    .B(net19149),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27328_ (.A1(_03252_),
    .A2(net19160),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input215 (.I(text_in[60]),
    .Z(net215));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27330_ (.A1(_03293_),
    .A2(net17257),
    .B(net19985),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27331_ (.A1(_03290_),
    .A2(_03296_),
    .B(net20200),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27332_ (.A1(_03281_),
    .A2(_03297_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27333_ (.A1(_03287_),
    .A2(net19155),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27334_ (.A1(net19155),
    .A2(_16026_[0]),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27335_ (.A1(_03299_),
    .A2(_03300_),
    .B(net19975),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27336_ (.A1(_03301_),
    .A2(net20410),
    .Z(_03302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27337_ (.A1(net19659),
    .A2(_16003_[0]),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27338_ (.A1(_03227_),
    .A2(net19163),
    .A3(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27339_ (.A1(net19667),
    .A2(_16005_[0]),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27340_ (.A1(_03305_),
    .A2(net19163),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27341_ (.A1(_03304_),
    .A2(_03306_),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27342_ (.A1(_03268_),
    .A2(net19985),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27343_ (.A1(net19665),
    .A2(net17977),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27344_ (.I(_03309_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27345_ (.A1(_03310_),
    .A2(net19155),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27346_ (.I(_03311_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27347_ (.A1(_03308_),
    .A2(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27348_ (.A1(_03307_),
    .A2(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input214 (.I(net595),
    .Z(net214));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27350_ (.A1(_03302_),
    .A2(_03314_),
    .B(net19962),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27351_ (.A1(_03230_),
    .A2(net19985),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27352_ (.A1(_03317_),
    .A2(_03311_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27353_ (.A1(net19655),
    .A2(net17974),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27354_ (.A1(net17718),
    .A2(_03319_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27355_ (.A1(_03320_),
    .A2(net19155),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27356_ (.A1(_03321_),
    .A2(net19981),
    .A3(net17260),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27357_ (.A1(_03318_),
    .A2(net20202),
    .A3(_03322_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27358_ (.A1(_03316_),
    .A2(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _27359_ (.I(_03263_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27360_ (.A1(_03298_),
    .A2(_03324_),
    .A3(net20199),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27361_ (.A1(_03265_),
    .A2(_03326_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27362_ (.I(_03170_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27363_ (.A1(_03327_),
    .A2(net17428),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27364_ (.A1(_03313_),
    .A2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27365_ (.A1(_03311_),
    .A2(net19975),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27366_ (.A1(net19155),
    .A2(_16033_[0]),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27367_ (.I(_03235_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input213 (.I(text_in[59]),
    .Z(net213));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27369_ (.A1(_03332_),
    .A2(net19155),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27370_ (.A1(_03330_),
    .A2(_03331_),
    .A3(_03334_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27371_ (.A1(_03329_),
    .A2(_03335_),
    .A3(net20210),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27372_ (.A1(_03158_),
    .A2(net18561),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27373_ (.A1(_03252_),
    .A2(_03151_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27374_ (.I(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27375_ (.A1(net19671),
    .A2(net19667),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27376_ (.A1(_03339_),
    .A2(net19140),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27377_ (.A1(_03337_),
    .A2(_03341_),
    .A3(net19978),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27378_ (.A1(_03286_),
    .A2(net19154),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27379_ (.A1(_03343_),
    .A2(_03192_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27380_ (.A1(net19168),
    .A2(net19667),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input212 (.I(text_in[58]),
    .Z(net212));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27382_ (.A1(_03345_),
    .A2(net17729),
    .B(net19975),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27383_ (.A1(_03344_),
    .A2(_03347_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27384_ (.A1(_03342_),
    .A2(_03348_),
    .A3(net19962),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27385_ (.A1(_03336_),
    .A2(_03349_),
    .A3(net20411),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27386_ (.A1(net18567),
    .A2(net19670),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27387_ (.I(_03351_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input211 (.I(text_in[57]),
    .Z(net211));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27389_ (.A1(_03352_),
    .A2(net19142),
    .B(net19170),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27390_ (.A1(_03299_),
    .A2(net18560),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27391_ (.A1(_03354_),
    .A2(net19989),
    .A3(_03355_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27392_ (.A1(_03340_),
    .A2(net19155),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27393_ (.A1(_03357_),
    .A2(_03086_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27394_ (.A1(_03158_),
    .A2(net17718),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27395_ (.A1(_03358_),
    .A2(_03359_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input210 (.I(text_in[56]),
    .Z(net210));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27397_ (.A1(_03360_),
    .A2(net19981),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27398_ (.A1(_03356_),
    .A2(_03362_),
    .A3(net20205),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27399_ (.A1(net19662),
    .A2(_16010_[0]),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27400_ (.A1(_03364_),
    .A2(net19156),
    .B(net19975),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27401_ (.A1(_03201_),
    .A2(net19160),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27402_ (.A1(net19656),
    .A2(net17979),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27403_ (.A1(_03366_),
    .A2(net17713),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input209 (.I(net556),
    .Z(net209));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27405_ (.A1(_03365_),
    .A2(_03368_),
    .B(net20205),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27406_ (.A1(net17426),
    .A2(net19160),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27407_ (.A1(_03371_),
    .A2(_03235_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _27408_ (.I(_16017_[0]),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27409_ (.A1(net19662),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27410_ (.A1(_03374_),
    .A2(net19167),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27411_ (.A1(_03372_),
    .A2(net19981),
    .A3(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27412_ (.A1(_03370_),
    .A2(_03376_),
    .B(net20408),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27413_ (.A1(_03363_),
    .A2(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27414_ (.A1(_03350_),
    .A2(net20199),
    .A3(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27415_ (.I(_03254_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27416_ (.A1(_03380_),
    .A2(net17731),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27417_ (.A1(_03157_),
    .A2(net19985),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27418_ (.A1(_03381_),
    .A2(_03382_),
    .B(_03210_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27419_ (.I(_16005_[0]),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27420_ (.A1(net19667),
    .A2(_03384_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27421_ (.A1(_03385_),
    .A2(net19155),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27422_ (.A1(_03386_),
    .A2(net17428),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27423_ (.A1(_03368_),
    .A2(_03387_),
    .A3(net19977),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27424_ (.A1(_03383_),
    .A2(_03388_),
    .B(net20408),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27425_ (.A1(_03327_),
    .A2(net17721),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27426_ (.A1(_03390_),
    .A2(_03225_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27427_ (.A1(net19169),
    .A2(_03340_),
    .B(net19975),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27428_ (.A1(_03391_),
    .A2(_03392_),
    .Z(_03393_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27429_ (.A1(_03163_),
    .A2(_03294_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27430_ (.I(_03394_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27431_ (.A1(_03198_),
    .A2(_03159_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27432_ (.A1(_03395_),
    .A2(_03396_),
    .A3(net19986),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27433_ (.A1(_03393_),
    .A2(_03210_),
    .A3(_03397_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27434_ (.A1(_03389_),
    .A2(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27435_ (.A1(_03243_),
    .A2(net19149),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27436_ (.A1(_03400_),
    .A2(_03159_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27437_ (.A1(_03250_),
    .A2(net17732),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27438_ (.A1(_03401_),
    .A2(_03210_),
    .A3(_03402_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27439_ (.A1(_03403_),
    .A2(net19972),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27440_ (.A1(net18567),
    .A2(net19664),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27441_ (.A1(_03198_),
    .A2(_03405_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27442_ (.A1(_03395_),
    .A2(net20205),
    .A3(_03406_),
    .Z(_03407_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27443_ (.I(_16029_[0]),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27444_ (.A1(net20205),
    .A2(_03408_),
    .A3(net19160),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27445_ (.A1(_03229_),
    .A2(net19154),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27446_ (.A1(_03410_),
    .A2(net17725),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27447_ (.A1(_03409_),
    .A2(_03411_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27448_ (.A1(_03412_),
    .A2(net19986),
    .B(_03257_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27449_ (.A1(_03404_),
    .A2(_03407_),
    .B(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27450_ (.A1(_03399_),
    .A2(_03414_),
    .A3(net20406),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27451_ (.A1(_03379_),
    .A2(_03415_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27452_ (.A1(net19663),
    .A2(net17730),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27453_ (.A1(_03158_),
    .A2(net17413),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27454_ (.A1(_03145_),
    .A2(_03417_),
    .B(net20206),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27455_ (.A1(_03384_),
    .A2(net17730),
    .Z(_03419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27456_ (.A1(net19657),
    .A2(_03419_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27457_ (.A1(net17416),
    .A2(net17252),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27458_ (.A1(net17253),
    .A2(_03421_),
    .A3(net19977),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27459_ (.A1(_03418_),
    .A2(_03422_),
    .B(_03257_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27460_ (.I(_03286_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27461_ (.A1(_03424_),
    .A2(_03249_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27462_ (.A1(net19159),
    .A2(_16035_[0]),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27463_ (.A1(_03426_),
    .A2(net19984),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27464_ (.I(_16024_[0]),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27465_ (.A1(net19170),
    .A2(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27466_ (.A1(_03233_),
    .A2(_03429_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _27467_ (.A1(_03425_),
    .A2(_03427_),
    .B1(net17251),
    .B2(net19981),
    .C(net20205),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27468_ (.A1(_03423_),
    .A2(_03431_),
    .B(net20406),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27469_ (.A1(net18120),
    .A2(_03192_),
    .A3(net19165),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _27470_ (.A1(net17971),
    .A2(net19165),
    .B(_03433_),
    .C(net19985),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _27471_ (.A1(_03424_),
    .A2(net19167),
    .A3(_03291_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27472_ (.A1(net19661),
    .A2(net17735),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27473_ (.A1(net17724),
    .A2(_03436_),
    .A3(net19167),
    .Z(_03437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27474_ (.A1(_03435_),
    .A2(_03437_),
    .B(net19979),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27475_ (.A1(_03434_),
    .A2(net20210),
    .A3(_03438_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27476_ (.A1(net18127),
    .A2(net19165),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27477_ (.A1(_03440_),
    .A2(net18560),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27478_ (.A1(net17412),
    .A2(net19977),
    .A3(net17418),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27479_ (.A1(net17972),
    .A2(net19155),
    .B(net19975),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27480_ (.A1(net17421),
    .A2(net17432),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27481_ (.A1(_03443_),
    .A2(_03444_),
    .B(net20210),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27482_ (.A1(_03442_),
    .A2(_03445_),
    .B(net20411),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27483_ (.A1(_03439_),
    .A2(_03446_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27484_ (.A1(_03432_),
    .A2(_03447_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27485_ (.I(_03245_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27486_ (.A1(_03449_),
    .A2(_03338_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27487_ (.A1(_03425_),
    .A2(net17205),
    .B(net19981),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input208 (.I(text_in[54]),
    .Z(net208));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input207 (.I(text_in[53]),
    .Z(net207));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27490_ (.A1(net17719),
    .A2(net17423),
    .A3(net19170),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27491_ (.A1(net17419),
    .A2(net19989),
    .A3(_03454_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27492_ (.A1(_03451_),
    .A2(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27493_ (.A1(_03456_),
    .A2(net20210),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27494_ (.A1(_03405_),
    .A2(net17435),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27495_ (.A1(net19143),
    .A2(net17720),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27496_ (.A1(_03459_),
    .A2(net19162),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _27497_ (.A1(net19165),
    .A2(_03458_),
    .B(_03460_),
    .C(net19977),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27498_ (.A1(net17416),
    .A2(net17429),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27499_ (.A1(net17430),
    .A2(net19987),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27500_ (.A1(_03462_),
    .A2(_03463_),
    .B(net20210),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27501_ (.A1(_03461_),
    .A2(_03464_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27502_ (.A1(_03457_),
    .A2(_03465_),
    .A3(net20411),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27503_ (.A1(_03162_),
    .A2(net19162),
    .A3(net17717),
    .Z(_03467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27504_ (.A1(net19667),
    .A2(net17973),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27505_ (.I(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27506_ (.A1(net18563),
    .A2(_03469_),
    .B(net19975),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27507_ (.A1(_03467_),
    .A2(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27508_ (.A1(_03243_),
    .A2(net19149),
    .A3(net17420),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27509_ (.A1(net17434),
    .A2(net17722),
    .A3(net19162),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27510_ (.A1(_03473_),
    .A2(_03472_),
    .B(net19976),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27511_ (.A1(_03471_),
    .A2(_03474_),
    .B(_03210_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27512_ (.A1(_03416_),
    .A2(net19160),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27513_ (.A1(_03476_),
    .A2(net18126),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27514_ (.A1(_03477_),
    .A2(net19989),
    .A3(_03321_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27515_ (.A1(net17719),
    .A2(net19170),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27516_ (.I(net19144),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27517_ (.A1(_03468_),
    .A2(net19158),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27518_ (.A1(_03479_),
    .A2(_03480_),
    .B(_03481_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27519_ (.I(_03319_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27520_ (.A1(net17411),
    .A2(net19155),
    .B(net19989),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27521_ (.A1(_03482_),
    .A2(_03484_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27522_ (.A1(_03478_),
    .A2(_03485_),
    .A3(net20205),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27523_ (.A1(_03475_),
    .A2(net20203),
    .A3(_03486_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27524_ (.A1(_03466_),
    .A2(_03487_),
    .A3(net20406),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27525_ (.A1(_03448_),
    .A2(_03488_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27526_ (.A1(_03410_),
    .A2(net17432),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27527_ (.A1(_03250_),
    .A2(_03206_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27528_ (.A1(_03489_),
    .A2(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27529_ (.A1(_03491_),
    .A2(net19986),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27530_ (.A1(net17436),
    .A2(net19155),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27531_ (.A1(_03493_),
    .A2(_03148_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27532_ (.A1(_03196_),
    .A2(_03494_),
    .A3(net19974),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27533_ (.A1(_03492_),
    .A2(_03495_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27534_ (.A1(_03496_),
    .A2(net19962),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27535_ (.A1(_03192_),
    .A2(net19140),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27536_ (.A1(_03498_),
    .A2(net19157),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27537_ (.A1(_03499_),
    .A2(net19987),
    .A3(net17425),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27538_ (.A1(_03276_),
    .A2(net19155),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27539_ (.A1(_03501_),
    .A2(net17714),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27540_ (.A1(_03372_),
    .A2(_03502_),
    .A3(net19981),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27541_ (.A1(_03500_),
    .A2(_03503_),
    .A3(net20205),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27542_ (.A1(_03497_),
    .A2(_03504_),
    .A3(net20200),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27543_ (.A1(net18127),
    .A2(net19165),
    .A3(net17435),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27544_ (.A1(_03499_),
    .A2(_03506_),
    .A3(net19986),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27545_ (.A1(net18127),
    .A2(net18559),
    .A3(net19152),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27546_ (.A1(_03508_),
    .A2(net19973),
    .A3(net17259),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27547_ (.A1(_03507_),
    .A2(_03509_),
    .A3(net20210),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27548_ (.A1(_03458_),
    .A2(net19152),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27549_ (.A1(_03476_),
    .A2(net17429),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27550_ (.A1(_03511_),
    .A2(_03512_),
    .A3(net19986),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27551_ (.A1(net19140),
    .A2(_03436_),
    .A3(net19157),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27552_ (.A1(net17440),
    .A2(net17432),
    .A3(net19167),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27553_ (.A1(_03514_),
    .A2(_03515_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27554_ (.A1(_03516_),
    .A2(net19973),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27555_ (.A1(_03513_),
    .A2(net19962),
    .A3(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27556_ (.A1(_03510_),
    .A2(_03518_),
    .A3(net20411),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27557_ (.A1(_03505_),
    .A2(_03519_),
    .A3(net20199),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27558_ (.I(_03344_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27559_ (.A1(_03304_),
    .A2(net19988),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27560_ (.A1(_03521_),
    .A2(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27561_ (.A1(_03227_),
    .A2(_03319_),
    .B(net19153),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27562_ (.A1(_03493_),
    .A2(net17250),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _27563_ (.A1(_03524_),
    .A2(net19985),
    .A3(_03525_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27564_ (.A1(_03523_),
    .A2(_03526_),
    .B(_03210_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27565_ (.A1(_03276_),
    .A2(net19160),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _27566_ (.I(_03528_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27567_ (.A1(_03529_),
    .A2(_03420_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27568_ (.A1(_03411_),
    .A2(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27569_ (.A1(_03531_),
    .A2(net19988),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27570_ (.A1(_03470_),
    .A2(net20205),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27571_ (.A1(_03532_),
    .A2(_03533_),
    .B(net20408),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27572_ (.A1(_03527_),
    .A2(_03534_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27573_ (.A1(net17726),
    .A2(net19155),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _27574_ (.A1(_03210_),
    .A2(_03424_),
    .A3(_03536_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27575_ (.A1(_03168_),
    .A2(net20205),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27576_ (.A1(_03537_),
    .A2(_03538_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _27577_ (.A1(_03210_),
    .A2(net19149),
    .A3(net17432),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27578_ (.I(_03271_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27579_ (.A1(_03540_),
    .A2(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27580_ (.A1(_03539_),
    .A2(_03542_),
    .B(net20204),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27581_ (.A1(_03371_),
    .A2(_03420_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27582_ (.A1(net18562),
    .A2(net19149),
    .A3(net17433),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27583_ (.A1(_03544_),
    .A2(_03545_),
    .A3(net20205),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27584_ (.A1(_03483_),
    .A2(net19165),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27585_ (.A1(_03472_),
    .A2(net19963),
    .A3(_03547_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27586_ (.A1(_03546_),
    .A2(_03548_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27587_ (.A1(_03549_),
    .A2(net19985),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27588_ (.A1(_03543_),
    .A2(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27589_ (.A1(_03535_),
    .A2(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27590_ (.A1(_03552_),
    .A2(net20407),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27591_ (.A1(_03520_),
    .A2(_03553_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27592_ (.A1(_03405_),
    .A2(_03243_),
    .A3(net19166),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27593_ (.A1(_03401_),
    .A2(_03554_),
    .A3(net19986),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27594_ (.A1(_03529_),
    .A2(net19985),
    .A3(_03224_),
    .Z(_03556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27595_ (.A1(_03555_),
    .A2(_03210_),
    .A3(_03556_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27596_ (.A1(_03433_),
    .A2(_03406_),
    .A3(net19986),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27597_ (.A1(net18123),
    .A2(net18118),
    .A3(net19151),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27598_ (.A1(net18123),
    .A2(net19165),
    .A3(_03159_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27599_ (.A1(_03559_),
    .A2(_03560_),
    .A3(net19974),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27600_ (.A1(_03558_),
    .A2(_03561_),
    .A3(net20210),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27601_ (.A1(_03557_),
    .A2(_03562_),
    .A3(net20200),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27602_ (.A1(_03440_),
    .A2(net17721),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27603_ (.A1(_03313_),
    .A2(_03564_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27604_ (.I(_03450_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27605_ (.A1(_03274_),
    .A2(net18127),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27606_ (.A1(_03566_),
    .A2(_03567_),
    .A3(net19973),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27607_ (.A1(_03565_),
    .A2(_03568_),
    .A3(net20210),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27608_ (.A1(_03483_),
    .A2(net19170),
    .B(net19985),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27609_ (.I(_03287_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27610_ (.A1(_03571_),
    .A2(net19168),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27611_ (.I(_03572_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27612_ (.A1(_03570_),
    .A2(_03573_),
    .A3(_03321_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27613_ (.A1(net17432),
    .A2(net17428),
    .A3(net19149),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27614_ (.A1(_03277_),
    .A2(net19986),
    .A3(_03575_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27615_ (.A1(_03574_),
    .A2(_03576_),
    .A3(net19962),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27616_ (.A1(_03569_),
    .A2(_03577_),
    .A3(net20411),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27617_ (.A1(_03563_),
    .A2(_03578_),
    .A3(net20199),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27618_ (.A1(_03235_),
    .A2(_03351_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27619_ (.A1(_03580_),
    .A2(net19150),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27620_ (.A1(_03529_),
    .A2(net19143),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27621_ (.A1(_03581_),
    .A2(_03582_),
    .B(net19988),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27622_ (.A1(_03196_),
    .A2(_03293_),
    .B(net19969),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27623_ (.A1(_03583_),
    .A2(_03584_),
    .B(_03220_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27624_ (.A1(net18127),
    .A2(net17439),
    .B(net19166),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27625_ (.A1(_03586_),
    .A2(net17206),
    .B(net19970),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27626_ (.I(_03345_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27627_ (.A1(_03197_),
    .A2(_03449_),
    .B(_03588_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27628_ (.A1(_03589_),
    .A2(net19986),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27629_ (.A1(_03587_),
    .A2(_03590_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27630_ (.A1(_03591_),
    .A2(_03257_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27631_ (.A1(_03585_),
    .A2(_03592_),
    .A3(net20205),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27632_ (.A1(net17722),
    .A2(net19162),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27633_ (.A1(net19149),
    .A2(net17712),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27634_ (.A1(_03594_),
    .A2(net19985),
    .A3(_03595_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27635_ (.A1(_03596_),
    .A2(_03257_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27636_ (.A1(net17258),
    .A2(net19969),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27637_ (.A1(_03529_),
    .A2(net18123),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27638_ (.A1(_03598_),
    .A2(_03599_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27639_ (.A1(_03597_),
    .A2(_03600_),
    .B(net20209),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27640_ (.A1(_03339_),
    .A2(net17724),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27641_ (.A1(_03317_),
    .A2(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27642_ (.A1(_03366_),
    .A2(_03386_),
    .A3(net19985),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27643_ (.A1(_03603_),
    .A2(net20202),
    .A3(_03604_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27644_ (.A1(_03601_),
    .A2(_03605_),
    .B(_03325_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27645_ (.A1(_03593_),
    .A2(_03606_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27646_ (.A1(_03579_),
    .A2(_03607_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27647_ (.A1(_03374_),
    .A2(net19164),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _27648_ (.A1(net18122),
    .A2(net17716),
    .B1(_03608_),
    .B2(net17437),
    .C(net19980),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27649_ (.A1(net18564),
    .A2(net19163),
    .B(net19975),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27650_ (.A1(_03581_),
    .A2(_03610_),
    .B(net20205),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27651_ (.A1(_03609_),
    .A2(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27652_ (.A1(_03386_),
    .A2(net18119),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27653_ (.A1(_03613_),
    .A2(net17245),
    .B(net19982),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _27654_ (.A1(net17260),
    .A2(net17417),
    .B(_03481_),
    .C(net19989),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27655_ (.A1(_03614_),
    .A2(net20207),
    .A3(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27656_ (.A1(_03612_),
    .A2(_03616_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27657_ (.A1(_03617_),
    .A2(net20409),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27658_ (.A1(net19667),
    .A2(net17729),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27659_ (.A1(net17255),
    .A2(net19975),
    .A3(_03619_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27660_ (.A1(_03620_),
    .A2(net19964),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27661_ (.A1(net17249),
    .A2(net19990),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27662_ (.A1(_03524_),
    .A2(_03622_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27663_ (.A1(_03621_),
    .A2(_03623_),
    .B(net20409),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27664_ (.A1(net17254),
    .A2(net17424),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27665_ (.A1(_03226_),
    .A2(_03625_),
    .A3(_03165_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27666_ (.A1(net17248),
    .A2(net17728),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27667_ (.I(_03419_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27668_ (.A1(_03476_),
    .A2(_03628_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27669_ (.A1(_03627_),
    .A2(_03629_),
    .A3(net19983),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27670_ (.A1(_03626_),
    .A2(_03630_),
    .A3(net19964),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27671_ (.A1(_03624_),
    .A2(_03631_),
    .B(net20406),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27672_ (.A1(_03632_),
    .A2(_03618_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27673_ (.A1(net17436),
    .A2(_03468_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _27674_ (.A1(net17207),
    .A2(net17727),
    .B1(_03634_),
    .B2(net19156),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27675_ (.A1(_03635_),
    .A2(net19982),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27676_ (.A1(net19167),
    .A2(net17735),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _27677_ (.A1(_03410_),
    .A2(net19980),
    .A3(_03637_),
    .B(net20205),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27678_ (.I(_03638_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27679_ (.A1(_03636_),
    .A2(_03639_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27680_ (.A1(_03234_),
    .A2(net17731),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27681_ (.A1(_03420_),
    .A2(net19164),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27682_ (.A1(_03641_),
    .A2(net19985),
    .A3(_03642_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27683_ (.I(_03371_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27684_ (.A1(_03330_),
    .A2(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27685_ (.A1(_03643_),
    .A2(_03645_),
    .A3(net19968),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27686_ (.A1(_03640_),
    .A2(net20409),
    .A3(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27687_ (.A1(net18117),
    .A2(net17413),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27688_ (.A1(net17256),
    .A2(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27689_ (.A1(net17438),
    .A2(net19167),
    .B(net19985),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27690_ (.A1(_03410_),
    .A2(net17427),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27691_ (.A1(_03650_),
    .A2(_03651_),
    .B(net19968),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27692_ (.A1(_03649_),
    .A2(_03652_),
    .B(net20409),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27693_ (.A1(_03501_),
    .A2(_03235_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27694_ (.A1(_03250_),
    .A2(net17436),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27695_ (.A1(net17204),
    .A2(_03655_),
    .A3(net19983),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27696_ (.A1(net19169),
    .A2(net19671),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27697_ (.A1(_03199_),
    .A2(net19990),
    .A3(_03657_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27698_ (.A1(_03656_),
    .A2(_03658_),
    .A3(net19964),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27699_ (.A1(_03653_),
    .A2(_03659_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27700_ (.A1(_03647_),
    .A2(_03660_),
    .A3(net20406),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27701_ (.A1(_03633_),
    .A2(_03661_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27702_ (.A1(net18116),
    .A2(net19164),
    .A3(net17728),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27703_ (.A1(_03662_),
    .A2(net19980),
    .A3(net17261),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27704_ (.A1(net17422),
    .A2(net19141),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27705_ (.A1(net17723),
    .A2(_03420_),
    .A3(net19155),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27706_ (.A1(_03664_),
    .A2(net19989),
    .A3(_03665_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27707_ (.A1(_03663_),
    .A2(_03666_),
    .A3(net20207),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27708_ (.A1(_03250_),
    .A2(net18124),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27709_ (.A1(net17715),
    .A2(net17414),
    .A3(net19158),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27710_ (.A1(_03668_),
    .A2(net19990),
    .A3(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27711_ (.A1(_03430_),
    .A2(_03168_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27712_ (.A1(_03671_),
    .A2(net19984),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27713_ (.A1(_03670_),
    .A2(_03672_),
    .A3(net19967),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27714_ (.A1(_03667_),
    .A2(_03673_),
    .A3(net20409),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27715_ (.A1(net19144),
    .A2(net17723),
    .A3(net19155),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27716_ (.A1(net18558),
    .A2(_03628_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27717_ (.A1(net17246),
    .A2(_03675_),
    .A3(_03676_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27718_ (.A1(net19666),
    .A2(_03373_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27719_ (.A1(net17733),
    .A2(_03678_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27720_ (.A1(_03679_),
    .A2(net19169),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27721_ (.A1(net17420),
    .A2(_03239_),
    .A3(net19155),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27722_ (.A1(_03680_),
    .A2(_03681_),
    .A3(net19990),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27723_ (.A1(_03677_),
    .A2(net20207),
    .A3(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27724_ (.A1(_03580_),
    .A2(net19161),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27725_ (.A1(_16022_[0]),
    .A2(_16031_[0]),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27726_ (.A1(net19150),
    .A2(_03685_),
    .B(net19975),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27727_ (.A1(_03684_),
    .A2(_03686_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27728_ (.A1(net17717),
    .A2(net17720),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27729_ (.A1(_03688_),
    .A2(net19161),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27730_ (.A1(_03689_),
    .A2(net19980),
    .A3(_03124_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27731_ (.A1(_03687_),
    .A2(_03690_),
    .A3(net19968),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27732_ (.A1(_03683_),
    .A2(_03691_),
    .A3(net20201),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27733_ (.A1(_03674_),
    .A2(_03692_),
    .B(net20406),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27734_ (.A1(_03332_),
    .A2(net17247),
    .B(_03536_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27735_ (.A1(_03694_),
    .A2(net19975),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27736_ (.A1(_03454_),
    .A2(net19989),
    .B(_03210_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27737_ (.A1(_03695_),
    .A2(_03696_),
    .B(_03257_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27738_ (.A1(net19155),
    .A2(_16023_[0]),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27739_ (.A1(_03698_),
    .A2(net19985),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27740_ (.A1(_03699_),
    .A2(_03654_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27741_ (.A1(_03634_),
    .A2(net19164),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _27742_ (.A1(_03701_),
    .A2(_03392_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27743_ (.A1(_03700_),
    .A2(_03702_),
    .B(net19964),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27744_ (.A1(_03697_),
    .A2(_03703_),
    .B(_03325_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27745_ (.A1(_03357_),
    .A2(net17428),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27746_ (.A1(_03192_),
    .A2(net19168),
    .A3(_03340_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27747_ (.A1(_03705_),
    .A2(_03706_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27748_ (.A1(_03707_),
    .A2(net19984),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27749_ (.A1(net18124),
    .A2(net19159),
    .A3(_03619_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27750_ (.A1(_03706_),
    .A2(_03709_),
    .A3(net19990),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27751_ (.A1(_03708_),
    .A2(_03710_),
    .A3(net19965),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27752_ (.A1(_03233_),
    .A2(net19142),
    .B(_03331_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27753_ (.A1(_03712_),
    .A2(net19984),
    .B(net19966),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27754_ (.I(_03367_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27755_ (.A1(net17410),
    .A2(net19158),
    .Z(_03715_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27756_ (.A1(_03524_),
    .A2(_03715_),
    .B(net19990),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27757_ (.A1(_03713_),
    .A2(_03716_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27758_ (.A1(_03711_),
    .A2(_03717_),
    .A3(net20201),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27759_ (.A1(_03704_),
    .A2(_03718_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _27760_ (.A1(_03693_),
    .A2(_03719_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27761_ (.I(_03386_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27762_ (.A1(_03405_),
    .A2(net19160),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27763_ (.A1(_03720_),
    .A2(_03721_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27764_ (.A1(_03722_),
    .A2(net20205),
    .A3(net17721),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _27765_ (.A1(_03283_),
    .A2(_03714_),
    .A3(net19155),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27766_ (.A1(net17721),
    .A2(net17734),
    .A3(net19153),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27767_ (.A1(_03724_),
    .A2(_03725_),
    .B(net20205),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27768_ (.A1(_03723_),
    .A2(_03726_),
    .B(net19988),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27769_ (.A1(net17976),
    .A2(net19150),
    .B(_03210_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27770_ (.A1(_03728_),
    .A2(_03684_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27771_ (.A1(_03203_),
    .A2(net18121),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27772_ (.A1(_03730_),
    .A2(_03530_),
    .A3(net19963),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27773_ (.A1(_03729_),
    .A2(_03731_),
    .A3(net19976),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27774_ (.A1(_03727_),
    .A2(net20204),
    .A3(_03732_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27775_ (.A1(_03598_),
    .A2(_03395_),
    .A3(_03165_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27776_ (.A1(net17711),
    .A2(net19162),
    .B(net19969),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27777_ (.A1(_03735_),
    .A2(_03306_),
    .B(net20205),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27778_ (.A1(_03734_),
    .A2(_03736_),
    .B(net20204),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27779_ (.A1(_03380_),
    .A2(net18123),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27780_ (.A1(_03327_),
    .A2(net17714),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27781_ (.A1(_03738_),
    .A2(net19976),
    .A3(_03739_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27782_ (.A1(net17717),
    .A2(net17432),
    .B(net19162),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27783_ (.A1(net19162),
    .A2(_16031_[0]),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _27784_ (.A1(_03741_),
    .A2(net19975),
    .A3(_03742_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27785_ (.A1(_03740_),
    .A2(_03743_),
    .A3(net20208),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27786_ (.A1(_03737_),
    .A2(_03744_),
    .B(net20407),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27787_ (.A1(_03733_),
    .A2(_03745_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27788_ (.A1(net17436),
    .A2(_03678_),
    .B(net19164),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27789_ (.A1(_03747_),
    .A2(_03274_),
    .B(net19975),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27790_ (.A1(_03493_),
    .A2(_03608_),
    .A3(net19985),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27791_ (.A1(_03748_),
    .A2(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27792_ (.A1(_03750_),
    .A2(net20209),
    .B(_03257_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27793_ (.A1(net19146),
    .A2(net19149),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27794_ (.A1(_03554_),
    .A2(net19970),
    .A3(_03752_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27795_ (.A1(_03203_),
    .A2(net18123),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27796_ (.A1(_03433_),
    .A2(_03754_),
    .B(net19971),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27797_ (.A1(_03753_),
    .A2(_03755_),
    .B(_03210_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27798_ (.A1(_03751_),
    .A2(_03756_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27799_ (.A1(_03380_),
    .A2(net17728),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27800_ (.A1(net17415),
    .A2(net17721),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27801_ (.A1(_03758_),
    .A2(net19976),
    .A3(_03759_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27802_ (.A1(net19151),
    .A2(net17428),
    .B(net19969),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27803_ (.A1(_03761_),
    .A2(_03599_),
    .B(net20205),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27804_ (.A1(_03760_),
    .A2(_03762_),
    .B(net20408),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27805_ (.A1(_03441_),
    .A2(net19985),
    .A3(_03681_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27806_ (.A1(_03328_),
    .A2(_03545_),
    .A3(net19976),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27807_ (.A1(_03764_),
    .A2(_03765_),
    .A3(net20208),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27808_ (.A1(_03763_),
    .A2(_03766_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27809_ (.A1(_03757_),
    .A2(_03767_),
    .A3(net20407),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27810_ (.A1(_03746_),
    .A2(_03768_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27811_ (.A1(\sa03_sr[1] ),
    .A2(\sa10_sub[1] ),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27812_ (.A1(_03769_),
    .A2(_00811_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27813_ (.A1(_12833_),
    .A2(_00807_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27814_ (.A1(_03771_),
    .A2(_03770_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27815_ (.I(\sa32_sub[7] ),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27816_ (.A1(_12811_),
    .A2(_03773_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27817_ (.A1(net21271),
    .A2(\sa32_sub[7] ),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27818_ (.A1(_03774_),
    .A2(_03775_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27819_ (.A1(_03776_),
    .A2(net21009),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27820_ (.A1(_03773_),
    .A2(net21271),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27821_ (.A1(_12811_),
    .A2(net21260),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27822_ (.A1(_03778_),
    .A2(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27823_ (.A1(_03780_),
    .A2(net21270),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27824_ (.A1(_03777_),
    .A2(_03781_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27825_ (.A1(_03772_),
    .A2(_03782_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27826_ (.A1(_03769_),
    .A2(_00807_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27827_ (.A1(_12833_),
    .A2(_00811_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27828_ (.A1(_03785_),
    .A2(_03784_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27829_ (.A1(_03780_),
    .A2(net21009),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27830_ (.A1(_03776_),
    .A2(net21270),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27831_ (.A1(_03787_),
    .A2(_03788_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27832_ (.A1(_03789_),
    .A2(_03786_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _27833_ (.A1(_03783_),
    .A2(_03790_),
    .B(net21488),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27834_ (.I(\text_in_r[9] ),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27835_ (.A1(_03792_),
    .A2(net21493),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _27836_ (.A1(net20198),
    .A2(net20930),
    .B(net21136),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27837_ (.A1(_03783_),
    .A2(_03790_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27838_ (.A1(_03795_),
    .A2(_10378_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27839_ (.I(net21136),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27840_ (.I(_03793_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27841_ (.A1(_03796_),
    .A2(_03797_),
    .A3(_03798_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27842_ (.A1(_03799_),
    .A2(_03794_),
    .ZN(_16043_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27843_ (.A1(_12762_),
    .A2(_12780_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27844_ (.A1(\sa03_sr[0] ),
    .A2(\sa10_sub[0] ),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27845_ (.A1(_03800_),
    .A2(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27846_ (.A1(_03802_),
    .A2(net20974),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27847_ (.A1(_03800_),
    .A2(net21315),
    .A3(_03801_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27848_ (.A1(_03803_),
    .A2(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27849_ (.A1(_03805_),
    .A2(_03776_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27850_ (.A1(_03803_),
    .A2(_03804_),
    .A3(_03780_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _27851_ (.A1(_03806_),
    .A2(_03807_),
    .B(net21483),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27852_ (.I(\text_in_r[8] ),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27853_ (.A1(_03809_),
    .A2(net21485),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27854_ (.A1(_03808_),
    .A2(_03810_),
    .B(net21137),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27855_ (.A1(_03806_),
    .A2(_03807_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27856_ (.A1(_03812_),
    .A2(_10378_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27857_ (.I(net21137),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27858_ (.I(_03810_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27859_ (.A1(_03813_),
    .A2(_03814_),
    .A3(_03815_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27860_ (.A1(_03816_),
    .A2(_03811_),
    .ZN(_16048_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27861_ (.A1(_12840_),
    .A2(_12842_),
    .A3(net21440),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27862_ (.A1(_12841_),
    .A2(_12839_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27863_ (.A1(net21381),
    .A2(\sa32_sub[2] ),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27864_ (.A1(_03818_),
    .A2(_12864_),
    .A3(_03819_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27865_ (.A1(_03817_),
    .A2(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27866_ (.A1(_03821_),
    .A2(net20895),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27867_ (.A1(_03817_),
    .A2(_03820_),
    .A3(net20893),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _27868_ (.A1(_03822_),
    .A2(_03823_),
    .B(net21488),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27869_ (.I(\text_in_r[10] ),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27870_ (.A1(_03825_),
    .A2(net21498),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _27871_ (.A1(_03826_),
    .A2(_03824_),
    .B(net21154),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27872_ (.A1(_03822_),
    .A2(_03823_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27873_ (.A1(_03828_),
    .A2(net21091),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27874_ (.I(_03826_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27875_ (.A1(_03830_),
    .A2(net21118),
    .A3(_03829_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27876_ (.A1(_03831_),
    .A2(_03827_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _27877_ (.I(net19649),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input206 (.I(text_in[52]),
    .Z(net206));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27879_ (.A1(_03793_),
    .A2(_03791_),
    .B(_03797_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27880_ (.A1(_03796_),
    .A2(net21136),
    .A3(_03798_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27881_ (.A1(_03834_),
    .A2(_03835_),
    .ZN(_16038_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input205 (.I(text_in[51]),
    .Z(net205));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27883_ (.I(_16039_[0]),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27884_ (.A1(net19651),
    .A2(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27885_ (.A1(_12882_),
    .A2(_00890_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27886_ (.A1(\sa10_sub[3] ),
    .A2(\sa03_sr[3] ),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27887_ (.A1(_03838_),
    .A2(_03839_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27888_ (.I(_03840_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27889_ (.A1(net20997),
    .A2(net20966),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27890_ (.A1(net21267),
    .A2(net21258),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27891_ (.A1(_03842_),
    .A2(_03843_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27892_ (.A1(_03841_),
    .A2(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27893_ (.I(_03844_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27894_ (.A1(_03846_),
    .A2(_03840_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _27895_ (.A1(_03845_),
    .A2(_03847_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27896_ (.A1(net21266),
    .A2(_00881_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27897_ (.A1(_03848_),
    .A2(_03849_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27898_ (.A1(net20993),
    .A2(_00881_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27899_ (.A1(_03845_),
    .A2(_03847_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27900_ (.A1(_03851_),
    .A2(_03852_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27901_ (.A1(_03850_),
    .A2(_03853_),
    .A3(net21090),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27902_ (.A1(net21484),
    .A2(\text_in_r[11] ),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27903_ (.A1(_03854_),
    .A2(_03855_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27904_ (.I(net21153),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27905_ (.A1(_03856_),
    .A2(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27906_ (.A1(_03854_),
    .A2(net21153),
    .A3(_03855_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27907_ (.A1(_03858_),
    .A2(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input204 (.I(text_in[50]),
    .Z(net204));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _27909_ (.A1(_03837_),
    .A2(net18549),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27910_ (.A1(net20971),
    .A2(_00916_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27911_ (.I(_12955_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27912_ (.A1(net21266),
    .A2(net21258),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27913_ (.A1(_03864_),
    .A2(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _27914_ (.A1(net21266),
    .A2(net21258),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27915_ (.A1(_03867_),
    .A2(_12955_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27916_ (.A1(_03866_),
    .A2(_03868_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27917_ (.A1(_03863_),
    .A2(_03869_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27918_ (.A1(_03863_),
    .A2(_03869_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27919_ (.A1(_03870_),
    .A2(net21095),
    .A3(_03871_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27920_ (.A1(net21497),
    .A2(\text_in_r[12] ),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27921_ (.A1(_03872_),
    .A2(_03873_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27922_ (.A1(_03874_),
    .A2(net21152),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27923_ (.I(net21152),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27924_ (.A1(_03872_),
    .A2(_03876_),
    .A3(_03873_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27925_ (.A1(_03875_),
    .A2(_03877_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27926_ (.A1(_03862_),
    .A2(net19640),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _27927_ (.I(_16040_[0]),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27928_ (.A1(_03880_),
    .A2(net19650),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27929_ (.A1(net515),
    .A2(net18549),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _27930_ (.I(_03882_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27931_ (.A1(net19129),
    .A2(net18384),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27932_ (.A1(_03883_),
    .A2(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27933_ (.I(_16049_[0]),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27934_ (.A1(net19132),
    .A2(_03886_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _27935_ (.I(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27936_ (.A1(_03856_),
    .A2(net21153),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27937_ (.A1(_03854_),
    .A2(_03857_),
    .A3(_03855_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27938_ (.A1(_03889_),
    .A2(_03890_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input203 (.I(text_in[4]),
    .Z(net203));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input202 (.I(text_in[49]),
    .Z(net202));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27941_ (.A1(_03888_),
    .A2(net18539),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27942_ (.A1(_03879_),
    .A2(_03885_),
    .A3(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27943_ (.A1(net19126),
    .A2(_03833_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27944_ (.I(_03896_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input201 (.I(text_in[48]),
    .Z(net201));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27946_ (.A1(_03897_),
    .A2(net18543),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27947_ (.I(_03899_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27948_ (.I(_03881_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27949_ (.A1(_03901_),
    .A2(net18543),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27950_ (.A1(net20197),
    .A2(net19961),
    .A3(_03880_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27951_ (.A1(net18549),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27952_ (.A1(_03902_),
    .A2(_03904_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27953_ (.A1(_03874_),
    .A2(_03876_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27954_ (.A1(_03872_),
    .A2(net21152),
    .A3(_03873_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27955_ (.A1(_03906_),
    .A2(_03907_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input200 (.I(text_in[47]),
    .Z(net200));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input199 (.I(text_in[46]),
    .Z(net199));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27958_ (.A1(_03900_),
    .A2(_03905_),
    .B(net19637),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27959_ (.A1(net21262),
    .A2(_00921_),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27960_ (.A1(_03912_),
    .A2(_13004_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27961_ (.A1(_03912_),
    .A2(_13004_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _27962_ (.A1(_03913_),
    .A2(_03914_),
    .A3(net21092),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27963_ (.A1(net21498),
    .A2(\text_in_r[13] ),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27964_ (.A1(_03915_),
    .A2(_03916_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27965_ (.A1(_03917_),
    .A2(\u0.tmp_w[13] ),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _27966_ (.I(\u0.tmp_w[13] ),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27967_ (.A1(_03915_),
    .A2(_03919_),
    .A3(_03916_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27968_ (.A1(_03918_),
    .A2(_03920_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input198 (.I(text_in[45]),
    .Z(net198));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27970_ (.A1(_03895_),
    .A2(_03911_),
    .A3(net19626),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _27971_ (.A1(_03808_),
    .A2(_03810_),
    .B(_03814_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27972_ (.A1(_03813_),
    .A2(net21137),
    .A3(_03815_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27973_ (.A1(_03925_),
    .A2(_03924_),
    .ZN(_16037_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _27974_ (.A1(net19126),
    .A2(net19124),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input197 (.I(text_in[44]),
    .Z(net197));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27976_ (.A1(net19135),
    .A2(net19650),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27977_ (.A1(_03926_),
    .A2(net18525),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input196 (.I(text_in[43]),
    .Z(net196));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27979_ (.A1(_03929_),
    .A2(net18554),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27980_ (.A1(_03928_),
    .A2(net18532),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _27981_ (.I(_03932_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27982_ (.A1(_03933_),
    .A2(net18528),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input195 (.I(text_in[42]),
    .Z(net195));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27984_ (.A1(_03931_),
    .A2(_03934_),
    .A3(net19636),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _27985_ (.A1(net18538),
    .A2(net471),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27986_ (.A1(_03833_),
    .A2(_16053_[0]),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27987_ (.A1(_03937_),
    .A2(net18114),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input194 (.I(text_in[41]),
    .Z(net194));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input193 (.I(text_in[40]),
    .Z(net193));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input192 (.I(text_in[3]),
    .Z(net192));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27991_ (.A1(net19652),
    .A2(net18380),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27992_ (.A1(_03884_),
    .A2(net18554),
    .A3(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27993_ (.A1(_03939_),
    .A2(net19640),
    .A3(_03944_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _27994_ (.I(_03921_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input191 (.I(text_in[39]),
    .Z(net191));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _27996_ (.A1(_03936_),
    .A2(_03945_),
    .A3(net19116),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _27997_ (.A1(\sa10_sub[6] ),
    .A2(\sa32_sub[6] ),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _27998_ (.A1(_03949_),
    .A2(_01000_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _27999_ (.A1(_03949_),
    .A2(_01000_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28000_ (.A1(_03950_),
    .A2(_03951_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28001_ (.A1(net20940),
    .A2(_03952_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28002_ (.A1(_03953_),
    .A2(net21095),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28003_ (.A1(net21095),
    .A2(\text_in_r[14] ),
    .B(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28004_ (.I(\u0.tmp_w[14] ),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28005_ (.A1(_03955_),
    .A2(_03956_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28006_ (.A1(_03955_),
    .A2(_03956_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28007_ (.A1(_03957_),
    .A2(_03958_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input190 (.I(text_in[38]),
    .Z(net190));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28009_ (.A1(_03923_),
    .A2(_03948_),
    .A3(net19954),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28010_ (.I(_16055_[0]),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28011_ (.A1(_03962_),
    .A2(net20197),
    .A3(net19959),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28012_ (.A1(_03883_),
    .A2(net17702),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28013_ (.A1(net20197),
    .A2(net19957),
    .A3(_16044_[0]),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28014_ (.A1(net18532),
    .A2(net18112),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28015_ (.A1(net19123),
    .A2(net19650),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28016_ (.I(_03967_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _28017_ (.A1(_03968_),
    .A2(_03966_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28018_ (.A1(_03964_),
    .A2(_03969_),
    .A3(net19634),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28019_ (.A1(_03965_),
    .A2(net18549),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _28020_ (.I(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28021_ (.I(_16046_[0]),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28022_ (.A1(net19650),
    .A2(net18111),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28023_ (.A1(_03972_),
    .A2(net17699),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28024_ (.A1(_03833_),
    .A2(net19123),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28025_ (.A1(_03976_),
    .A2(net18532),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28026_ (.A1(_03975_),
    .A2(net19640),
    .A3(net18110),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28027_ (.A1(_03970_),
    .A2(_03978_),
    .A3(net19116),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28028_ (.A1(net19650),
    .A2(net18382),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28029_ (.A1(net18108),
    .A2(net18543),
    .B(net19630),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28030_ (.A1(net19650),
    .A2(_16053_[0]),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28031_ (.A1(net18106),
    .A2(net18553),
    .A3(net18521),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28032_ (.A1(_03981_),
    .A2(_03983_),
    .A3(_03899_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28033_ (.A1(net19125),
    .A2(net19650),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input189 (.I(text_in[37]),
    .Z(net189));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28035_ (.A1(net18113),
    .A2(net18535),
    .A3(net18517),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28036_ (.A1(net19650),
    .A2(_03962_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28037_ (.A1(net18519),
    .A2(net18554),
    .A3(net17697),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input188 (.I(text_in[36]),
    .Z(net188));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28039_ (.A1(net19631),
    .A2(_03989_),
    .A3(_03987_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28040_ (.A1(_03984_),
    .A2(net19626),
    .A3(_03991_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _28041_ (.I(_03959_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input187 (.I(text_in[35]),
    .Z(net187));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28043_ (.A1(_03979_),
    .A2(_03992_),
    .A3(net19623),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _28044_ (.A1(net21258),
    .A2(net20892),
    .A3(net20939),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28045_ (.A1(net21489),
    .A2(\text_in_r[15] ),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28046_ (.A1(_03996_),
    .A2(net21092),
    .B(_03997_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28047_ (.A1(\u0.tmp_w[15] ),
    .A2(_03998_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input186 (.I(text_in[34]),
    .Z(net186));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28049_ (.A1(net20403),
    .A2(_03961_),
    .A3(_03995_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input185 (.I(text_in[33]),
    .Z(net185));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28051_ (.A1(_03833_),
    .A2(net18381),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28052_ (.I(_16044_[0]),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28053_ (.A1(net19650),
    .A2(_04004_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28054_ (.A1(_04003_),
    .A2(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28055_ (.A1(_04006_),
    .A2(net18543),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input184 (.I(text_in[32]),
    .Z(net184));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28057_ (.A1(net19651),
    .A2(net18384),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28058_ (.A1(net18521),
    .A2(net18553),
    .A3(_04009_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28059_ (.A1(net19130),
    .A2(net18382),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _28060_ (.A1(_04011_),
    .A2(net18553),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _28061_ (.A1(net19645),
    .A2(net17243),
    .A3(_04010_),
    .A4(_04012_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input183 (.I(text_in[31]),
    .Z(net183));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28063_ (.A1(net20197),
    .A2(_16040_[0]),
    .A3(net19960),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28064_ (.A1(net18532),
    .A2(net18100),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28065_ (.A1(_16062_[0]),
    .A2(net18533),
    .B(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input182 (.I(text_in[30]),
    .Z(net182));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28067_ (.A1(_04017_),
    .A2(net19634),
    .B(net19117),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28068_ (.A1(_04013_),
    .A2(_04019_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28069_ (.A1(net19650),
    .A2(_16044_[0]),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28070_ (.A1(_04021_),
    .A2(net18549),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28071_ (.I(_16051_[0]),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28072_ (.A1(net19957),
    .A2(net20197),
    .A3(_04023_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28073_ (.A1(_04022_),
    .A2(net616),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input181 (.I(text_in[2]),
    .Z(net181));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28075_ (.A1(net18108),
    .A2(net18543),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28076_ (.A1(_04025_),
    .A2(net19640),
    .A3(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28077_ (.A1(_04005_),
    .A2(net18549),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28078_ (.A1(_03980_),
    .A2(net18557),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28079_ (.A1(_04029_),
    .A2(_04030_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input180 (.I(text_in[29]),
    .Z(net180));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28081_ (.A1(_03888_),
    .A2(net18537),
    .B(net19640),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28082_ (.A1(_04031_),
    .A2(_04033_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input179 (.I(text_in[28]),
    .Z(net179));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28084_ (.A1(_04028_),
    .A2(_04034_),
    .A3(net19117),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28085_ (.A1(_04020_),
    .A2(net19954),
    .A3(_04036_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28086_ (.I(_04003_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input178 (.I(text_in[27]),
    .Z(net178));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28088_ (.A1(_04038_),
    .A2(net18541),
    .B(net19630),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28089_ (.A1(_04040_),
    .A2(_03983_),
    .B(net19121),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28090_ (.A1(net19650),
    .A2(net18379),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28091_ (.A1(_04003_),
    .A2(_04042_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28092_ (.A1(_04043_),
    .A2(net18532),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28093_ (.A1(_04044_),
    .A2(net17409),
    .A3(net19639),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28094_ (.A1(_04041_),
    .A2(_04045_),
    .B(net19953),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28095_ (.A1(net20197),
    .A2(net19961),
    .A3(_16049_[0]),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28096_ (.A1(net19135),
    .A2(net19127),
    .B(net18551),
    .C(net18097),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28097_ (.A1(net19136),
    .A2(net19650),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input177 (.I(text_in[26]),
    .Z(net177));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28099_ (.A1(net613),
    .A2(net18532),
    .A3(net18514),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28100_ (.A1(_04048_),
    .A2(net19642),
    .A3(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _28101_ (.I(_03980_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28102_ (.A1(net19130),
    .A2(_03836_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28103_ (.A1(_04053_),
    .A2(_04054_),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28104_ (.A1(_04055_),
    .A2(net18541),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input176 (.I(text_in[25]),
    .Z(net176));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28106_ (.A1(net409),
    .A2(net18553),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28107_ (.A1(_04058_),
    .A2(net19630),
    .A3(_04056_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28108_ (.A1(_04052_),
    .A2(_04059_),
    .A3(net19115),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28109_ (.A1(_04060_),
    .A2(_04046_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _28110_ (.I(_03999_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28111_ (.A1(_04037_),
    .A2(_04061_),
    .A3(net20196),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28112_ (.A1(_04001_),
    .A2(_04063_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input175 (.I(net602),
    .Z(net175));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28114_ (.A1(net18109),
    .A2(net18543),
    .B(net19640),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28115_ (.I(_03904_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28116_ (.A1(_04066_),
    .A2(net18103),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28117_ (.A1(_03833_),
    .A2(net19134),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28118_ (.I(_04068_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28119_ (.A1(_04069_),
    .A2(net18542),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28120_ (.A1(_04065_),
    .A2(_04067_),
    .A3(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28121_ (.A1(net18529),
    .A2(net18552),
    .A3(net17698),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28122_ (.A1(_03884_),
    .A2(net18526),
    .A3(net18540),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28123_ (.A1(_04072_),
    .A2(_04073_),
    .A3(net19647),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28124_ (.A1(_04071_),
    .A2(_04074_),
    .A3(net19118),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28125_ (.A1(net17408),
    .A2(net19640),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28126_ (.A1(net18520),
    .A2(net18541),
    .A3(net18106),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28127_ (.A1(_04076_),
    .A2(_04077_),
    .B(_03946_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _28128_ (.I(_16053_[0]),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28129_ (.A1(net19127),
    .A2(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28130_ (.A1(_04080_),
    .A2(net17708),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28131_ (.A1(_04081_),
    .A2(net18553),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28132_ (.I(_16041_[0]),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28133_ (.A1(net20197),
    .A2(net19958),
    .A3(net18092),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28134_ (.A1(net18532),
    .A2(_04084_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _28135_ (.I(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28136_ (.A1(net17242),
    .A2(net17696),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28137_ (.A1(_04082_),
    .A2(_04087_),
    .A3(net19638),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28138_ (.A1(_04078_),
    .A2(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28139_ (.A1(_04089_),
    .A2(_04075_),
    .B(net19955),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28140_ (.A1(_03982_),
    .A2(_04047_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _28141_ (.A1(_04091_),
    .A2(net18549),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28142_ (.I(_16065_[0]),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28143_ (.A1(net19624),
    .A2(net18549),
    .A3(_04093_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28144_ (.A1(_04092_),
    .A2(_04094_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28145_ (.A1(_04095_),
    .A2(net19633),
    .B(net19953),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28146_ (.A1(_04072_),
    .A2(net19637),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28147_ (.A1(net19136),
    .A2(_03833_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28148_ (.A1(_03933_),
    .A2(net18513),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _28149_ (.A1(_04097_),
    .A2(_04099_),
    .A3(net19118),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28150_ (.A1(_03972_),
    .A2(net18107),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28151_ (.A1(_03884_),
    .A2(net18522),
    .A3(net18543),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28152_ (.A1(_03946_),
    .A2(net19630),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28153_ (.A1(_04101_),
    .A2(_04102_),
    .A3(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _28154_ (.A1(_04096_),
    .A2(_04100_),
    .A3(_04104_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28155_ (.A1(_04090_),
    .A2(_04105_),
    .B(net20403),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28156_ (.A1(_04038_),
    .A2(net18541),
    .B(net19640),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _28157_ (.A1(net18536),
    .A2(_16069_[0]),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _28158_ (.I(_03985_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28159_ (.A1(_04109_),
    .A2(net18541),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28160_ (.A1(_04107_),
    .A2(_04108_),
    .A3(_04110_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28161_ (.A1(_04066_),
    .A2(net17696),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28162_ (.A1(net17243),
    .A2(_04112_),
    .A3(net19646),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28163_ (.A1(_04111_),
    .A2(_04113_),
    .A3(net19626),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28164_ (.A1(net18549),
    .A2(_03833_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28165_ (.A1(_04115_),
    .A2(net18104),
    .B(net19630),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28166_ (.A1(_04049_),
    .A2(net18532),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28167_ (.A1(_04117_),
    .A2(_03926_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28168_ (.A1(_04116_),
    .A2(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28169_ (.A1(_04068_),
    .A2(net18541),
    .A3(net17699),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28170_ (.A1(net18520),
    .A2(net17707),
    .A3(net18554),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28171_ (.A1(_04120_),
    .A2(_04121_),
    .A3(net19635),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28172_ (.A1(_04119_),
    .A2(_04122_),
    .A3(net19116),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28173_ (.A1(_04114_),
    .A2(_04123_),
    .A3(net19955),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28174_ (.A1(net19650),
    .A2(net18381),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28175_ (.A1(_04125_),
    .A2(net18548),
    .B(net19630),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input174 (.I(text_in[23]),
    .Z(net174));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28177_ (.A1(_04126_),
    .A2(_04082_),
    .B(net19626),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28178_ (.A1(net18553),
    .A2(net17701),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _28179_ (.A1(_04109_),
    .A2(_04129_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28180_ (.A1(net19654),
    .A2(_04079_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28181_ (.A1(_04131_),
    .A2(net18546),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28182_ (.A1(_04130_),
    .A2(net19635),
    .A3(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28183_ (.A1(_04128_),
    .A2(_04133_),
    .B(net19953),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28184_ (.A1(_03883_),
    .A2(_04003_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28185_ (.A1(_04068_),
    .A2(net18535),
    .A3(net17710),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28186_ (.A1(_04135_),
    .A2(_04136_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28187_ (.A1(_04137_),
    .A2(net19631),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28188_ (.A1(net19137),
    .A2(net19135),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28189_ (.A1(_04139_),
    .A2(net18522),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28190_ (.A1(_04140_),
    .A2(net18549),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28191_ (.A1(_04016_),
    .A2(_03968_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28192_ (.A1(_04141_),
    .A2(_04142_),
    .A3(net19640),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28193_ (.A1(_04138_),
    .A2(_04143_),
    .A3(net19626),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28194_ (.A1(_04134_),
    .A2(_04144_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28195_ (.A1(_04124_),
    .A2(net20196),
    .A3(_04145_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28196_ (.A1(_04106_),
    .A2(_04146_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28197_ (.A1(net18532),
    .A2(net418),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28198_ (.I(_03963_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _28199_ (.A1(_04148_),
    .A2(_04147_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28200_ (.A1(net19126),
    .A2(_03833_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28201_ (.A1(_03971_),
    .A2(_04150_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input173 (.I(text_in[22]),
    .Z(net173));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28203_ (.A1(_04149_),
    .A2(_04151_),
    .B(net19633),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28204_ (.A1(_04003_),
    .A2(net18557),
    .A3(_04005_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input172 (.I(text_in[21]),
    .Z(net172));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28206_ (.A1(_04051_),
    .A2(_04154_),
    .A3(net19640),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28207_ (.A1(_04153_),
    .A2(_04156_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28208_ (.A1(_04157_),
    .A2(net19624),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28209_ (.A1(_04011_),
    .A2(net18526),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28210_ (.A1(_04159_),
    .A2(net18553),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28211_ (.A1(net18513),
    .A2(net17708),
    .A3(net18547),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28212_ (.A1(_04160_),
    .A2(_04161_),
    .A3(net19630),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28213_ (.A1(_03938_),
    .A2(net18549),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28214_ (.I(net17697),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28215_ (.A1(_04163_),
    .A2(_04164_),
    .B(net19640),
    .C(_03966_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28216_ (.A1(_04162_),
    .A2(_04165_),
    .A3(net19116),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28217_ (.A1(_04158_),
    .A2(_04166_),
    .A3(net19956),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28218_ (.A1(net20197),
    .A2(net19958),
    .A3(net18378),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28219_ (.I(_04168_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28220_ (.A1(_03932_),
    .A2(_04169_),
    .B(net19630),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28221_ (.A1(_03896_),
    .A2(net18549),
    .A3(net18098),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28222_ (.A1(_04170_),
    .A2(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28223_ (.A1(net18522),
    .A2(net18540),
    .A3(_04024_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28224_ (.A1(net17709),
    .A2(net18550),
    .A3(net614),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28225_ (.A1(_04173_),
    .A2(_04174_),
    .B(net19633),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28226_ (.A1(_04172_),
    .A2(_04175_),
    .B(net19120),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28227_ (.A1(net20197),
    .A2(net19958),
    .A3(net18111),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28228_ (.A1(net18555),
    .A2(_04177_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28229_ (.A1(_04178_),
    .A2(net18518),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28230_ (.A1(_04044_),
    .A2(_04179_),
    .A3(net19641),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28231_ (.A1(_04178_),
    .A2(net18524),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28232_ (.A1(net18098),
    .A2(_04168_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28233_ (.A1(_04182_),
    .A2(net18544),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28234_ (.A1(_04181_),
    .A2(_04183_),
    .A3(net19632),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28235_ (.A1(_04180_),
    .A2(_04184_),
    .A3(net19627),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28236_ (.A1(_04176_),
    .A2(_04185_),
    .A3(net19621),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28237_ (.A1(_04167_),
    .A2(_04186_),
    .A3(net20402),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28238_ (.I(_04151_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28239_ (.A1(_16071_[0]),
    .A2(net18532),
    .B(net19640),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28240_ (.A1(_04188_),
    .A2(_04189_),
    .B(_03946_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _28241_ (.A1(net18536),
    .A2(_16060_[0]),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28242_ (.A1(_04191_),
    .A2(net19640),
    .A3(_03966_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input171 (.I(text_in[20]),
    .Z(net171));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28244_ (.A1(_04190_),
    .A2(_04192_),
    .B(net19620),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28245_ (.A1(net17692),
    .A2(net17244),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28246_ (.A1(_04195_),
    .A2(_03879_),
    .B(net19627),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28247_ (.I(_04163_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28248_ (.A1(_04083_),
    .A2(_03973_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28249_ (.A1(net19650),
    .A2(_04198_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28250_ (.A1(_04197_),
    .A2(net17401),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28251_ (.A1(_04200_),
    .A2(net19633),
    .A3(_04092_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28252_ (.A1(_04201_),
    .A2(_04196_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28253_ (.A1(_04202_),
    .A2(_04194_),
    .B(net20402),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28254_ (.A1(_03926_),
    .A2(net18515),
    .A3(net18555),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28255_ (.A1(_04204_),
    .A2(net19640),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28256_ (.A1(net18545),
    .A2(net18091),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28257_ (.A1(_04205_),
    .A2(_04206_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28258_ (.A1(net18515),
    .A2(_04054_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28259_ (.A1(_04208_),
    .A2(net18544),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28260_ (.A1(net19652),
    .A2(_03886_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28261_ (.A1(_04210_),
    .A2(net612),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28262_ (.A1(_04211_),
    .A2(net18549),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28263_ (.A1(_04209_),
    .A2(_04212_),
    .A3(net19632),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28264_ (.A1(_04207_),
    .A2(net19628),
    .A3(_04213_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28265_ (.A1(net18530),
    .A2(net18556),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28266_ (.A1(_04215_),
    .A2(net18523),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28267_ (.A1(_04216_),
    .A2(net19633),
    .A3(_04051_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28268_ (.A1(net18533),
    .A2(_16062_[0]),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28269_ (.A1(net17705),
    .A2(_04022_),
    .B(_04218_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28270_ (.A1(_04219_),
    .A2(net19643),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28271_ (.A1(_04217_),
    .A2(_04220_),
    .A3(net19112),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28272_ (.A1(_04214_),
    .A2(_04221_),
    .A3(net19621),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28273_ (.A1(_04222_),
    .A2(_04203_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28274_ (.A1(_04223_),
    .A2(_04187_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28275_ (.A1(_03972_),
    .A2(_03943_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28276_ (.A1(net18105),
    .A2(net18535),
    .A3(net617),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28277_ (.A1(_04224_),
    .A2(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28278_ (.A1(_04226_),
    .A2(net19640),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28279_ (.A1(_03937_),
    .A2(net17706),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28280_ (.A1(_03931_),
    .A2(_04228_),
    .A3(net19636),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28281_ (.A1(_04227_),
    .A2(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28282_ (.A1(_04230_),
    .A2(net19623),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28283_ (.A1(_04178_),
    .A2(net17696),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28284_ (.A1(net18383),
    .A2(net19653),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28285_ (.A1(net18529),
    .A2(net18541),
    .A3(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28286_ (.A1(_04232_),
    .A2(_04234_),
    .A3(net19640),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28287_ (.A1(_04068_),
    .A2(net18535),
    .A3(_04210_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28288_ (.A1(net17710),
    .A2(net18554),
    .A3(net17704),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28289_ (.A1(_04236_),
    .A2(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28290_ (.A1(_04238_),
    .A2(net19631),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28291_ (.A1(_04235_),
    .A2(_04239_),
    .A3(net19953),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28292_ (.A1(_04231_),
    .A2(net19116),
    .A3(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28293_ (.A1(_03904_),
    .A2(net19630),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28294_ (.A1(net18531),
    .A2(net18546),
    .A3(net18523),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28295_ (.A1(_04242_),
    .A2(_04243_),
    .B(_03993_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28296_ (.A1(net19125),
    .A2(net19134),
    .B(net18525),
    .C(net18535),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28297_ (.A1(net18529),
    .A2(net17708),
    .A3(net18553),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28298_ (.A1(_04245_),
    .A2(_04246_),
    .A3(net19640),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28299_ (.A1(_04244_),
    .A2(_04247_),
    .B(net19118),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28300_ (.A1(_04245_),
    .A2(net19640),
    .A3(net17700),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28301_ (.A1(net18532),
    .A2(_04024_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28302_ (.I(_04250_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28303_ (.A1(net17240),
    .A2(net18086),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28304_ (.A1(_04130_),
    .A2(_04252_),
    .A3(net19635),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28305_ (.A1(_04249_),
    .A2(net19623),
    .A3(_04253_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28306_ (.A1(_04248_),
    .A2(_04254_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28307_ (.A1(_04241_),
    .A2(_04255_),
    .A3(net20196),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28308_ (.A1(_04118_),
    .A2(_04010_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28309_ (.A1(_04257_),
    .A2(net19645),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28310_ (.A1(_03937_),
    .A2(net17701),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28311_ (.A1(_03976_),
    .A2(_04042_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28312_ (.A1(_04260_),
    .A2(net18554),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28313_ (.A1(_04259_),
    .A2(_04261_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28314_ (.A1(_04262_),
    .A2(net19634),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28315_ (.A1(_04263_),
    .A2(net19116),
    .A3(_04258_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28316_ (.A1(_04170_),
    .A2(net19625),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28317_ (.A1(net18549),
    .A2(_04024_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28318_ (.I(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28319_ (.A1(_04267_),
    .A2(net17401),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28320_ (.A1(_04092_),
    .A2(_04268_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28321_ (.A1(_04269_),
    .A2(net19640),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28322_ (.A1(_04265_),
    .A2(_04270_),
    .B(net19953),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28323_ (.A1(_04264_),
    .A2(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28324_ (.A1(_04199_),
    .A2(net18549),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28325_ (.A1(_04273_),
    .A2(_04148_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28326_ (.A1(_03976_),
    .A2(_03881_),
    .A3(net18541),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28327_ (.A1(_04274_),
    .A2(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28328_ (.A1(_04276_),
    .A2(net19115),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28329_ (.I(_04042_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28330_ (.A1(_04278_),
    .A2(net18549),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28331_ (.A1(_04173_),
    .A2(_03946_),
    .A3(_04279_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28332_ (.A1(_04277_),
    .A2(_04280_),
    .B(net19642),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28333_ (.A1(net18096),
    .A2(net18543),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _28334_ (.A1(_04282_),
    .A2(_04150_),
    .A3(_03946_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28335_ (.A1(_03902_),
    .A2(net19624),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28336_ (.A1(_04283_),
    .A2(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28337_ (.I(net618),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28338_ (.A1(net19624),
    .A2(net18549),
    .A3(_04286_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28339_ (.A1(_04030_),
    .A2(net19630),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28340_ (.A1(_04287_),
    .A2(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28341_ (.A1(_04285_),
    .A2(_04289_),
    .B(_03993_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28342_ (.A1(_04281_),
    .A2(_04290_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28343_ (.A1(_04272_),
    .A2(_04291_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28344_ (.A1(_04292_),
    .A2(net20403),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28345_ (.A1(_04256_),
    .A2(_04293_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28346_ (.A1(_04056_),
    .A2(_03931_),
    .B(net19636),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28347_ (.A1(_03985_),
    .A2(_04139_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28348_ (.A1(_04295_),
    .A2(net18532),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28349_ (.A1(net17239),
    .A2(net18527),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28350_ (.A1(_04297_),
    .A2(_04296_),
    .B(net19640),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28351_ (.A1(_04294_),
    .A2(_04298_),
    .B(net19953),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28352_ (.A1(_03933_),
    .A2(net17701),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28353_ (.A1(_04115_),
    .A2(net19630),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28354_ (.A1(_04300_),
    .A2(_04301_),
    .B(net19953),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28355_ (.A1(net18513),
    .A2(net18543),
    .A3(net18103),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28356_ (.A1(_04072_),
    .A2(_04303_),
    .A3(net19630),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28357_ (.A1(_04302_),
    .A2(_04304_),
    .B(_04062_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28358_ (.A1(_04305_),
    .A2(_04299_),
    .B(net19120),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28359_ (.A1(_04007_),
    .A2(net19640),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28360_ (.A1(_04215_),
    .A2(net18103),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28361_ (.A1(_04307_),
    .A2(_04308_),
    .B(_03993_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28362_ (.A1(_04022_),
    .A2(_03896_),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _28363_ (.A1(_04310_),
    .A2(net19640),
    .A3(_04149_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28364_ (.A1(_04309_),
    .A2(_04311_),
    .B(net20402),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28365_ (.A1(net18544),
    .A2(_04208_),
    .B(_04296_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28366_ (.A1(_04313_),
    .A2(net19632),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28367_ (.I(_04099_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28368_ (.A1(_04205_),
    .A2(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28369_ (.A1(_04314_),
    .A2(net19621),
    .A3(_04316_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28370_ (.A1(_04317_),
    .A2(_04312_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28371_ (.A1(_04306_),
    .A2(_04318_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28372_ (.A1(net18543),
    .A2(net18093),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28373_ (.A1(net18555),
    .A2(net18102),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28374_ (.A1(_04320_),
    .A2(_04321_),
    .A3(net19640),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28375_ (.A1(_04322_),
    .A2(_03993_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28376_ (.A1(_04029_),
    .A2(net19630),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28377_ (.A1(net17239),
    .A2(net18518),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28378_ (.A1(_04324_),
    .A2(_04325_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28379_ (.A1(_04323_),
    .A2(_04326_),
    .B(_04062_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28380_ (.I(net18102),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _28381_ (.A1(net17403),
    .A2(net17691),
    .B(_03983_),
    .C(net19640),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28382_ (.A1(_04163_),
    .A2(net19630),
    .A3(net17405),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28383_ (.A1(_04330_),
    .A2(net19953),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28384_ (.A1(_04331_),
    .A2(_04329_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28385_ (.A1(_04327_),
    .A2(_04332_),
    .B(net19627),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28386_ (.A1(_04098_),
    .A2(net18556),
    .A3(net18522),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28387_ (.A1(_04334_),
    .A2(_04102_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28388_ (.A1(net17397),
    .A2(net17694),
    .B(net19640),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _28389_ (.A1(net19648),
    .A2(_04335_),
    .B(_04336_),
    .C(net19953),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28390_ (.A1(_04279_),
    .A2(net19630),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28391_ (.A1(_04328_),
    .A2(net18550),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28392_ (.I(_04339_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28393_ (.A1(_04340_),
    .A2(_04044_),
    .A3(_04338_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28394_ (.A1(_03988_),
    .A2(net18532),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28395_ (.A1(net17394),
    .A2(net17705),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28396_ (.A1(_04025_),
    .A2(_04343_),
    .A3(net19643),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28397_ (.A1(_04341_),
    .A2(_04344_),
    .B(_03993_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28398_ (.A1(_04337_),
    .A2(_04345_),
    .B(_04062_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28399_ (.A1(_04346_),
    .A2(_04333_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28400_ (.A1(_04347_),
    .A2(_04319_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28401_ (.A1(net17698),
    .A2(net18553),
    .A3(net17701),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28402_ (.A1(_03981_),
    .A2(_03899_),
    .A3(_04348_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28403_ (.A1(net18099),
    .A2(net18540),
    .A3(net531),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28404_ (.I(_04198_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28405_ (.A1(net18549),
    .A2(_04177_),
    .A3(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28406_ (.A1(_04350_),
    .A2(_04352_),
    .A3(net19630),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28407_ (.A1(_04349_),
    .A2(net19114),
    .A3(_04353_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28408_ (.I(_03937_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28409_ (.A1(_04261_),
    .A2(net19640),
    .A3(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28410_ (.A1(_03833_),
    .A2(net18104),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28411_ (.A1(net17402),
    .A2(net19630),
    .A3(_04357_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28412_ (.A1(_04356_),
    .A2(net19626),
    .A3(_04358_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28413_ (.A1(_04354_),
    .A2(_04359_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28414_ (.A1(_04360_),
    .A2(net19623),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28415_ (.A1(net17405),
    .A2(net18511),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28416_ (.A1(_04362_),
    .A2(_04339_),
    .B(net19639),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28417_ (.A1(_03883_),
    .A2(_04054_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28418_ (.A1(net18532),
    .A2(_04168_),
    .B(net19630),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28419_ (.A1(_04364_),
    .A2(_04365_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28420_ (.A1(_04363_),
    .A2(net19625),
    .A3(_04366_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28421_ (.A1(net17693),
    .A2(net18551),
    .B(net19640),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28422_ (.I(_03977_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28423_ (.A1(_04369_),
    .A2(net18512),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28424_ (.A1(_04368_),
    .A2(_04370_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28425_ (.A1(net19126),
    .A2(net18550),
    .B(net19630),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28426_ (.A1(_04296_),
    .A2(_04372_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28427_ (.A1(_04371_),
    .A2(_04373_),
    .A3(net19113),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28428_ (.A1(_04367_),
    .A2(_04374_),
    .A3(net19953),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28429_ (.A1(_04361_),
    .A2(_04375_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28430_ (.A1(_04376_),
    .A2(net20196),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28431_ (.A1(_04107_),
    .A2(net17404),
    .B(_03993_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28432_ (.A1(net18105),
    .A2(net18535),
    .A3(net18113),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28433_ (.A1(_04379_),
    .A2(net19640),
    .A3(net17238),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28434_ (.A1(_04378_),
    .A2(_04380_),
    .B(net19626),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28435_ (.A1(_03972_),
    .A2(net17707),
    .Z(_04382_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28436_ (.A1(_04251_),
    .A2(_03985_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28437_ (.A1(_04382_),
    .A2(_04383_),
    .B(net19636),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28438_ (.A1(net18554),
    .A2(net19134),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28439_ (.A1(_03934_),
    .A2(_04385_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28440_ (.A1(_04386_),
    .A2(net19644),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28441_ (.A1(_04384_),
    .A2(_04387_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28442_ (.A1(_04388_),
    .A2(net19623),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28443_ (.A1(_04381_),
    .A2(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28444_ (.A1(_03883_),
    .A2(net18097),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28445_ (.A1(net18086),
    .A2(net18539),
    .A3(net17702),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28446_ (.A1(_04391_),
    .A2(net19634),
    .A3(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28447_ (.A1(net18105),
    .A2(net18532),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28448_ (.A1(net18380),
    .A2(net18537),
    .B(_04394_),
    .C(net19640),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28449_ (.A1(_04393_),
    .A2(_04395_),
    .A3(net19953),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28450_ (.A1(_03888_),
    .A2(net18554),
    .B(net19640),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28451_ (.A1(_04394_),
    .A2(_04148_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28452_ (.A1(_04397_),
    .A2(_04398_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28453_ (.A1(net18524),
    .A2(net18545),
    .A3(net17692),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28454_ (.A1(_03983_),
    .A2(_04400_),
    .A3(net19640),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28455_ (.A1(_04399_),
    .A2(_04401_),
    .A3(net19623),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28456_ (.A1(_04396_),
    .A2(_04402_),
    .A3(net19626),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28457_ (.A1(_04390_),
    .A2(_04403_),
    .A3(net20403),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28458_ (.A1(_04377_),
    .A2(_04404_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28459_ (.A1(net17703),
    .A2(net615),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28460_ (.A1(net18089),
    .A2(net17393),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28461_ (.A1(_04338_),
    .A2(_04405_),
    .A3(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28462_ (.A1(_04053_),
    .A2(_04080_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28463_ (.A1(_04408_),
    .A2(net18553),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28464_ (.A1(_04251_),
    .A2(net17696),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28465_ (.A1(_04409_),
    .A2(_04410_),
    .A3(net19645),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28466_ (.A1(_04407_),
    .A2(_04411_),
    .A3(net19626),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28467_ (.A1(_04115_),
    .A2(net18382),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28468_ (.A1(_04338_),
    .A2(_03862_),
    .A3(_04413_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28469_ (.A1(_04295_),
    .A2(net18549),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28470_ (.A1(_16058_[0]),
    .A2(_16067_[0]),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28471_ (.A1(net18536),
    .A2(_04416_),
    .B(net19630),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28472_ (.A1(_04415_),
    .A2(_04417_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28473_ (.A1(_04414_),
    .A2(net19112),
    .A3(_04418_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28474_ (.A1(_04412_),
    .A2(_04419_),
    .A3(net19623),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28475_ (.A1(net17241),
    .A2(net18085),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28476_ (.A1(net17406),
    .A2(net18516),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28477_ (.A1(_04421_),
    .A2(_04422_),
    .A3(net19640),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28478_ (.A1(net18085),
    .A2(_04357_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28479_ (.A1(_04424_),
    .A2(net18536),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28480_ (.A1(_04425_),
    .A2(net19630),
    .A3(_04191_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28481_ (.A1(_04423_),
    .A2(_04426_),
    .A3(net19112),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28482_ (.A1(net17695),
    .A2(_04068_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28483_ (.A1(net18101),
    .A2(net18532),
    .A3(net17400),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28484_ (.A1(_04429_),
    .A2(net19640),
    .A3(_04428_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28485_ (.A1(_04098_),
    .A2(net18549),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28486_ (.A1(net18084),
    .A2(net18099),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28487_ (.A1(_04432_),
    .A2(_04033_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28488_ (.A1(_04430_),
    .A2(_04433_),
    .A3(net19626),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28489_ (.A1(_04427_),
    .A2(net19953),
    .A3(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28490_ (.A1(_04435_),
    .A2(_04420_),
    .A3(net20196),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28491_ (.A1(_04342_),
    .A2(_04068_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28492_ (.A1(_03926_),
    .A2(_04068_),
    .A3(net18554),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28493_ (.A1(_04437_),
    .A2(_04438_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28494_ (.A1(_04439_),
    .A2(net19631),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28495_ (.A1(net18516),
    .A2(_04357_),
    .A3(net18535),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28496_ (.A1(_04441_),
    .A2(_04438_),
    .A3(net19640),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28497_ (.A1(_04440_),
    .A2(_04442_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28498_ (.A1(_04443_),
    .A2(net19116),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28499_ (.A1(_03969_),
    .A2(net19636),
    .A3(_04108_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28500_ (.I(_04233_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28501_ (.A1(_04446_),
    .A2(net18542),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28502_ (.A1(net17398),
    .A2(net19644),
    .A3(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28503_ (.A1(_04445_),
    .A2(_04448_),
    .A3(net19626),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28504_ (.A1(_04449_),
    .A2(net19623),
    .A3(_04444_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28505_ (.A1(_04109_),
    .A2(net17397),
    .B(_04282_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28506_ (.A1(_04451_),
    .A2(net19630),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28507_ (.A1(_04154_),
    .A2(net19640),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28508_ (.A1(_04452_),
    .A2(_04453_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28509_ (.A1(_04454_),
    .A2(net19626),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28510_ (.I(_16059_[0]),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28511_ (.A1(net18554),
    .A2(_04456_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _28512_ (.A1(_04109_),
    .A2(net17399),
    .B(_04457_),
    .C(net19640),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28513_ (.A1(net18086),
    .A2(net18553),
    .A3(net462),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28514_ (.A1(_04459_),
    .A2(_04070_),
    .A3(net19635),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28515_ (.A1(_04458_),
    .A2(_04460_),
    .A3(net19116),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28516_ (.A1(_04455_),
    .A2(_04461_),
    .A3(net19954),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28517_ (.A1(_04450_),
    .A2(net20403),
    .A3(_04462_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28518_ (.A1(_04436_),
    .A2(_04463_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _28519_ (.A1(net18090),
    .A2(net18110),
    .B1(net17407),
    .B2(_04446_),
    .C(net19630),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28520_ (.A1(_04278_),
    .A2(net18534),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28521_ (.A1(net18549),
    .A2(_16067_[0]),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _28522_ (.A1(_04465_),
    .A2(net19640),
    .A3(_04466_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28523_ (.A1(net17395),
    .A2(net18543),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28524_ (.A1(_04467_),
    .A2(_04468_),
    .B(net19119),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28525_ (.A1(_04464_),
    .A2(_04469_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28526_ (.A1(_04324_),
    .A2(_03899_),
    .A3(_04072_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28527_ (.A1(net18094),
    .A2(net18556),
    .B(net19630),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28528_ (.A1(_04472_),
    .A2(_04012_),
    .B(net19624),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28529_ (.A1(_04471_),
    .A2(_04473_),
    .B(net19622),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28530_ (.A1(_04470_),
    .A2(_04474_),
    .B(net20402),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28531_ (.A1(_04431_),
    .A2(_04086_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28532_ (.A1(net19624),
    .A2(_04009_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28533_ (.A1(_04476_),
    .A2(_04477_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28534_ (.A1(net18115),
    .A2(net18545),
    .A3(_04009_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28535_ (.A1(net18087),
    .A2(net18551),
    .A3(net18095),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28536_ (.A1(_04479_),
    .A2(_04480_),
    .B(net19627),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28537_ (.A1(_04478_),
    .A2(_04481_),
    .B(net19641),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28538_ (.A1(net18381),
    .A2(net18548),
    .B(_03946_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28539_ (.A1(_04483_),
    .A2(_04415_),
    .B(net19640),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28540_ (.A1(net18088),
    .A2(net18114),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28541_ (.A1(_04485_),
    .A2(net19113),
    .A3(_04268_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28542_ (.A1(_04484_),
    .A2(_04486_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28543_ (.A1(_04482_),
    .A2(_03993_),
    .A3(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28544_ (.A1(_04475_),
    .A2(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28545_ (.A1(_03902_),
    .A2(net19640),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28546_ (.A1(_04131_),
    .A2(net18557),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28547_ (.A1(_04490_),
    .A2(_04491_),
    .B(net19119),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28548_ (.A1(net18547),
    .A2(_04081_),
    .B(_04022_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28549_ (.A1(_04493_),
    .A2(net19638),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28550_ (.A1(_04492_),
    .A2(_04494_),
    .B(_03993_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28551_ (.A1(net18543),
    .A2(net19124),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28552_ (.A1(_04334_),
    .A2(net19639),
    .A3(_04496_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28553_ (.A1(net18518),
    .A2(net18115),
    .A3(net18543),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28554_ (.A1(_04204_),
    .A2(_04498_),
    .B(net19639),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28555_ (.A1(_04497_),
    .A2(_04499_),
    .B(net19120),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28556_ (.A1(_04495_),
    .A2(_04500_),
    .B(_04062_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28557_ (.A1(_04369_),
    .A2(net18099),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28558_ (.A1(_04197_),
    .A2(_04009_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28559_ (.A1(_04502_),
    .A2(_04503_),
    .A3(net19633),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28560_ (.I(net17394),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28561_ (.A1(_04325_),
    .A2(net19642),
    .A3(_04505_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28562_ (.A1(_04504_),
    .A2(_04506_),
    .A3(_03946_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28563_ (.A1(_04216_),
    .A2(net19647),
    .A3(_04410_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28564_ (.A1(_04112_),
    .A2(net17396),
    .A3(net19637),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28565_ (.A1(_04508_),
    .A2(net19629),
    .A3(_04509_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28566_ (.A1(_04507_),
    .A2(_04510_),
    .A3(_03993_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28567_ (.A1(_04501_),
    .A2(_04511_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28568_ (.A1(_04489_),
    .A2(_04512_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28569_ (.A1(_01588_),
    .A2(_01564_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28570_ (.A1(_01562_),
    .A2(_01560_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28571_ (.A1(_04514_),
    .A2(_04513_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28572_ (.A1(net21368),
    .A2(_10351_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28573_ (.A1(net21099),
    .A2(_10342_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28574_ (.A1(_04516_),
    .A2(_04517_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28575_ (.A1(_04518_),
    .A2(_04515_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28576_ (.A1(_04517_),
    .A2(_04516_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28577_ (.A1(_04514_),
    .A2(_04513_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28578_ (.A1(_04520_),
    .A2(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28579_ (.A1(_04519_),
    .A2(_04522_),
    .A3(_10378_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28580_ (.I(net21226),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28581_ (.A1(_10378_),
    .A2(\text_in_r[97] ),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28582_ (.A1(_04523_),
    .A2(_04524_),
    .A3(_04525_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28583_ (.A1(_04520_),
    .A2(_04515_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28584_ (.A1(_04518_),
    .A2(_04521_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28585_ (.A1(_04527_),
    .A2(_04528_),
    .A3(_10378_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28586_ (.A1(net21501),
    .A2(\text_in_r[97] ),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28587_ (.A1(_04529_),
    .A2(net21226),
    .A3(net20965),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28588_ (.A1(_04526_),
    .A2(_04531_),
    .ZN(_16079_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28589_ (.A1(net21061),
    .A2(net605),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28590_ (.A1(net21098),
    .A2(net21372),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28591_ (.A1(_04533_),
    .A2(_04532_),
    .A3(net20969),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28592_ (.A1(net21300),
    .A2(_10395_),
    .A3(_10396_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28593_ (.A1(_04535_),
    .A2(_04534_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28594_ (.A1(net20921),
    .A2(_04536_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28595_ (.A1(_04534_),
    .A2(_04535_),
    .A3(_10351_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28596_ (.A1(_04538_),
    .A2(_04537_),
    .B(net21501),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28597_ (.I(\text_in_r[96] ),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28598_ (.A1(_04540_),
    .A2(net21501),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28599_ (.A1(net20401),
    .A2(net20929),
    .B(net21236),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28600_ (.A1(_04538_),
    .A2(_04537_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28601_ (.A1(net21079),
    .A2(_04543_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28602_ (.I(net21236),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28603_ (.I(_04541_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28604_ (.A1(net20195),
    .A2(_04545_),
    .A3(net20866),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28605_ (.A1(_04547_),
    .A2(_04542_),
    .ZN(_16082_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28606_ (.A1(net21311),
    .A2(net21367),
    .Z(_04548_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28607_ (.A1(net21311),
    .A2(net21367),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28608_ (.A1(_04548_),
    .A2(_04549_),
    .B(net21476),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28609_ (.A1(net21100),
    .A2(_10417_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28610_ (.A1(net21311),
    .A2(net21367),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28611_ (.A1(_04551_),
    .A2(_10450_),
    .A3(_04552_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28612_ (.A1(_04550_),
    .A2(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _28613_ (.A1(net21479),
    .A2(\sa10_sr[2] ),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28614_ (.I(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28615_ (.A1(_04554_),
    .A2(_04556_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28616_ (.A1(_04550_),
    .A2(_04553_),
    .A3(_04555_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28617_ (.A1(_04557_),
    .A2(_04558_),
    .B(net21501),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28618_ (.I(\text_in_r[98] ),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28619_ (.A1(_04560_),
    .A2(net21504),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28620_ (.I(net21217),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28621_ (.A1(_04559_),
    .A2(_04561_),
    .B(_04562_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28622_ (.A1(_04557_),
    .A2(_04558_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28623_ (.A1(_04564_),
    .A2(net21070),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28624_ (.I(_04561_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28625_ (.A1(_04565_),
    .A2(net21217),
    .A3(_04566_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28626_ (.A1(_04563_),
    .A2(_04567_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input170 (.I(text_in[1]),
    .Z(net170));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28628_ (.A1(_04541_),
    .A2(_04539_),
    .B(_04545_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28629_ (.A1(_04546_),
    .A2(net21236),
    .A3(_04544_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28630_ (.A1(_04570_),
    .A2(_04569_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input169 (.I(text_in[19]),
    .Z(net169));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28632_ (.A1(_04559_),
    .A2(_04561_),
    .B(net21217),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28633_ (.A1(_04565_),
    .A2(_04562_),
    .A3(_04566_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28634_ (.A1(_04572_),
    .A2(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input168 (.I(text_in[18]),
    .Z(net168));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input167 (.I(text_in[17]),
    .Z(net167));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28637_ (.A1(net19616),
    .A2(net19610),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28638_ (.A1(_10453_),
    .A2(net21365),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28639_ (.A1(_10457_),
    .A2(net21053),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28640_ (.A1(_04577_),
    .A2(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28641_ (.A1(_01634_),
    .A2(net20629),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28642_ (.I(_04579_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28643_ (.A1(net20423),
    .A2(_04581_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28644_ (.A1(_04580_),
    .A2(_04582_),
    .A3(net21075),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28645_ (.I(net21214),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _28646_ (.A1(net21077),
    .A2(\text_in_r[99] ),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28647_ (.A1(_04583_),
    .A2(_04584_),
    .A3(_04585_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28648_ (.A1(_01634_),
    .A2(_04581_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28649_ (.A1(net20423),
    .A2(net20629),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28650_ (.A1(_04587_),
    .A2(_04588_),
    .A3(net21075),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28651_ (.A1(net21501),
    .A2(\text_in_r[99] ),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28652_ (.A1(_04589_),
    .A2(net21214),
    .A3(_04590_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28653_ (.A1(_04586_),
    .A2(_04591_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28654_ (.A1(_04576_),
    .A2(net19097),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28655_ (.A1(_04525_),
    .A2(net21226),
    .A3(_04523_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28656_ (.A1(_04529_),
    .A2(_04524_),
    .A3(_04530_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28657_ (.A1(_04594_),
    .A2(_04595_),
    .ZN(_16074_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _28658_ (.A1(net19610),
    .A2(net19602),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28659_ (.A1(_04596_),
    .A2(net19606),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28660_ (.A1(_04593_),
    .A2(_04597_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28661_ (.A1(net19602),
    .A2(net19614),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input166 (.I(text_in[16]),
    .Z(net166));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28663_ (.A1(net18953),
    .A2(net19606),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28664_ (.A1(_04599_),
    .A2(_04601_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28665_ (.A1(_04589_),
    .A2(_04584_),
    .A3(_04590_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28666_ (.A1(_04583_),
    .A2(net21214),
    .A3(_04585_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28667_ (.A1(_04603_),
    .A2(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input165 (.I(net592),
    .Z(net165));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input164 (.I(text_in[14]),
    .Z(net164));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28670_ (.A1(_04602_),
    .A2(net19088),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28671_ (.A1(_04598_),
    .A2(_04608_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28672_ (.A1(net20912),
    .A2(net20804),
    .B(net21078),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28673_ (.A1(net20912),
    .A2(_01654_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28674_ (.I(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28675_ (.A1(net21501),
    .A2(\text_in_r[100] ),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28676_ (.A1(_04610_),
    .A2(_04612_),
    .B(_04613_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28677_ (.I(net21213),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28678_ (.A1(_04614_),
    .A2(_04615_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28679_ (.A1(net20912),
    .A2(_01654_),
    .Z(_04617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28680_ (.A1(_04617_),
    .A2(net21078),
    .A3(_04611_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28681_ (.A1(_04618_),
    .A2(net21213),
    .A3(_04613_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28682_ (.A1(_04616_),
    .A2(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input163 (.I(net600),
    .Z(net163));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28684_ (.A1(_04609_),
    .A2(net19588),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input162 (.I(text_in[12]),
    .Z(net162));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input161 (.I(text_in[127]),
    .Z(net161));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _28687_ (.I(_16089_[0]),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28688_ (.A1(net20194),
    .A2(_04625_),
    .A3(net19952),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28689_ (.A1(net19111),
    .A2(net19107),
    .A3(_04626_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input160 (.I(text_in[126]),
    .Z(net160));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28691_ (.A1(_04627_),
    .A2(net19588),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28692_ (.A1(net19619),
    .A2(net19612),
    .A3(net19608),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28693_ (.I(_04630_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28694_ (.A1(net19602),
    .A2(net19606),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input159 (.I(text_in[125]),
    .Z(net159));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28696_ (.A1(_04632_),
    .A2(net19082),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28697_ (.A1(_04631_),
    .A2(_04634_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _28698_ (.A1(net21302),
    .A2(\sa20_sr[5] ),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28699_ (.A1(_04636_),
    .A2(net21472),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28700_ (.A1(_04636_),
    .A2(net21472),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28701_ (.A1(_04637_),
    .A2(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28702_ (.A1(net21473),
    .A2(\sa10_sr[5] ),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28703_ (.A1(_04639_),
    .A2(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28704_ (.I(_04640_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28705_ (.A1(_04637_),
    .A2(_04642_),
    .A3(_04638_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28706_ (.A1(_04641_),
    .A2(_04643_),
    .A3(net21065),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28707_ (.A1(net21494),
    .A2(\text_in_r[101] ),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28708_ (.A1(_04644_),
    .A2(_04645_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28709_ (.I(net21212),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28710_ (.A1(_04646_),
    .A2(_04647_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28711_ (.A1(_04644_),
    .A2(net21212),
    .A3(_04645_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28712_ (.A1(_04648_),
    .A2(_04649_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _28713_ (.I(_04650_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input158 (.I(text_in[124]),
    .Z(net158));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28715_ (.A1(_04629_),
    .A2(_04635_),
    .B(_04651_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28716_ (.A1(_04622_),
    .A2(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28717_ (.A1(net19606),
    .A2(net19610),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28718_ (.A1(_04655_),
    .A2(net19082),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28719_ (.A1(_04656_),
    .A2(_04630_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28720_ (.A1(_04657_),
    .A2(net19593),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28721_ (.I(_16076_[0]),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28722_ (.A1(_04574_),
    .A2(_04659_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28723_ (.A1(_04660_),
    .A2(net19097),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _28724_ (.I(_04661_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28725_ (.A1(net19612),
    .A2(_04625_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28726_ (.A1(_04662_),
    .A2(_04663_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28727_ (.A1(_04664_),
    .A2(_04658_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28728_ (.I(_16080_[0]),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28729_ (.A1(net18506),
    .A2(net19606),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input157 (.I(text_in[123]),
    .Z(net157));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28731_ (.A1(_04667_),
    .A2(net19103),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28732_ (.A1(_04631_),
    .A2(_04669_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28733_ (.A1(_04576_),
    .A2(net19082),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28734_ (.A1(_04614_),
    .A2(net21213),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28735_ (.A1(_04618_),
    .A2(_04615_),
    .A3(_04613_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28736_ (.A1(_04672_),
    .A2(_04673_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input156 (.I(text_in[122]),
    .Z(net156));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28738_ (.A1(net18505),
    .A2(net19581),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input155 (.I(text_in[121]),
    .Z(net155));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input154 (.I(text_in[120]),
    .Z(net154));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28741_ (.A1(_04670_),
    .A2(_04676_),
    .B(net19945),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28742_ (.A1(_04679_),
    .A2(_04665_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28743_ (.A1(\sa30_sr[5] ),
    .A2(\sa20_sr[6] ),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28744_ (.A1(\sa00_sr[6] ),
    .A2(_04681_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28745_ (.A1(net21472),
    .A2(net21416),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28746_ (.A1(_04682_),
    .A2(_04683_),
    .Z(_04684_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28747_ (.A1(_04682_),
    .A2(_04683_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28748_ (.A1(net21494),
    .A2(\text_in_r[102] ),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _28749_ (.A1(_04684_),
    .A2(net21494),
    .A3(_04685_),
    .B(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28750_ (.A1(_04687_),
    .A2(\u0.w[0][6] ),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28751_ (.A1(_04687_),
    .A2(\u0.w[0][6] ),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28752_ (.A1(_04688_),
    .A2(_04689_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _28753_ (.I(_04690_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input153 (.I(net567),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28755_ (.A1(_04680_),
    .A2(_04654_),
    .B(net20192),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28756_ (.I(_16075_[0]),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28757_ (.A1(net19614),
    .A2(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28758_ (.I(_16083_[0]),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28759_ (.A1(net19606),
    .A2(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28760_ (.A1(_04695_),
    .A2(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28761_ (.A1(_04698_),
    .A2(net19109),
    .B(net19588),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28762_ (.A1(net19614),
    .A2(_04596_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28763_ (.A1(_04660_),
    .A2(net19082),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28764_ (.A1(_04700_),
    .A2(_04701_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28765_ (.A1(_04699_),
    .A2(_04702_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28766_ (.A1(net19602),
    .A2(net511),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28767_ (.A1(net19603),
    .A2(net19617),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28768_ (.A1(_04704_),
    .A2(net19072),
    .A3(net19090),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28769_ (.A1(net19619),
    .A2(net19608),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28770_ (.A1(net19616),
    .A2(net19617),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28771_ (.A1(_04707_),
    .A2(_04708_),
    .A3(net19097),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28772_ (.A1(_04706_),
    .A2(_04709_),
    .A3(net19599),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28773_ (.A1(_04703_),
    .A2(_04710_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input152 (.I(text_in[119]),
    .Z(net152));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28775_ (.A1(_04711_),
    .A2(net19950),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28776_ (.A1(net19615),
    .A2(net18955),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28777_ (.A1(net18080),
    .A2(_04714_),
    .A3(net19107),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28778_ (.A1(net19606),
    .A2(net18955),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28779_ (.A1(net19611),
    .A2(_16083_[0]),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28780_ (.A1(_04716_),
    .A2(net18497),
    .A3(net19083),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28781_ (.A1(_04715_),
    .A2(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input151 (.I(text_in[118]),
    .Z(net151));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28783_ (.A1(_04719_),
    .A2(net19579),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input150 (.I(net601),
    .Z(net150));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28785_ (.A1(net19618),
    .A2(net19611),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28786_ (.A1(net18954),
    .A2(net19606),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input149 (.I(text_in[116]),
    .Z(net149));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28788_ (.A1(net19066),
    .A2(net493),
    .A3(net19082),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input148 (.I(text_in[115]),
    .Z(net148));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28790_ (.A1(net19613),
    .A2(_04659_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28791_ (.A1(_04728_),
    .A2(net19097),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28792_ (.A1(_04726_),
    .A2(net19588),
    .A3(net17688),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28793_ (.A1(_04721_),
    .A2(_04651_),
    .A3(_04730_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input147 (.I(text_in[114]),
    .Z(net147));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28795_ (.A1(_04713_),
    .A2(_04731_),
    .A3(net20400),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28796_ (.A1(_04733_),
    .A2(_04693_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28797_ (.A1(\sa30_sr[6] ),
    .A2(net20915),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _28798_ (.A1(_13742_),
    .A2(net21362),
    .A3(_04735_),
    .Z(_04736_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28799_ (.A1(net21493),
    .A2(\text_in_r[103] ),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28800_ (.A1(_04736_),
    .A2(net21065),
    .B(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _28801_ (.A1(\u0.w[0][7] ),
    .A2(_04738_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input146 (.I(net574),
    .Z(net146));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28803_ (.A1(net20190),
    .A2(_04734_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28804_ (.A1(net19615),
    .A2(net18952),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28805_ (.A1(_04742_),
    .A2(net19103),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28806_ (.A1(_04743_),
    .A2(net19581),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28807_ (.A1(_04744_),
    .A2(_04598_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28808_ (.A1(net19606),
    .A2(_16085_[0]),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28809_ (.A1(_04742_),
    .A2(_04746_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28810_ (.A1(_04747_),
    .A2(net19088),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28811_ (.A1(_04748_),
    .A2(net19588),
    .A3(net17689),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input145 (.I(net543),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28813_ (.A1(_04745_),
    .A2(_04749_),
    .A3(net19586),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28814_ (.A1(net19619),
    .A2(net19603),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28815_ (.A1(net18954),
    .A2(net19614),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28816_ (.A1(_04752_),
    .A2(_04753_),
    .A3(net19094),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28817_ (.A1(_04754_),
    .A2(net19571),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28818_ (.A1(net19075),
    .A2(net18497),
    .A3(net19098),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _28819_ (.A1(_04755_),
    .A2(_04756_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input144 (.I(text_in[111]),
    .Z(net144));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28821_ (.A1(_04669_),
    .A2(net19588),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28822_ (.A1(_04695_),
    .A2(_04601_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input143 (.I(text_in[110]),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28824_ (.A1(_04760_),
    .A2(net19088),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28825_ (.A1(_04759_),
    .A2(_04762_),
    .B(_04651_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28826_ (.A1(_04757_),
    .A2(_04763_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28827_ (.A1(_04751_),
    .A2(_04764_),
    .B(net20400),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28828_ (.I(_16085_[0]),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28829_ (.A1(_04766_),
    .A2(net19612),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28830_ (.A1(_04767_),
    .A2(net19097),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28831_ (.A1(net19619),
    .A2(net19604),
    .A3(net19608),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28832_ (.A1(_04768_),
    .A2(net19062),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28833_ (.I(_04601_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28834_ (.A1(net18070),
    .A2(net19093),
    .B(net19588),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28835_ (.A1(_04770_),
    .A2(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28836_ (.A1(_04717_),
    .A2(net19082),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28837_ (.I(_04774_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28838_ (.A1(net17685),
    .A2(net19062),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28839_ (.A1(_04771_),
    .A2(net19098),
    .B(net19571),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28840_ (.A1(_04776_),
    .A2(net17684),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input142 (.I(net598),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28842_ (.A1(_04773_),
    .A2(_04778_),
    .A3(net19945),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28843_ (.A1(net19614),
    .A2(net18506),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28844_ (.A1(_04769_),
    .A2(net19094),
    .A3(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28845_ (.A1(_04593_),
    .A2(_04716_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28846_ (.A1(net19614),
    .A2(net18953),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28847_ (.I(_04784_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28848_ (.A1(_04785_),
    .A2(net19087),
    .B(net19588),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28849_ (.A1(net17683),
    .A2(_04783_),
    .A3(_04786_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28850_ (.A1(net19082),
    .A2(_16096_[0]),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28851_ (.A1(_04753_),
    .A2(net19082),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28852_ (.A1(_04788_),
    .A2(net18062),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28853_ (.A1(_04790_),
    .A2(net19588),
    .B(net19945),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28854_ (.A1(_04787_),
    .A2(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28855_ (.A1(_04780_),
    .A2(_04792_),
    .B(net20192),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _28856_ (.I(_04739_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28857_ (.A1(_04765_),
    .A2(_04793_),
    .B(_04794_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28858_ (.A1(_04795_),
    .A2(_04741_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28859_ (.A1(_04708_),
    .A2(net19089),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28860_ (.A1(net19606),
    .A2(_04694_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28861_ (.A1(_04796_),
    .A2(_04797_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28862_ (.A1(_04662_),
    .A2(net18494),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28863_ (.A1(_04798_),
    .A2(_04799_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input141 (.I(text_in[109]),
    .Z(net141));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28865_ (.A1(_04800_),
    .A2(net19597),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _28866_ (.I(_04789_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28867_ (.A1(_04803_),
    .A2(net19076),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28868_ (.A1(net19619),
    .A2(net19617),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28869_ (.A1(_04805_),
    .A2(net19075),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input140 (.I(text_in[108]),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28871_ (.A1(_04806_),
    .A2(net19110),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input139 (.I(text_in[107]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28873_ (.A1(_04804_),
    .A2(_04808_),
    .A3(net19571),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28874_ (.A1(_04802_),
    .A2(_04810_),
    .A3(_04651_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input138 (.I(text_in[106]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28876_ (.A1(net513),
    .A2(net19101),
    .A3(net18495),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28877_ (.A1(net19086),
    .A2(net18952),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28878_ (.A1(_04814_),
    .A2(net19607),
    .B(net19588),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28879_ (.A1(_04813_),
    .A2(_04815_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28880_ (.A1(_04632_),
    .A2(_04663_),
    .A3(net19108),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28881_ (.A1(_04805_),
    .A2(net19606),
    .A3(net19091),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input137 (.I(text_in[105]),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28883_ (.A1(_04817_),
    .A2(_04818_),
    .A3(net19598),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28884_ (.A1(_04816_),
    .A2(_04820_),
    .A3(net19950),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28885_ (.A1(_04811_),
    .A2(_04821_),
    .A3(net20193),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28886_ (.A1(_04752_),
    .A2(net19082),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28887_ (.A1(_04823_),
    .A2(net19073),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28888_ (.A1(net19097),
    .A2(net19611),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28889_ (.A1(_04825_),
    .A2(_04707_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28890_ (.A1(_04824_),
    .A2(net19580),
    .A3(net18061),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28891_ (.A1(net18510),
    .A2(net523),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28892_ (.A1(net19068),
    .A2(_04667_),
    .A3(net19087),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28893_ (.A1(_04828_),
    .A2(net19595),
    .A3(_04829_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28894_ (.A1(_04827_),
    .A2(_04830_),
    .A3(net19945),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28895_ (.A1(_04743_),
    .A2(net19588),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28896_ (.A1(_04723_),
    .A2(net19097),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28897_ (.A1(net18491),
    .A2(net19079),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28898_ (.A1(_04832_),
    .A2(_04834_),
    .B(net19945),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _28899_ (.I(_04729_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28900_ (.A1(_04836_),
    .A2(net18082),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28901_ (.A1(net17683),
    .A2(_04837_),
    .A3(net19573),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28902_ (.A1(_04835_),
    .A2(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28903_ (.A1(_04831_),
    .A2(_04839_),
    .A3(net20400),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28904_ (.A1(_04822_),
    .A2(_04840_),
    .A3(_04794_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28905_ (.A1(net19068),
    .A2(_04601_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input136 (.I(text_in[104]),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28907_ (.A1(_04842_),
    .A2(net19086),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28908_ (.A1(_04716_),
    .A2(net18075),
    .A3(net19098),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28909_ (.A1(_04844_),
    .A2(_04845_),
    .A3(net19595),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _28910_ (.A1(net19095),
    .A2(_04667_),
    .A3(net19107),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28911_ (.A1(net19071),
    .A2(net18499),
    .A3(net19083),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input135 (.I(text_in[103]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28913_ (.A1(_04847_),
    .A2(_04848_),
    .A3(net19580),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28914_ (.A1(_04846_),
    .A2(_04850_),
    .A3(net19951),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28915_ (.I(_04671_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28916_ (.A1(net18059),
    .A2(_04597_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28917_ (.A1(_04661_),
    .A2(net19571),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28918_ (.A1(_04853_),
    .A2(_04854_),
    .B(net19950),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28919_ (.A1(_04626_),
    .A2(net19082),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _28920_ (.I(_16077_[0]),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28921_ (.A1(net19614),
    .A2(net18490),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28922_ (.A1(_04856_),
    .A2(net18058),
    .B(net19574),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28923_ (.A1(_04813_),
    .A2(_04859_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28924_ (.A1(_04855_),
    .A2(_04860_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28925_ (.A1(_04851_),
    .A2(_04861_),
    .B(net20400),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28926_ (.A1(net19097),
    .A2(net19606),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28927_ (.A1(_04863_),
    .A2(net19608),
    .B(_04651_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28928_ (.A1(_04707_),
    .A2(_04752_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28929_ (.A1(_04865_),
    .A2(net19098),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28930_ (.A1(_04656_),
    .A2(_04714_),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28931_ (.A1(_04864_),
    .A2(_04866_),
    .A3(_04867_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28932_ (.A1(_04705_),
    .A2(net19082),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28933_ (.I(_04869_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28934_ (.A1(_04870_),
    .A2(net19067),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28935_ (.A1(_04871_),
    .A2(_04651_),
    .A3(_04847_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28936_ (.A1(_04868_),
    .A2(_04872_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _28937_ (.A1(_04650_),
    .A2(_16099_[0]),
    .A3(net19093),
    .Z(_04874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28938_ (.A1(_04597_),
    .A2(_04775_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28939_ (.A1(_04874_),
    .A2(_04875_),
    .A3(net19571),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input134 (.I(text_in[102]),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28941_ (.A1(_04876_),
    .A2(net20400),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28942_ (.A1(_04873_),
    .A2(net19588),
    .B(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28943_ (.A1(_04862_),
    .A2(_04879_),
    .B(net20190),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28944_ (.A1(_04841_),
    .A2(_04880_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28945_ (.A1(_04781_),
    .A2(net19106),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28946_ (.A1(_04881_),
    .A2(net19078),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28947_ (.A1(_04882_),
    .A2(net19577),
    .A3(_04748_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28948_ (.A1(_04746_),
    .A2(net19097),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28949_ (.A1(_04884_),
    .A2(net19578),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28950_ (.A1(net19077),
    .A2(net18065),
    .A3(net19106),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28951_ (.A1(net19612),
    .A2(net18951),
    .Z(_04887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28952_ (.A1(_04887_),
    .A2(net19082),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28953_ (.A1(_04885_),
    .A2(_04886_),
    .A3(_04888_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28954_ (.A1(_04883_),
    .A2(_04889_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28955_ (.A1(_04890_),
    .A2(net19583),
    .B(net20400),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28956_ (.A1(_04656_),
    .A2(net18071),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28957_ (.A1(net652),
    .A2(net18493),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _28958_ (.A1(_04892_),
    .A2(_04893_),
    .A3(net19950),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28959_ (.A1(net19945),
    .A2(net19588),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28960_ (.A1(_04599_),
    .A2(net19097),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28961_ (.A1(_04896_),
    .A2(_04746_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28962_ (.A1(_04869_),
    .A2(_04887_),
    .B(net19588),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28963_ (.A1(_04897_),
    .A2(_04898_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28964_ (.A1(_04894_),
    .A2(_04895_),
    .B(_04899_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _28965_ (.A1(_04900_),
    .A2(_04891_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28966_ (.A1(_04724_),
    .A2(net19082),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28967_ (.A1(_04902_),
    .A2(net19095),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28968_ (.A1(net19071),
    .A2(_04784_),
    .A3(net19107),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28969_ (.A1(_04903_),
    .A2(_04904_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28970_ (.A1(_04905_),
    .A2(net19577),
    .B(net19950),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input133 (.I(text_in[101]),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28972_ (.A1(net18503),
    .A2(net19106),
    .A3(net18082),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28973_ (.A1(_04630_),
    .A2(net19092),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28974_ (.A1(_04908_),
    .A2(net18487),
    .B(net19588),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28975_ (.A1(_04906_),
    .A2(_04910_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28976_ (.A1(_04865_),
    .A2(net19591),
    .A3(net19099),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28977_ (.A1(net19588),
    .A2(_04663_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _28978_ (.A1(_04667_),
    .A2(net19082),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28979_ (.A1(_04913_),
    .A2(_04914_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28980_ (.A1(_04915_),
    .A2(net19945),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28981_ (.A1(_04912_),
    .A2(_04916_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28982_ (.A1(_04769_),
    .A2(net18067),
    .B(net19094),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28983_ (.A1(_04755_),
    .A2(_04918_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28984_ (.A1(_04917_),
    .A2(_04919_),
    .B(net20400),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _28985_ (.A1(_04911_),
    .A2(_04920_),
    .B(net20187),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _28986_ (.A1(_04921_),
    .A2(_04901_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28987_ (.A1(_16103_[0]),
    .A2(net19093),
    .B(net19945),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28988_ (.A1(_04866_),
    .A2(_04923_),
    .B(net19576),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _28989_ (.A1(_04666_),
    .A2(_04857_),
    .Z(_04925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _28990_ (.I(net18056),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28991_ (.A1(_04863_),
    .A2(_04926_),
    .B(_04651_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28992_ (.A1(net19095),
    .A2(net19111),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28993_ (.A1(_04928_),
    .A2(net19107),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _28994_ (.A1(_04927_),
    .A2(_04875_),
    .A3(_04929_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28995_ (.A1(_04924_),
    .A2(_04930_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28996_ (.A1(net19091),
    .A2(_04797_),
    .B(_04651_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _28997_ (.A1(net652),
    .A2(net18064),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _28998_ (.A1(_04932_),
    .A2(_04933_),
    .B(net19588),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _28999_ (.A1(net19082),
    .A2(_16094_[0]),
    .Z(_04935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29000_ (.A1(_04909_),
    .A2(_04935_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29001_ (.A1(_04936_),
    .A2(net19950),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29002_ (.A1(_04934_),
    .A2(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29003_ (.A1(_04931_),
    .A2(_04938_),
    .A3(net20400),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29004_ (.A1(_04896_),
    .A2(net19075),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29005_ (.A1(_04940_),
    .A2(net19590),
    .A3(net18072),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29006_ (.A1(_04836_),
    .A2(net19063),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29007_ (.A1(net18950),
    .A2(net19092),
    .B(net19588),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29008_ (.A1(_04942_),
    .A2(_04943_),
    .B(net19584),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29009_ (.A1(_04941_),
    .A2(_04944_),
    .B(net20400),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29010_ (.A1(_04823_),
    .A2(_04695_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29011_ (.A1(net18493),
    .A2(net18077),
    .A3(net19109),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29012_ (.A1(_04946_),
    .A2(_04947_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29013_ (.A1(_04948_),
    .A2(net19588),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29014_ (.A1(net19074),
    .A2(_04752_),
    .A3(net19098),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29015_ (.A1(net19107),
    .A2(_16099_[0]),
    .Z(_04951_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29016_ (.A1(_04950_),
    .A2(net19579),
    .A3(_04951_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29017_ (.A1(_04949_),
    .A2(_04952_),
    .A3(_04651_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29018_ (.A1(_04945_),
    .A2(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29019_ (.A1(_04939_),
    .A2(_04954_),
    .B(net20187),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29020_ (.A1(_04922_),
    .A2(_04955_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29021_ (.A1(_04881_),
    .A2(net18082),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29022_ (.A1(net19950),
    .A2(net19571),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29023_ (.A1(_04903_),
    .A2(_04956_),
    .A3(_04957_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29024_ (.A1(_04958_),
    .A2(net20400),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29025_ (.I(_04797_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29026_ (.A1(_04836_),
    .A2(_04960_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29027_ (.A1(_04708_),
    .A2(net19091),
    .A3(_04697_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29028_ (.A1(_04961_),
    .A2(_04962_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29029_ (.A1(_04963_),
    .A2(_04895_),
    .Z(_04964_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29030_ (.A1(_04959_),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29031_ (.A1(_04704_),
    .A2(_04708_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29032_ (.A1(_04966_),
    .A2(net19091),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29033_ (.A1(net19095),
    .A2(net514),
    .A3(net19109),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29034_ (.A1(_04967_),
    .A2(_04968_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29035_ (.A1(_04969_),
    .A2(net19579),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29036_ (.I(net18074),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29037_ (.A1(_04971_),
    .A2(net19098),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29038_ (.I(_04972_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29039_ (.A1(_04871_),
    .A2(_04973_),
    .A3(net19589),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29040_ (.A1(_04970_),
    .A2(_04974_),
    .A3(net19583),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29041_ (.A1(_04965_),
    .A2(_04975_),
    .B(net20188),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _29042_ (.A1(net19095),
    .A2(_04708_),
    .A3(_04697_),
    .A4(net19109),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29043_ (.A1(_04805_),
    .A2(net19607),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29044_ (.A1(_04803_),
    .A2(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29045_ (.A1(_04979_),
    .A2(net19579),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29046_ (.A1(net19615),
    .A2(_04696_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29047_ (.I(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29048_ (.A1(_04701_),
    .A2(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29049_ (.A1(_04983_),
    .A2(net19599),
    .A3(_04709_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29050_ (.A1(_04977_),
    .A2(_04980_),
    .B(_04984_),
    .C(net19950),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29051_ (.A1(_04902_),
    .A2(net18071),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29052_ (.A1(_04986_),
    .A2(net19598),
    .A3(_04817_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _29053_ (.A1(_04966_),
    .A2(net19588),
    .A3(_04863_),
    .Z(_04988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29054_ (.A1(_04987_),
    .A2(_04988_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29055_ (.A1(_04989_),
    .A2(net19587),
    .B(net20400),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29056_ (.A1(_04985_),
    .A2(_04990_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29057_ (.A1(_04976_),
    .A2(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29058_ (.A1(_04925_),
    .A2(net19606),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29059_ (.A1(net19097),
    .A2(_04993_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29060_ (.A1(_04994_),
    .A2(net18071),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29061_ (.A1(_04875_),
    .A2(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29062_ (.A1(_04996_),
    .A2(net19576),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29063_ (.A1(_04898_),
    .A2(_04651_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29064_ (.A1(_04997_),
    .A2(_04998_),
    .B(net20400),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29065_ (.A1(_04824_),
    .A2(_04783_),
    .A3(net19580),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29066_ (.A1(net653),
    .A2(net18079),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29067_ (.I(_04746_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29068_ (.A1(_05002_),
    .A2(net19097),
    .B(net19571),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29069_ (.A1(_04825_),
    .A2(net19608),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29070_ (.A1(_05001_),
    .A2(_05003_),
    .A3(_05004_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29071_ (.A1(_05005_),
    .A2(_05000_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29072_ (.A1(_05006_),
    .A2(net19946),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29073_ (.A1(_05007_),
    .A2(_04999_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29074_ (.A1(_04852_),
    .A2(net18080),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29075_ (.A1(net508),
    .A2(_04663_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29076_ (.A1(_05009_),
    .A2(_05010_),
    .A3(_04651_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29077_ (.A1(_05002_),
    .A2(net19097),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29078_ (.A1(_04892_),
    .A2(net19950),
    .A3(_05012_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29079_ (.A1(_05011_),
    .A2(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29080_ (.A1(_05014_),
    .A2(net19572),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29081_ (.I(net19064),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29082_ (.A1(net18069),
    .A2(_05016_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29083_ (.A1(_05017_),
    .A2(_04972_),
    .B(net19582),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29084_ (.I(_04777_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _29085_ (.A1(net18080),
    .A2(net19105),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29086_ (.A1(_05020_),
    .A2(_04651_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29087_ (.A1(_05019_),
    .A2(_05021_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29088_ (.A1(_05018_),
    .A2(_05022_),
    .B(_04691_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29089_ (.A1(_05015_),
    .A2(_05023_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29090_ (.A1(_05008_),
    .A2(_05024_),
    .A3(net20189),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29091_ (.A1(_04992_),
    .A2(_05025_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29092_ (.A1(_04871_),
    .A2(_04950_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29093_ (.A1(_05026_),
    .A2(net19572),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29094_ (.A1(_04599_),
    .A2(_04707_),
    .A3(net19085),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29095_ (.A1(_04752_),
    .A2(_04695_),
    .A3(net19098),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29096_ (.A1(_05028_),
    .A2(_05029_),
    .A3(net19595),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29097_ (.A1(_05027_),
    .A2(_04691_),
    .A3(_05030_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29098_ (.A1(_04769_),
    .A2(net19588),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29099_ (.A1(net19571),
    .A2(_04716_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29100_ (.A1(_05032_),
    .A2(_05033_),
    .B(net18488),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29101_ (.A1(_04782_),
    .A2(net19588),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29102_ (.A1(_04915_),
    .A2(_04691_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29103_ (.A1(_05034_),
    .A2(_05035_),
    .A3(_05036_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29104_ (.A1(_05031_),
    .A2(_05037_),
    .B(_04651_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29105_ (.A1(net17686),
    .A2(net19575),
    .A3(net18070),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29106_ (.A1(_05039_),
    .A2(net20400),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29107_ (.I(_04833_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29108_ (.A1(_05041_),
    .A2(net19075),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29109_ (.A1(_05042_),
    .A2(_04867_),
    .A3(net19572),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29110_ (.A1(_05040_),
    .A2(_05043_),
    .B(_04651_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29111_ (.A1(_04856_),
    .A2(net18076),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29112_ (.A1(_04770_),
    .A2(_05045_),
    .A3(net19572),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _29113_ (.I(_04753_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29114_ (.A1(_05047_),
    .A2(net19100),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29115_ (.A1(net17680),
    .A2(_04748_),
    .A3(net17678),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29116_ (.A1(_05046_),
    .A2(_05049_),
    .A3(net20400),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29117_ (.A1(_05044_),
    .A2(_05050_),
    .B(net20190),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29118_ (.A1(_05038_),
    .A2(_05051_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29119_ (.I(_16087_[0]),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29120_ (.A1(_05053_),
    .A2(net19101),
    .B(_05048_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29121_ (.A1(_05054_),
    .A2(net19947),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29122_ (.A1(_04762_),
    .A2(net18500),
    .A3(_04651_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29123_ (.A1(_05055_),
    .A2(net19573),
    .A3(_05056_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29124_ (.A1(net17687),
    .A2(net19071),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29125_ (.A1(_05058_),
    .A2(_05028_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29126_ (.A1(_04651_),
    .A2(net19588),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29127_ (.A1(_05059_),
    .A2(net19061),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29128_ (.A1(_04768_),
    .A2(net19079),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29129_ (.A1(_04707_),
    .A2(net19605),
    .A3(net19082),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29130_ (.A1(_05062_),
    .A2(_05063_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29131_ (.A1(_05064_),
    .A2(_04895_),
    .B(_04691_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29132_ (.A1(_05057_),
    .A2(_05061_),
    .A3(_05065_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29133_ (.A1(net18502),
    .A2(net19101),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29134_ (.A1(_04858_),
    .A2(net19082),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29135_ (.A1(_05068_),
    .A2(net19588),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29136_ (.A1(_05067_),
    .A2(_05069_),
    .B(_04651_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29137_ (.A1(_04914_),
    .A2(_05047_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29138_ (.A1(net18083),
    .A2(_05071_),
    .A3(net19573),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29139_ (.A1(_05070_),
    .A2(_05072_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29140_ (.A1(_04870_),
    .A2(_04663_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29141_ (.A1(_04825_),
    .A2(net19589),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29142_ (.A1(_05074_),
    .A2(_05075_),
    .B(net19945),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29143_ (.A1(net19067),
    .A2(net19093),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29144_ (.A1(_05077_),
    .A2(net18498),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29145_ (.A1(_05078_),
    .A2(net19591),
    .A3(_04847_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29146_ (.A1(_05076_),
    .A2(_05079_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29147_ (.A1(_05073_),
    .A2(_05080_),
    .A3(_04691_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29148_ (.A1(_05066_),
    .A2(_05081_),
    .A3(net20190),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29149_ (.A1(_05052_),
    .A2(_05082_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29150_ (.A1(_04826_),
    .A2(net19588),
    .A3(_04914_),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29151_ (.A1(net19111),
    .A2(_04746_),
    .B(net19090),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _29152_ (.A1(_05084_),
    .A2(net19588),
    .A3(_04701_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _29153_ (.A1(_05085_),
    .A2(_05083_),
    .A3(net20400),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29154_ (.A1(_05048_),
    .A2(net19588),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29155_ (.I(_05068_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29156_ (.A1(_05088_),
    .A2(net19065),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29157_ (.A1(_05089_),
    .A2(_05087_),
    .B(_04691_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29158_ (.A1(net18080),
    .A2(_04695_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29159_ (.A1(net19082),
    .A2(_05091_),
    .B(_04888_),
    .C(net19571),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29160_ (.A1(_05092_),
    .A2(_05090_),
    .B(net19946),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _29161_ (.A1(_05093_),
    .A2(_05086_),
    .B(net20189),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29162_ (.A1(net18509),
    .A2(net18497),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29163_ (.A1(net18505),
    .A2(net19096),
    .B(net19600),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29164_ (.A1(_05095_),
    .A2(net19109),
    .B(_05096_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29165_ (.A1(net19109),
    .A2(net19602),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29166_ (.A1(_05028_),
    .A2(net19579),
    .A3(_05098_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29167_ (.A1(_05099_),
    .A2(net20400),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29168_ (.A1(_05097_),
    .A2(_05100_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29169_ (.A1(net19063),
    .A2(net19084),
    .A3(net18071),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29170_ (.A1(_04881_),
    .A2(_04926_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29171_ (.A1(_05102_),
    .A2(_05103_),
    .A3(net19595),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29172_ (.I(_04663_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29173_ (.A1(_04669_),
    .A2(_05105_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29174_ (.A1(_05106_),
    .A2(net17690),
    .A3(net19581),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29175_ (.A1(_05104_),
    .A2(_05107_),
    .B(net20400),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29176_ (.A1(_05101_),
    .A2(_05108_),
    .B(net19950),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29177_ (.A1(_05094_),
    .A2(_05109_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29178_ (.A1(_04724_),
    .A2(_04663_),
    .Z(_05111_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29179_ (.A1(_05111_),
    .A2(net19089),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29180_ (.A1(_04662_),
    .A2(net18497),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29181_ (.A1(_05113_),
    .A2(_05112_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29182_ (.A1(_05114_),
    .A2(_05060_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29183_ (.A1(net20400),
    .A2(_05115_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29184_ (.A1(_04597_),
    .A2(net19089),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29185_ (.A1(net19110),
    .A2(net18504),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _29186_ (.A1(_05117_),
    .A2(_05118_),
    .B(net19950),
    .C(net19597),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29187_ (.A1(_05119_),
    .A2(_05116_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29188_ (.I(_04994_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29189_ (.A1(_05117_),
    .A2(net18508),
    .B(net19581),
    .C(_05121_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29190_ (.A1(net18078),
    .A2(net19104),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29191_ (.A1(_04832_),
    .A2(_05123_),
    .B(_04651_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29192_ (.A1(_05122_),
    .A2(_05124_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29193_ (.A1(_05125_),
    .A2(_05120_),
    .B(_04794_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29194_ (.A1(net18507),
    .A2(net18066),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _29195_ (.A1(_04651_),
    .A2(_04598_),
    .A3(_05127_),
    .A4(net19581),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29196_ (.A1(net18055),
    .A2(net19104),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29197_ (.A1(_05117_),
    .A2(net17677),
    .B(_05060_),
    .C(_05129_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29198_ (.A1(_05128_),
    .A2(_05130_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29199_ (.I(_04634_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29200_ (.A1(_05132_),
    .A2(net18071),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29201_ (.A1(net652),
    .A2(net19081),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29202_ (.A1(_05133_),
    .A2(_05134_),
    .A3(net19599),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29203_ (.A1(net19109),
    .A2(net19617),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29204_ (.A1(net18501),
    .A2(net19579),
    .A3(_05136_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29205_ (.A1(_05135_),
    .A2(_05137_),
    .B(_04651_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29206_ (.A1(_05131_),
    .A2(_05138_),
    .B(net20193),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29207_ (.A1(_05139_),
    .A2(_05126_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29208_ (.A1(_05140_),
    .A2(_05110_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29209_ (.A1(_05004_),
    .A2(net19574),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29210_ (.A1(_04803_),
    .A2(net17681),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29211_ (.A1(_05141_),
    .A2(net18500),
    .A3(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29212_ (.A1(_05041_),
    .A2(net19070),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29213_ (.A1(net18055),
    .A2(net19088),
    .B(net19581),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29214_ (.A1(_05144_),
    .A2(_05145_),
    .B(net19948),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29215_ (.A1(_05143_),
    .A2(_05146_),
    .B(net20192),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29216_ (.A1(net19080),
    .A2(net19101),
    .A3(net19079),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29217_ (.A1(net17391),
    .A2(net18496),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29218_ (.A1(_05148_),
    .A2(_05149_),
    .B(net19588),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29219_ (.A1(_05020_),
    .A2(net19588),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29220_ (.A1(_04936_),
    .A2(_05151_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29221_ (.A1(_05150_),
    .A2(_05152_),
    .B(net19948),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29222_ (.A1(_05153_),
    .A2(_05147_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29223_ (.A1(_04797_),
    .A2(net19088),
    .Z(_05155_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29224_ (.I(_05012_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29225_ (.A1(_05155_),
    .A2(_05156_),
    .B(net19949),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29226_ (.A1(net18063),
    .A2(net19102),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29227_ (.A1(_05157_),
    .A2(_05158_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29228_ (.A1(_05159_),
    .A2(net19594),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29229_ (.A1(_16092_[0]),
    .A2(_16101_[0]),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29230_ (.A1(net19085),
    .A2(_05161_),
    .B(_04651_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29231_ (.A1(_04896_),
    .A2(_04707_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29232_ (.A1(_05162_),
    .A2(_05163_),
    .B(net19595),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29233_ (.A1(net18070),
    .A2(net19097),
    .B(net19945),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29234_ (.A1(_04856_),
    .A2(_04767_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29235_ (.A1(_05165_),
    .A2(_04929_),
    .A3(_05166_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29236_ (.A1(_05164_),
    .A2(_05167_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29237_ (.A1(_04803_),
    .A2(net19071),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29238_ (.A1(net18073),
    .A2(net19101),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29239_ (.A1(_05169_),
    .A2(_05170_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29240_ (.A1(_05171_),
    .A2(net19061),
    .B(net20400),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29241_ (.A1(_05160_),
    .A2(_05168_),
    .A3(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29242_ (.A1(_05154_),
    .A2(_05173_),
    .A3(_04794_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29243_ (.A1(net19102),
    .A2(net18496),
    .B(_05004_),
    .C(net17679),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29244_ (.A1(net18491),
    .A2(net19593),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29245_ (.A1(_05176_),
    .A2(net18081),
    .B(net19948),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29246_ (.A1(_05175_),
    .A2(net19594),
    .B(_05177_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _29247_ (.A1(_04966_),
    .A2(net19088),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29248_ (.A1(_05179_),
    .A2(net18489),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29249_ (.A1(_05180_),
    .A2(net19573),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29250_ (.A1(_04856_),
    .A2(net19069),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29251_ (.A1(_05179_),
    .A2(net19594),
    .A3(_05182_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29252_ (.A1(_05181_),
    .A2(_05183_),
    .A3(net19948),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29253_ (.A1(_05178_),
    .A2(_05184_),
    .A3(net20192),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29254_ (.A1(net18068),
    .A2(net19588),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29255_ (.A1(_05062_),
    .A2(_05186_),
    .B(net19945),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29256_ (.A1(_04918_),
    .A2(net19573),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29257_ (.A1(_05187_),
    .A2(_05188_),
    .B(net20191),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29258_ (.I(_16093_[0]),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29259_ (.A1(_05190_),
    .A2(net19108),
    .B(net19588),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29260_ (.A1(_05133_),
    .A2(_05191_),
    .B(_04651_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29261_ (.A1(_05111_),
    .A2(net19089),
    .B(net18492),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29262_ (.A1(_05193_),
    .A2(net19596),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29263_ (.A1(_05192_),
    .A2(_05194_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29264_ (.A1(_05189_),
    .A2(_05195_),
    .B(_04794_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29265_ (.A1(_05185_),
    .A2(_05196_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29266_ (.A1(_05174_),
    .A2(_05197_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29267_ (.A1(net18502),
    .A2(net19100),
    .A3(net18498),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29268_ (.A1(net18060),
    .A2(_04769_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29269_ (.A1(_05199_),
    .A2(_05198_),
    .A3(net19947),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29270_ (.A1(_05009_),
    .A2(_04837_),
    .A3(_04651_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29271_ (.A1(net19592),
    .A2(_05200_),
    .A3(_05201_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29272_ (.A1(_04940_),
    .A2(_05166_),
    .A3(_04651_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29273_ (.A1(_04856_),
    .A2(_04651_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29274_ (.A1(_05062_),
    .A2(_05204_),
    .B(net19592),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29275_ (.A1(_05203_),
    .A2(_05205_),
    .B(net20400),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29276_ (.A1(_05206_),
    .A2(_05202_),
    .B(_04794_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29277_ (.A1(net19082),
    .A2(net19608),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29278_ (.A1(_05042_),
    .A2(_05208_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29279_ (.A1(_05209_),
    .A2(net19590),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29280_ (.A1(_05132_),
    .A2(_04700_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29281_ (.A1(_05211_),
    .A2(net19580),
    .A3(_04950_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29282_ (.A1(_05210_),
    .A2(_05212_),
    .A3(net19946),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29283_ (.A1(net19084),
    .A2(_04978_),
    .B(_05020_),
    .C(net19579),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29284_ (.A1(net19063),
    .A2(net19105),
    .B(net19571),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29285_ (.A1(net18503),
    .A2(net18057),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29286_ (.A1(_05215_),
    .A2(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29287_ (.A1(_05214_),
    .A2(net19585),
    .A3(_05217_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29288_ (.A1(_05213_),
    .A2(_05218_),
    .A3(net20400),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29289_ (.A1(_05219_),
    .A2(_05207_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _29290_ (.A1(net18060),
    .A2(net19079),
    .B1(net17392),
    .B2(net18495),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29291_ (.A1(_05221_),
    .A2(net19590),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29292_ (.A1(net19108),
    .A2(_16101_[0]),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29293_ (.A1(_04884_),
    .A2(_05223_),
    .A3(net19588),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29294_ (.A1(net17682),
    .A2(net19093),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29295_ (.A1(_05224_),
    .A2(_05225_),
    .B(net19946),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29296_ (.A1(_05222_),
    .A2(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29297_ (.A1(_05077_),
    .A2(net19070),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29298_ (.A1(_05228_),
    .A2(net19588),
    .A3(_04847_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29299_ (.A1(net19101),
    .A2(_05053_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29300_ (.A1(_04786_),
    .A2(_05230_),
    .B(_04651_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29301_ (.A1(_05229_),
    .A2(_05231_),
    .B(_04691_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29302_ (.A1(_05227_),
    .A2(_05232_),
    .B(net20190),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29303_ (.A1(_04823_),
    .A2(_04805_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29304_ (.A1(_04995_),
    .A2(_05234_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29305_ (.A1(_05235_),
    .A2(net19595),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29306_ (.A1(_04700_),
    .A2(_04716_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29307_ (.A1(_05237_),
    .A2(net19089),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29308_ (.A1(_04662_),
    .A2(_04982_),
    .B(net19600),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29309_ (.A1(_05239_),
    .A2(_05238_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29310_ (.A1(net19951),
    .A2(_05240_),
    .A3(_05236_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29311_ (.I(_05163_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29312_ (.A1(_05242_),
    .A2(_04814_),
    .B(net19595),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29313_ (.A1(net18491),
    .A2(_05068_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29314_ (.A1(_05244_),
    .A2(_05033_),
    .B(net19945),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29315_ (.A1(_05243_),
    .A2(_05245_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29316_ (.A1(_05246_),
    .A2(_05241_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29317_ (.A1(net20193),
    .A2(_05247_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29318_ (.A1(_05233_),
    .A2(_05248_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29319_ (.A1(_05249_),
    .A2(_05220_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29320_ (.A1(_02288_),
    .A2(net20873),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29321_ (.A1(_11215_),
    .A2(_02285_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29322_ (.A1(_05250_),
    .A2(_05251_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29323_ (.I(_05252_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29324_ (.A1(_11156_),
    .A2(net21358),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29325_ (.A1(_11152_),
    .A2(net21046),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29326_ (.A1(_05254_),
    .A2(_05255_),
    .Z(_05256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29327_ (.A1(_05253_),
    .A2(_05256_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29328_ (.A1(_05254_),
    .A2(_05255_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29329_ (.A1(_05252_),
    .A2(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29330_ (.A1(_05257_),
    .A2(net21068),
    .A3(_05259_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29331_ (.A1(net21504),
    .A2(\text_in_r[65] ),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29332_ (.A1(net19944),
    .A2(net21199),
    .A3(net20964),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29333_ (.A1(_05253_),
    .A2(_05258_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29334_ (.A1(_05256_),
    .A2(_05252_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29335_ (.A1(_05263_),
    .A2(_05264_),
    .A3(net21068),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29336_ (.A1(net21068),
    .A2(\text_in_r[65] ),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29337_ (.A1(net19943),
    .A2(_07791_),
    .A3(net20928),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29338_ (.A1(_05267_),
    .A2(_05262_),
    .ZN(_16111_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29339_ (.A1(_11193_),
    .A2(_11195_),
    .A3(net21287),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29340_ (.A1(net21043),
    .A2(net21041),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29341_ (.A1(net21411),
    .A2(net21360),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29342_ (.A1(_05269_),
    .A2(net20968),
    .A3(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29343_ (.A1(_05268_),
    .A2(_05271_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29344_ (.A1(_05272_),
    .A2(net20910),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29345_ (.A1(_05268_),
    .A2(_05271_),
    .A3(net20911),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29346_ (.A1(_05273_),
    .A2(_05274_),
    .B(net21501),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29347_ (.I(\text_in_r[64] ),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29348_ (.A1(_05276_),
    .A2(net21501),
    .Z(_05277_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29349_ (.A1(net20399),
    .A2(net20927),
    .B(net21208),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29350_ (.A1(_05273_),
    .A2(_05274_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29351_ (.A1(_05279_),
    .A2(net21068),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29352_ (.I(_05277_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29353_ (.A1(net20186),
    .A2(net21109),
    .A3(net20865),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29354_ (.A1(_05278_),
    .A2(_05282_),
    .ZN(_16114_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29355_ (.A1(net21296),
    .A2(\sa21_sr[2] ),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29356_ (.A1(net21296),
    .A2(\sa21_sr[2] ),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29357_ (.A1(_05283_),
    .A2(_05284_),
    .B(net21465),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29358_ (.A1(net21045),
    .A2(_11216_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29359_ (.A1(net21296),
    .A2(\sa21_sr[2] ),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29360_ (.A1(_05286_),
    .A2(_11250_),
    .A3(_05287_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29361_ (.A1(_05285_),
    .A2(_05288_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _29362_ (.A1(net21466),
    .A2(\sa11_sr[2] ),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29363_ (.I(_05290_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29364_ (.A1(_05289_),
    .A2(_05291_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29365_ (.A1(_05285_),
    .A2(_05288_),
    .A3(_05290_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29366_ (.A1(_05292_),
    .A2(_05293_),
    .B(net21501),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29367_ (.I(\text_in_r[66] ),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29368_ (.A1(_05295_),
    .A2(net21501),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _29369_ (.A1(_05294_),
    .A2(_05296_),
    .B(net21189),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29370_ (.A1(_05292_),
    .A2(_05293_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29371_ (.A1(_05298_),
    .A2(net21068),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29372_ (.I(_05296_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29373_ (.A1(_05299_),
    .A2(_07796_),
    .A3(_05300_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29374_ (.A1(_05297_),
    .A2(_05301_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _29375_ (.I(_05302_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input132 (.I(net573),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29377_ (.A1(_05275_),
    .A2(_05277_),
    .B(_07782_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29378_ (.A1(_05280_),
    .A2(net21208),
    .A3(_05281_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29379_ (.A1(_05304_),
    .A2(_05305_),
    .ZN(_16105_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input131 (.I(text_in[0]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input130 (.I(net560),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29382_ (.A1(_05303_),
    .A2(net19565),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29383_ (.A1(_11257_),
    .A2(net21353),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29384_ (.A1(_11253_),
    .A2(net21034),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29385_ (.A1(_05308_),
    .A2(_05309_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29386_ (.A1(net20420),
    .A2(_05310_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29387_ (.I(_05310_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29388_ (.A1(net20419),
    .A2(_05312_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29389_ (.A1(_05311_),
    .A2(_05313_),
    .A3(net21068),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29390_ (.A1(net21503),
    .A2(\text_in_r[67] ),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29391_ (.A1(_05314_),
    .A2(_07801_),
    .A3(_05315_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29392_ (.A1(net20420),
    .A2(_05312_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29393_ (.A1(net20419),
    .A2(_05310_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29394_ (.A1(_05317_),
    .A2(net21068),
    .A3(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _29395_ (.A1(net21070),
    .A2(\text_in_r[67] ),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29396_ (.A1(_05319_),
    .A2(net21188),
    .A3(_05320_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29397_ (.A1(_05316_),
    .A2(_05321_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input129 (.I(ld),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29399_ (.A1(_05307_),
    .A2(net19038),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29400_ (.A1(net21351),
    .A2(_11301_),
    .Z(_05325_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29401_ (.A1(_05325_),
    .A2(net20803),
    .B(net21067),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29402_ (.A1(_05325_),
    .A2(net20803),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29403_ (.I(_05327_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29404_ (.A1(net21505),
    .A2(\text_in_r[68] ),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29405_ (.A1(_05326_),
    .A2(_05328_),
    .B(_05329_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29406_ (.A1(net20184),
    .A2(net21187),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29407_ (.A1(_05325_),
    .A2(net20803),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29408_ (.A1(_05332_),
    .A2(net21067),
    .A3(_05327_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29409_ (.A1(net20398),
    .A2(_07808_),
    .A3(net20963),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29410_ (.A1(_05331_),
    .A2(_05334_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input128 (.I(key[9]),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29412_ (.A1(net18054),
    .A2(net19559),
    .Z(_05337_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29413_ (.I(_16112_[0]),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29414_ (.A1(net19567),
    .A2(_05338_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29415_ (.A1(_05314_),
    .A2(net21188),
    .A3(_05315_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29416_ (.A1(_05319_),
    .A2(_07801_),
    .A3(_05320_),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29417_ (.A1(_05340_),
    .A2(_05341_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input127 (.I(net548),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29419_ (.A1(_05339_),
    .A2(net19022),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29420_ (.A1(net19060),
    .A2(net19057),
    .A3(net19566),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29421_ (.A1(_05344_),
    .A2(net18484),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _29422_ (.A1(net21290),
    .A2(\sa21_sr[5] ),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29423_ (.A1(_05347_),
    .A2(net21460),
    .Z(_05348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29424_ (.A1(_05347_),
    .A2(net21460),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29425_ (.A1(_05348_),
    .A2(_05349_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29426_ (.A1(net21461),
    .A2(\sa11_sr[5] ),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29427_ (.A1(_05350_),
    .A2(_05351_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29428_ (.A1(_05350_),
    .A2(_05351_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29429_ (.A1(net21505),
    .A2(\text_in_r[69] ),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _29430_ (.A1(_05352_),
    .A2(net21505),
    .A3(_05353_),
    .B(_05354_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29431_ (.A1(_05355_),
    .A2(net21186),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29432_ (.A1(_05355_),
    .A2(net21186),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29433_ (.A1(_05356_),
    .A2(_05357_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input126 (.I(key[98]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29435_ (.A1(_05337_),
    .A2(_05346_),
    .B(net20182),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29436_ (.A1(_05302_),
    .A2(net19565),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29437_ (.A1(net19020),
    .A2(net19052),
    .Z(_05362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29438_ (.A1(net19060),
    .A2(net19566),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29439_ (.A1(_05362_),
    .A2(net18483),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29440_ (.A1(_05330_),
    .A2(_07808_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29441_ (.A1(_05333_),
    .A2(net21187),
    .A3(_05329_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29442_ (.A1(_05365_),
    .A2(_05366_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input125 (.I(key[97]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input124 (.I(net554),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _29445_ (.I(_16121_[0]),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29446_ (.A1(_05370_),
    .A2(_05303_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input123 (.I(key[95]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29448_ (.I(_16108_[0]),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29449_ (.A1(_05373_),
    .A2(net19567),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29450_ (.A1(net17674),
    .A2(net19032),
    .A3(net17671),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29451_ (.A1(_05364_),
    .A2(net19554),
    .A3(_05375_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29452_ (.A1(net21289),
    .A2(net21348),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29453_ (.A1(\sa01_sr[6] ),
    .A2(_05377_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29454_ (.A1(net21460),
    .A2(net21404),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29455_ (.A1(_05378_),
    .A2(_05379_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29456_ (.A1(_05378_),
    .A2(_05379_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29457_ (.A1(net21505),
    .A2(\text_in_r[70] ),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _29458_ (.A1(_05380_),
    .A2(net21505),
    .A3(_05381_),
    .B(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29459_ (.A1(_05383_),
    .A2(net21185),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29460_ (.A1(_05383_),
    .A2(net21185),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29461_ (.A1(_05384_),
    .A2(_05385_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input122 (.I(key[94]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29463_ (.A1(_05360_),
    .A2(_05376_),
    .B(net20397),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29464_ (.A1(_05265_),
    .A2(net21199),
    .A3(_05266_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29465_ (.A1(_07791_),
    .A2(_05260_),
    .A3(_05261_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29466_ (.A1(_05389_),
    .A2(_05390_),
    .ZN(_16106_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29467_ (.A1(net19019),
    .A2(_05303_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29468_ (.A1(_05303_),
    .A2(net19570),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29469_ (.A1(_05391_),
    .A2(_05392_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29470_ (.A1(net19060),
    .A2(net19568),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input121 (.I(key[93]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29472_ (.A1(_05394_),
    .A2(net19050),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29473_ (.A1(_05393_),
    .A2(_05396_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29474_ (.A1(net19567),
    .A2(_05370_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input120 (.I(key[92]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input119 (.I(key[91]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29477_ (.A1(net18486),
    .A2(net17669),
    .B(net19046),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29478_ (.A1(_05397_),
    .A2(_05401_),
    .B(net19551),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29479_ (.A1(net19060),
    .A2(net19570),
    .A3(net19567),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input118 (.I(key[90]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29481_ (.A1(_05403_),
    .A2(net19023),
    .A3(net18485),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29482_ (.A1(net19567),
    .A2(net18374),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29483_ (.A1(net18482),
    .A2(net18049),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29484_ (.A1(_05407_),
    .A2(net19046),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input117 (.I(key[8]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29486_ (.A1(_05405_),
    .A2(_05408_),
    .A3(net19562),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input116 (.I(key[89]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input115 (.I(key[88]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29489_ (.A1(_05402_),
    .A2(_05410_),
    .A3(net20182),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29490_ (.A1(net21288),
    .A2(net20908),
    .Z(_05414_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _29491_ (.A1(_14478_),
    .A2(net689),
    .A3(_05414_),
    .Z(_05415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29492_ (.A1(net21501),
    .A2(\text_in_r[71] ),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29493_ (.A1(_05415_),
    .A2(net21078),
    .B(_05416_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _29494_ (.A1(net21184),
    .A2(_05417_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29495_ (.I(_05418_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29496_ (.A1(_05388_),
    .A2(_05413_),
    .B(_05419_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29497_ (.A1(net19060),
    .A2(_05303_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29498_ (.A1(net19567),
    .A2(net18376),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29499_ (.A1(_05421_),
    .A2(net19053),
    .A3(net18048),
    .Z(_05423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29500_ (.A1(_05303_),
    .A2(net18052),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29501_ (.A1(net19022),
    .A2(_05424_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29502_ (.A1(_05423_),
    .A2(net19561),
    .A3(_05425_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29503_ (.A1(net19022),
    .A2(_05374_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _29504_ (.I(_05427_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29505_ (.A1(net19056),
    .A2(net18377),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29506_ (.A1(_05428_),
    .A2(_05429_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _29507_ (.I(_16115_[0]),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29508_ (.A1(net19567),
    .A2(_05431_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29509_ (.A1(_05432_),
    .A2(net19022),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29510_ (.A1(net19567),
    .A2(net18377),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29511_ (.A1(net17389),
    .A2(net18044),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input114 (.I(key[87]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29513_ (.A1(_05430_),
    .A2(_05435_),
    .B(net19554),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29514_ (.A1(_05426_),
    .A2(_05437_),
    .B(net20183),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29515_ (.A1(net17672),
    .A2(net19038),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29516_ (.A1(net19060),
    .A2(_05303_),
    .A3(net19570),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29517_ (.A1(_05439_),
    .A2(net18471),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29518_ (.I(_16107_[0]),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29519_ (.A1(net19055),
    .A2(_05442_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29520_ (.A1(net19568),
    .A2(net18046),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29521_ (.A1(net17665),
    .A2(_05444_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input113 (.I(key[86]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29523_ (.A1(_05445_),
    .A2(net19027),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input112 (.I(key[85]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29525_ (.A1(_05441_),
    .A2(_05447_),
    .A3(net19559),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29526_ (.A1(_05302_),
    .A2(net19570),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29527_ (.A1(_05450_),
    .A2(net19038),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29528_ (.A1(net19019),
    .A2(net19566),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29529_ (.A1(_05451_),
    .A2(net18470),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input111 (.I(key[84]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29531_ (.A1(_05363_),
    .A2(_05392_),
    .A3(net19027),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29532_ (.A1(_05453_),
    .A2(_05455_),
    .A3(net19553),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 _29533_ (.I(_05358_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input110 (.I(key[83]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29535_ (.A1(_05449_),
    .A2(_05456_),
    .A3(net19934),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29536_ (.A1(_05438_),
    .A2(_05459_),
    .A3(net20397),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29537_ (.A1(_05420_),
    .A2(_05460_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29538_ (.A1(net18485),
    .A2(net19022),
    .A3(_05434_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29539_ (.A1(_05462_),
    .A2(net19559),
    .Z(_05463_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29540_ (.A1(_05303_),
    .A2(net18375),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _29541_ (.A1(_05464_),
    .A2(net19022),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29542_ (.I(_05361_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29543_ (.A1(_05466_),
    .A2(net19060),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29544_ (.A1(net20185),
    .A2(net19942),
    .A3(net18053),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29545_ (.A1(_05467_),
    .A2(net19046),
    .A3(_05468_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29546_ (.A1(_05463_),
    .A2(_05465_),
    .A3(_05469_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _29547_ (.A1(net20185),
    .A2(net19942),
    .A3(net18376),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29548_ (.A1(_05471_),
    .A2(net19038),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input109 (.I(key[82]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29550_ (.A1(net19047),
    .A2(_16128_[0]),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _29551_ (.A1(_05472_),
    .A2(_05474_),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input108 (.I(key[81]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29553_ (.A1(_05475_),
    .A2(net19549),
    .B(_05457_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29554_ (.A1(_05470_),
    .A2(_05477_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _29555_ (.A1(net19567),
    .A2(_16117_[0]),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _29556_ (.A1(_05479_),
    .A2(net19038),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29557_ (.A1(_05467_),
    .A2(net17664),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29558_ (.I(_05406_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29559_ (.A1(net17663),
    .A2(net19046),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29560_ (.A1(_05481_),
    .A2(net19562),
    .A3(_05483_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29561_ (.A1(_05482_),
    .A2(net19022),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29562_ (.A1(_05485_),
    .A2(net19546),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29563_ (.A1(_05467_),
    .A2(net17390),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29564_ (.A1(_05486_),
    .A2(_05487_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input107 (.I(key[80]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29566_ (.A1(_05484_),
    .A2(_05488_),
    .A3(net19935),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29567_ (.A1(_05478_),
    .A2(_05490_),
    .A3(net20397),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _29568_ (.I(_05443_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29569_ (.A1(_05492_),
    .A2(net17663),
    .B(net19050),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input106 (.I(key[7]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29571_ (.A1(_05344_),
    .A2(net19559),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29572_ (.A1(_05493_),
    .A2(_05495_),
    .B(net20182),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29573_ (.A1(_05394_),
    .A2(net19050),
    .A3(_05471_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29574_ (.A1(_05497_),
    .A2(net19559),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29575_ (.I(net17666),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29576_ (.A1(_05499_),
    .A2(net19029),
    .A3(net19020),
    .Z(_05500_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29577_ (.A1(_05498_),
    .A2(_05500_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29578_ (.A1(_05496_),
    .A2(_05501_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29579_ (.A1(net20185),
    .A2(net19942),
    .A3(net18372),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _29580_ (.I(_05503_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29581_ (.A1(_05504_),
    .A2(net19046),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29582_ (.A1(_05405_),
    .A2(net17386),
    .A3(net19562),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input105 (.I(key[79]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29584_ (.A1(_05427_),
    .A2(net19546),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29585_ (.A1(net19567),
    .A2(_16117_[0]),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29586_ (.A1(net18040),
    .A2(_05503_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29587_ (.A1(_05510_),
    .A2(net19039),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29588_ (.A1(_05508_),
    .A2(_05511_),
    .B(_05457_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29589_ (.A1(_05506_),
    .A2(_05512_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _29590_ (.I(_05386_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input104 (.I(key[78]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29592_ (.A1(_05502_),
    .A2(_05513_),
    .A3(net20179),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29593_ (.A1(_05491_),
    .A2(_05516_),
    .A3(net19940),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29594_ (.A1(_05461_),
    .A2(_05517_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29595_ (.A1(net19022),
    .A2(_05303_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input103 (.I(key[77]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29597_ (.A1(_05518_),
    .A2(net18483),
    .B(net19546),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29598_ (.A1(_05394_),
    .A2(_05452_),
    .A3(net19051),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29599_ (.A1(_05520_),
    .A2(_05521_),
    .B(net20183),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29600_ (.A1(_05339_),
    .A2(net19044),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29601_ (.A1(_05523_),
    .A2(net18478),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29602_ (.A1(_05428_),
    .A2(net18486),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29603_ (.A1(_05524_),
    .A2(_05525_),
    .A3(net19550),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29604_ (.A1(_05522_),
    .A2(_05526_),
    .B(_05514_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29605_ (.A1(_05421_),
    .A2(net19022),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29606_ (.A1(net19019),
    .A2(net19568),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29607_ (.A1(_05528_),
    .A2(_05529_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29608_ (.A1(_05505_),
    .A2(net19554),
    .Z(_05531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29609_ (.A1(_05530_),
    .A2(_05531_),
    .B(_05457_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29610_ (.A1(_05425_),
    .A2(net17668),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29611_ (.A1(_05469_),
    .A2(_05533_),
    .A3(net19562),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29612_ (.A1(_05532_),
    .A2(_05534_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input102 (.I(key[76]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29614_ (.A1(_05527_),
    .A2(_05535_),
    .B(net20180),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29615_ (.A1(net18477),
    .A2(net19049),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29616_ (.A1(net19568),
    .A2(_05442_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29617_ (.I(_05539_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _29618_ (.A1(_05538_),
    .A2(net17385),
    .B1(_05427_),
    .B2(_05504_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input101 (.I(key[75]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29620_ (.A1(_05541_),
    .A2(net19558),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29621_ (.A1(net19060),
    .A2(net19570),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input100 (.I(key[74]),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29623_ (.A1(_05544_),
    .A2(net18469),
    .B(net19025),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29624_ (.A1(_05472_),
    .A2(net19020),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29625_ (.A1(_05546_),
    .A2(net19559),
    .A3(_05547_),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29626_ (.A1(_05543_),
    .A2(net20182),
    .A3(_05548_),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29627_ (.A1(_05440_),
    .A2(net19030),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _29628_ (.I(_05422_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _29629_ (.A1(_05550_),
    .A2(_05551_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29630_ (.A1(net19567),
    .A2(net18373),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29631_ (.I(_05553_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input99 (.I(key[73]),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29633_ (.A1(_05554_),
    .A2(net19042),
    .B(net19546),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29634_ (.A1(_05552_),
    .A2(_05556_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29635_ (.A1(_05371_),
    .A2(net19022),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29636_ (.I(_05558_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29637_ (.A1(_05559_),
    .A2(net18468),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29638_ (.A1(_05529_),
    .A2(net19020),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input98 (.I(key[72]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29640_ (.A1(_05561_),
    .A2(net19046),
    .ZN(_05563_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input97 (.I(key[71]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29642_ (.A1(_05560_),
    .A2(_05563_),
    .A3(net19547),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29643_ (.A1(_05557_),
    .A2(_05565_),
    .A3(net19938),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29644_ (.A1(_05549_),
    .A2(net20179),
    .A3(_05566_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29645_ (.A1(_05537_),
    .A2(_05567_),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29646_ (.A1(_05398_),
    .A2(net19046),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29647_ (.I(_16109_[0]),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29648_ (.A1(_05303_),
    .A2(_05570_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29649_ (.A1(_05569_),
    .A2(net17659),
    .B(net19559),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29650_ (.A1(_05552_),
    .A2(_05572_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _29651_ (.I(_05324_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29652_ (.A1(_05574_),
    .A2(net18474),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29653_ (.A1(_05427_),
    .A2(net19559),
    .Z(_05576_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29654_ (.A1(_05575_),
    .A2(_05576_),
    .B(_05457_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29655_ (.A1(_05573_),
    .A2(_05577_),
    .B(net20397),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29656_ (.A1(_05425_),
    .A2(net18044),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29657_ (.A1(net19038),
    .A2(net19056),
    .A3(net19570),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29658_ (.A1(_05580_),
    .A2(net19546),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29659_ (.I(_05581_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29660_ (.A1(_05579_),
    .A2(_05582_),
    .A3(_05483_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29661_ (.A1(_05451_),
    .A2(net18047),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _29662_ (.A1(_05344_),
    .A2(net18480),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29663_ (.A1(_05584_),
    .A2(_05585_),
    .A3(net19562),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29664_ (.A1(_05583_),
    .A2(_05586_),
    .A3(net19935),
    .ZN(_05587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29665_ (.A1(_05578_),
    .A2(_05587_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29666_ (.A1(_05362_),
    .A2(_05429_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29667_ (.A1(_05589_),
    .A2(_05457_),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29668_ (.A1(net18050),
    .A2(_05561_),
    .B(net19034),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29669_ (.A1(_05590_),
    .A2(_05591_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29670_ (.A1(_05451_),
    .A2(_05421_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29671_ (.A1(_05593_),
    .A2(_05585_),
    .A3(net20183),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29672_ (.A1(_05592_),
    .A2(net19555),
    .A3(_05594_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _29673_ (.I(_16131_[0]),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29674_ (.A1(net19032),
    .A2(_05596_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29675_ (.A1(_05433_),
    .A2(_05403_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29676_ (.A1(_05457_),
    .A2(_05597_),
    .B(net17237),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input96 (.I(key[70]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29678_ (.A1(_05599_),
    .A2(net19563),
    .B(_05514_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29679_ (.A1(_05595_),
    .A2(_05601_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29680_ (.A1(_05588_),
    .A2(_05602_),
    .A3(net20181),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29681_ (.A1(_05568_),
    .A2(_05603_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29682_ (.A1(_05467_),
    .A2(_05468_),
    .B(net19046),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29683_ (.A1(_05604_),
    .A2(_05498_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29684_ (.A1(_05523_),
    .A2(net17674),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29685_ (.A1(net18475),
    .A2(_05363_),
    .A3(net19027),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input95 (.I(key[6]),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29687_ (.A1(_05606_),
    .A2(_05607_),
    .B(net19559),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29688_ (.A1(_05605_),
    .A2(_05609_),
    .B(net20182),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29689_ (.A1(net18484),
    .A2(net19050),
    .B(net19546),
    .ZN(_05611_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29690_ (.A1(net18471),
    .A2(net19026),
    .A3(net17669),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29691_ (.A1(_05611_),
    .A2(_05612_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29692_ (.A1(_05464_),
    .A2(net19015),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29693_ (.A1(_05614_),
    .A2(net19026),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29694_ (.A1(_05421_),
    .A2(net19051),
    .A3(net17673),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29695_ (.A1(_05615_),
    .A2(_05616_),
    .A3(net19552),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29696_ (.A1(_05613_),
    .A2(_05617_),
    .A3(net19933),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29697_ (.A1(_05610_),
    .A2(net20397),
    .A3(_05618_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _29698_ (.A1(_05479_),
    .A2(net19022),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29699_ (.A1(_05620_),
    .A2(net19021),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29700_ (.A1(_05471_),
    .A2(net19022),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29701_ (.A1(_05622_),
    .A2(net17671),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29702_ (.A1(_05621_),
    .A2(_05623_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29703_ (.A1(_05624_),
    .A2(net19559),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29704_ (.A1(net18481),
    .A2(net19022),
    .A3(net18040),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29705_ (.A1(net20185),
    .A2(net19942),
    .A3(net18371),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29706_ (.A1(net19015),
    .A2(net19039),
    .A3(_05627_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29707_ (.A1(_05626_),
    .A2(net19557),
    .A3(_05628_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29708_ (.A1(_05625_),
    .A2(_05629_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29709_ (.A1(_05630_),
    .A2(net19939),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29710_ (.A1(net19015),
    .A2(net18042),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29711_ (.A1(_05627_),
    .A2(net19039),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29712_ (.A1(_05632_),
    .A2(net19040),
    .B(_05633_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29713_ (.I(_05509_),
    .ZN(_05635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29714_ (.A1(net17657),
    .A2(net19040),
    .B(net19559),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29715_ (.A1(_05634_),
    .A2(_05636_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29716_ (.A1(_05529_),
    .A2(net19023),
    .A3(_05468_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29717_ (.A1(_05638_),
    .A2(_05511_),
    .A3(net19559),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29718_ (.A1(_05637_),
    .A2(_05639_),
    .A3(net20182),
    .ZN(_05640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29719_ (.A1(_05631_),
    .A2(_05514_),
    .A3(_05640_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29720_ (.A1(_05619_),
    .A2(_05641_),
    .A3(net20180),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29721_ (.A1(_05425_),
    .A2(_05467_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29722_ (.A1(_16128_[0]),
    .A2(net19047),
    .B(net19546),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29723_ (.A1(_05643_),
    .A2(_05644_),
    .B(net20182),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _29724_ (.A1(net19019),
    .A2(_05303_),
    .B(net19038),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29725_ (.A1(_05646_),
    .A2(net19020),
    .ZN(_05647_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29726_ (.A1(_05647_),
    .A2(net19551),
    .A3(net17662),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29727_ (.A1(_05645_),
    .A2(_05648_),
    .B(net20397),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29728_ (.A1(_05622_),
    .A2(_05444_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29729_ (.A1(_05396_),
    .A2(_05492_),
    .B(_05650_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29730_ (.A1(_05651_),
    .A2(net19552),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29731_ (.A1(net18475),
    .A2(_05452_),
    .A3(net19027),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29732_ (.A1(_05653_),
    .A2(net19559),
    .Z(_05654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29733_ (.A1(net19051),
    .A2(_05596_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29734_ (.A1(_05654_),
    .A2(_05655_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29735_ (.A1(_05652_),
    .A2(_05656_),
    .A3(net20182),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29736_ (.A1(_05649_),
    .A2(_05657_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29737_ (.A1(_05598_),
    .A2(net19546),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29738_ (.A1(_05391_),
    .A2(net18485),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29739_ (.A1(net18049),
    .A2(_05553_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29740_ (.A1(_05660_),
    .A2(_05661_),
    .B(net19028),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29741_ (.A1(_05659_),
    .A2(_05662_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29742_ (.A1(_05540_),
    .A2(net19045),
    .B(net19546),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29743_ (.A1(_05428_),
    .A2(_05468_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29744_ (.A1(_05665_),
    .A2(_05664_),
    .B(net20182),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29745_ (.A1(_05663_),
    .A2(_05666_),
    .B(_05514_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29746_ (.A1(_05345_),
    .A2(net19048),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29747_ (.A1(net19038),
    .A2(_16126_[0]),
    .Z(_05669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29748_ (.A1(_05668_),
    .A2(_05669_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29749_ (.A1(_05670_),
    .A2(net19553),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29750_ (.A1(net19048),
    .A2(_16135_[0]),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29751_ (.A1(_05607_),
    .A2(net19553),
    .A3(_05672_),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29752_ (.A1(_05671_),
    .A2(net20182),
    .A3(_05673_),
    .ZN(_05674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29753_ (.A1(_05667_),
    .A2(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29754_ (.A1(_05658_),
    .A2(_05675_),
    .A3(net19941),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29755_ (.A1(_05642_),
    .A2(_05676_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29756_ (.A1(net18466),
    .A2(net17673),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29757_ (.A1(_05451_),
    .A2(net18483),
    .ZN(_05678_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29758_ (.A1(_05677_),
    .A2(_05678_),
    .A3(net19561),
    .ZN(_05679_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29759_ (.I(_05424_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29760_ (.A1(_05680_),
    .A2(net19022),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29761_ (.A1(_05593_),
    .A2(_05681_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29762_ (.A1(_05682_),
    .A2(net19555),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29763_ (.A1(_05679_),
    .A2(_05683_),
    .A3(net20183),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29764_ (.A1(_05392_),
    .A2(net19049),
    .A3(_05444_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29765_ (.A1(net17667),
    .A2(net19025),
    .A3(net17661),
    .ZN(_05686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29766_ (.A1(_05685_),
    .A2(_05686_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29767_ (.A1(_05687_),
    .A2(net19552),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29768_ (.A1(_05422_),
    .A2(net19046),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29769_ (.A1(_05689_),
    .A2(net18480),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29770_ (.A1(net17670),
    .A2(_05468_),
    .A3(net19029),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29771_ (.A1(_05690_),
    .A2(net19560),
    .A3(_05691_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29772_ (.A1(_05688_),
    .A2(_05692_),
    .A3(_05457_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29773_ (.A1(_05684_),
    .A2(net20397),
    .A3(_05693_),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29774_ (.I(_05529_),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29775_ (.A1(_05558_),
    .A2(_05695_),
    .B(net19546),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29776_ (.A1(_05620_),
    .A2(net18048),
    .Z(_05697_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29777_ (.A1(_05696_),
    .A2(_05697_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _29778_ (.A1(_05452_),
    .A2(net18479),
    .A3(net19559),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29779_ (.A1(net19027),
    .A2(net19569),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29780_ (.A1(_05699_),
    .A2(_05700_),
    .B(net19934),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29781_ (.A1(_05698_),
    .A2(_05701_),
    .B(net20397),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29782_ (.A1(_05392_),
    .A2(_05444_),
    .Z(_05703_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29783_ (.A1(_05703_),
    .A2(_05646_),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29784_ (.A1(net19019),
    .A2(net19566),
    .B(net19569),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29785_ (.A1(_05705_),
    .A2(_05472_),
    .ZN(_05706_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29786_ (.A1(_05704_),
    .A2(net19559),
    .A3(_05706_),
    .ZN(_05707_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29787_ (.A1(net19055),
    .A2(_05431_),
    .Z(_05708_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29788_ (.I(_05708_),
    .ZN(_05709_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29789_ (.A1(_05439_),
    .A2(_05709_),
    .ZN(_05710_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29790_ (.A1(_05710_),
    .A2(_05455_),
    .A3(net19553),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29791_ (.A1(_05707_),
    .A2(_05711_),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29792_ (.A1(_05712_),
    .A2(net19934),
    .ZN(_05713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29793_ (.A1(_05702_),
    .A2(_05713_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29794_ (.A1(_05694_),
    .A2(_05714_),
    .A3(net19941),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29795_ (.A1(net17389),
    .A2(net18476),
    .Z(_05716_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29796_ (.I(_05681_),
    .ZN(_05717_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29797_ (.A1(_05716_),
    .A2(_05717_),
    .B(net20183),
    .ZN(_05718_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29798_ (.I(_05374_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29799_ (.A1(_05719_),
    .A2(net19041),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29800_ (.A1(_05358_),
    .A2(_05720_),
    .Z(_05721_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29801_ (.A1(_05721_),
    .A2(_05486_),
    .Z(_05722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29802_ (.A1(_05718_),
    .A2(_05722_),
    .B(_05514_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29803_ (.A1(_05574_),
    .A2(net17671),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29804_ (.A1(_05570_),
    .A2(_05338_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29805_ (.A1(_05725_),
    .A2(net19567),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29806_ (.A1(_05726_),
    .A2(net19035),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29807_ (.A1(_05727_),
    .A2(net17675),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29808_ (.A1(_05724_),
    .A2(net20183),
    .A3(_05728_),
    .ZN(_05729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29809_ (.A1(net17657),
    .A2(net19023),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29810_ (.A1(_05621_),
    .A2(_05457_),
    .A3(_05730_),
    .ZN(_05731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29811_ (.A1(_05729_),
    .A2(_05731_),
    .ZN(_05732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29812_ (.A1(_05732_),
    .A2(net19563),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29813_ (.A1(_05723_),
    .A2(_05733_),
    .ZN(_05734_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _29814_ (.I(_05307_),
    .ZN(_05735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _29815_ (.A1(_05735_),
    .A2(net17657),
    .B(net19035),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29816_ (.A1(_05439_),
    .A2(net17674),
    .ZN(_05737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29817_ (.A1(_05736_),
    .A2(_05737_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29818_ (.A1(_05738_),
    .A2(net19547),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29819_ (.A1(_05521_),
    .A2(_05462_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29820_ (.A1(_05740_),
    .A2(net19562),
    .ZN(_05741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29821_ (.A1(_05739_),
    .A2(net19938),
    .A3(_05741_),
    .ZN(_05742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29822_ (.A1(_05480_),
    .A2(_05726_),
    .ZN(_05743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29823_ (.A1(_05598_),
    .A2(_05743_),
    .ZN(_05744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29824_ (.A1(_05744_),
    .A2(net19559),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29825_ (.A1(_05628_),
    .A2(net19546),
    .B(_05457_),
    .ZN(_05746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29826_ (.A1(_05745_),
    .A2(_05746_),
    .B(net20397),
    .ZN(_05747_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29827_ (.A1(_05742_),
    .A2(_05747_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29828_ (.A1(_05734_),
    .A2(_05748_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29829_ (.A1(_05749_),
    .A2(net20181),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29830_ (.A1(_05715_),
    .A2(_05750_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29831_ (.A1(net18466),
    .A2(net18044),
    .B(net19554),
    .ZN(_05751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29832_ (.A1(_05751_),
    .A2(_05469_),
    .ZN(_05752_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29833_ (.A1(net18466),
    .A2(_05467_),
    .ZN(_05753_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29834_ (.A1(_05753_),
    .A2(net19554),
    .A3(_05606_),
    .ZN(_05754_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29835_ (.A1(_05752_),
    .A2(_05754_),
    .A3(net20183),
    .ZN(_05755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29836_ (.A1(_05569_),
    .A2(net17667),
    .ZN(_05756_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29837_ (.A1(_05481_),
    .A2(_05756_),
    .A3(net19560),
    .ZN(_05757_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29838_ (.A1(net17657),
    .A2(net19023),
    .B(net19559),
    .ZN(_05758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29839_ (.A1(_05518_),
    .A2(net18376),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29840_ (.A1(_05758_),
    .A2(_05511_),
    .A3(_05759_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29841_ (.A1(_05757_),
    .A2(_05760_),
    .A3(net19936),
    .ZN(_05761_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29842_ (.A1(_05755_),
    .A2(_05761_),
    .A3(net20397),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29843_ (.A1(_05593_),
    .A2(net18037),
    .A3(net19561),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29844_ (.A1(_05391_),
    .A2(_05363_),
    .ZN(_05764_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29845_ (.A1(_05764_),
    .A2(net19051),
    .ZN(_05765_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29846_ (.A1(net18467),
    .A2(net18047),
    .A3(net19033),
    .ZN(_05766_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29847_ (.A1(_05765_),
    .A2(_05766_),
    .A3(net19555),
    .ZN(_05767_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29848_ (.A1(_05763_),
    .A2(_05767_),
    .A3(net20183),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29849_ (.A1(_05421_),
    .A2(net19022),
    .A3(net19020),
    .ZN(_05769_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29850_ (.A1(_05589_),
    .A2(_05769_),
    .A3(net19561),
    .ZN(_05770_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _29851_ (.A1(net17664),
    .A2(net19559),
    .A3(net17663),
    .Z(_05771_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29852_ (.A1(_05770_),
    .A2(net19937),
    .A3(_05771_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29853_ (.A1(_05768_),
    .A2(_05514_),
    .A3(_05772_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29854_ (.A1(_05762_),
    .A2(_05773_),
    .A3(net19940),
    .ZN(_05774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29855_ (.A1(_05405_),
    .A2(net19559),
    .Z(_05775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29856_ (.A1(_05523_),
    .A2(net18043),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29857_ (.A1(_05775_),
    .A2(_05776_),
    .ZN(_05777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29858_ (.A1(_05571_),
    .A2(net19038),
    .ZN(_05778_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29859_ (.A1(_05778_),
    .A2(net19546),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29860_ (.A1(_05779_),
    .A2(net18038),
    .B(net20183),
    .ZN(_05780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29861_ (.A1(_05777_),
    .A2(_05780_),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29862_ (.A1(_05451_),
    .A2(net17674),
    .ZN(_05782_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29863_ (.A1(_05518_),
    .A2(net19546),
    .ZN(_05783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29864_ (.A1(_05782_),
    .A2(_05783_),
    .B(_05457_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29865_ (.A1(net18473),
    .A2(net19053),
    .A3(net18044),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29866_ (.A1(_05585_),
    .A2(_05785_),
    .A3(net19555),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29867_ (.A1(_05784_),
    .A2(_05786_),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29868_ (.A1(_05781_),
    .A2(net20179),
    .A3(_05787_),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29869_ (.A1(_05764_),
    .A2(net19027),
    .Z(_05789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29870_ (.A1(net17664),
    .A2(net19016),
    .ZN(_05790_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29871_ (.A1(_05789_),
    .A2(net19546),
    .A3(_05790_),
    .ZN(_05791_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29872_ (.A1(_05493_),
    .A2(_05455_),
    .A3(net19559),
    .ZN(_05792_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29873_ (.A1(_05791_),
    .A2(_05792_),
    .A3(net20182),
    .ZN(_05793_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29874_ (.I(_16119_[0]),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29875_ (.A1(_05794_),
    .A2(net19040),
    .B(net19546),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29876_ (.I(_05622_),
    .ZN(_05796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29877_ (.A1(_05795_),
    .A2(_05796_),
    .B(net20182),
    .ZN(_05797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29878_ (.A1(_05529_),
    .A2(net19015),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29879_ (.A1(_05798_),
    .A2(net19046),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29880_ (.A1(_05480_),
    .A2(_05529_),
    .ZN(_05800_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29881_ (.A1(_05799_),
    .A2(_05800_),
    .A3(net19554),
    .ZN(_05801_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29882_ (.A1(_05797_),
    .A2(_05801_),
    .B(_05514_),
    .ZN(_05802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29883_ (.A1(_05793_),
    .A2(_05802_),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29884_ (.A1(_05788_),
    .A2(net20181),
    .A3(_05803_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29885_ (.A1(_05774_),
    .A2(_05804_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29886_ (.A1(net19019),
    .A2(net19027),
    .B(net19546),
    .ZN(_05805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29887_ (.A1(_05789_),
    .A2(_05805_),
    .ZN(_05806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29888_ (.A1(_05806_),
    .A2(_05457_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _29889_ (.A1(_05705_),
    .A2(_05709_),
    .A3(net19027),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29890_ (.A1(net18054),
    .A2(_05544_),
    .B(net19546),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29891_ (.A1(_05808_),
    .A2(_05809_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29892_ (.A1(_05807_),
    .A2(_05810_),
    .ZN(_05811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29893_ (.I(_05394_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29894_ (.A1(_05778_),
    .A2(_05812_),
    .Z(_05813_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29895_ (.A1(_05813_),
    .A2(_05759_),
    .B(net19559),
    .ZN(_05814_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _29896_ (.A1(_05427_),
    .A2(_05492_),
    .B(net19559),
    .C(_05633_),
    .ZN(_05815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29897_ (.A1(_05815_),
    .A2(net20182),
    .ZN(_05816_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29898_ (.A1(_05814_),
    .A2(_05816_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29899_ (.A1(_05811_),
    .A2(_05817_),
    .B(net20397),
    .ZN(_05818_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29900_ (.A1(_05439_),
    .A2(net19547),
    .ZN(_05819_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29901_ (.A1(_05819_),
    .A2(_05736_),
    .B(_05457_),
    .ZN(_05820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29902_ (.A1(net18051),
    .A2(net19032),
    .B(_05523_),
    .ZN(_05821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29903_ (.A1(_05821_),
    .A2(net19547),
    .ZN(_05822_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29904_ (.A1(_05820_),
    .A2(_05822_),
    .B(net20397),
    .ZN(_05823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29905_ (.A1(net19028),
    .A2(net18373),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29906_ (.A1(_05467_),
    .A2(net17658),
    .ZN(_05825_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29907_ (.A1(_05486_),
    .A2(_05824_),
    .A3(_05825_),
    .ZN(_05826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29908_ (.A1(_05559_),
    .A2(net17676),
    .ZN(_05827_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29909_ (.A1(_05827_),
    .A2(net19562),
    .A3(_05408_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29910_ (.A1(_05826_),
    .A2(_05828_),
    .A3(net19935),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29911_ (.A1(_05823_),
    .A2(_05829_),
    .ZN(_05830_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29912_ (.A1(_05818_),
    .A2(net19940),
    .A3(_05830_),
    .ZN(_05831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29913_ (.A1(net19570),
    .A2(net19024),
    .B(net19546),
    .ZN(_05832_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29914_ (.A1(_05832_),
    .A2(_05453_),
    .B(net20182),
    .ZN(_05833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29915_ (.A1(_05428_),
    .A2(net18484),
    .ZN(_05834_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29916_ (.A1(_05620_),
    .A2(net18467),
    .ZN(_05835_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29917_ (.A1(_05834_),
    .A2(_05835_),
    .A3(net19552),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29918_ (.A1(_05833_),
    .A2(_05836_),
    .B(net20397),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29919_ (.A1(_05632_),
    .A2(net19042),
    .ZN(_05838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29920_ (.A1(_05775_),
    .A2(_05838_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29921_ (.A1(net18474),
    .A2(net19042),
    .A3(net17675),
    .ZN(_05840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29922_ (.A1(net17656),
    .A2(net19037),
    .B(net19559),
    .ZN(_05841_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29923_ (.A1(_05840_),
    .A2(_05841_),
    .B(_05457_),
    .ZN(_05842_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29924_ (.A1(_05839_),
    .A2(_05842_),
    .ZN(_05843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29925_ (.A1(_05837_),
    .A2(_05843_),
    .ZN(_05844_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29926_ (.A1(net18045),
    .A2(net19028),
    .B(net19548),
    .ZN(_05845_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29927_ (.A1(net18474),
    .A2(net19042),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29928_ (.A1(_05845_),
    .A2(_05846_),
    .B(_05457_),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29929_ (.A1(_05689_),
    .A2(_05371_),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29930_ (.A1(_05428_),
    .A2(net17387),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29931_ (.A1(_05848_),
    .A2(_05849_),
    .A3(net19554),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29932_ (.A1(_05847_),
    .A2(_05850_),
    .B(_05514_),
    .ZN(_05851_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29933_ (.A1(net18051),
    .A2(_05561_),
    .B(net19043),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29934_ (.I(net17236),
    .ZN(_05853_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29935_ (.A1(_05852_),
    .A2(net19563),
    .A3(_05853_),
    .ZN(_05854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29936_ (.A1(_05531_),
    .A2(net17384),
    .B(net20183),
    .ZN(_05855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29937_ (.A1(_05854_),
    .A2(_05855_),
    .ZN(_05856_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29938_ (.A1(_05851_),
    .A2(_05856_),
    .ZN(_05857_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29939_ (.A1(_05844_),
    .A2(_05857_),
    .A3(net20181),
    .ZN(_05858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29940_ (.A1(_05831_),
    .A2(_05858_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29941_ (.A1(_05467_),
    .A2(net19022),
    .A3(net18478),
    .ZN(_05859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29942_ (.A1(_05472_),
    .A2(net17382),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29943_ (.A1(_05859_),
    .A2(net19559),
    .A3(_05860_),
    .ZN(_05861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29944_ (.A1(net17656),
    .A2(net19042),
    .B(net19559),
    .ZN(_05862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29945_ (.A1(net19015),
    .A2(net19060),
    .ZN(_05863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29946_ (.A1(_05863_),
    .A2(net19037),
    .ZN(_05864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29947_ (.A1(_05862_),
    .A2(_05864_),
    .B(_05514_),
    .ZN(_05865_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29948_ (.A1(_05861_),
    .A2(_05865_),
    .B(net19932),
    .ZN(_05866_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29949_ (.A1(_05620_),
    .A2(net17668),
    .B(net19546),
    .ZN(_05867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29950_ (.A1(_05660_),
    .A2(net19031),
    .ZN(_05868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29951_ (.A1(_05867_),
    .A2(net17388),
    .A3(_05868_),
    .ZN(_05869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29952_ (.A1(_05451_),
    .A2(net18043),
    .ZN(_05870_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29953_ (.A1(net19567),
    .A2(net17655),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29954_ (.A1(net17657),
    .A2(_05871_),
    .B(net19036),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29955_ (.A1(_05870_),
    .A2(_05872_),
    .A3(net19546),
    .ZN(_05873_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29956_ (.A1(_05869_),
    .A2(_05514_),
    .A3(_05873_),
    .ZN(_05874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29957_ (.A1(_05866_),
    .A2(_05874_),
    .B(net20180),
    .ZN(_05875_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29958_ (.A1(_05393_),
    .A2(_05812_),
    .ZN(_05876_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29959_ (.A1(_05876_),
    .A2(net19042),
    .B(_05778_),
    .ZN(_05877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29960_ (.A1(_05551_),
    .A2(net19041),
    .B(net19546),
    .ZN(_05878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29961_ (.A1(_05877_),
    .A2(_05878_),
    .ZN(_05879_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29962_ (.A1(_05720_),
    .A2(net19546),
    .Z(_05880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29963_ (.A1(_05670_),
    .A2(_05880_),
    .B(_05514_),
    .ZN(_05881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29964_ (.A1(_05881_),
    .A2(_05879_),
    .ZN(_05882_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29965_ (.A1(_05464_),
    .A2(net18041),
    .B(net19054),
    .ZN(_05883_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29966_ (.A1(_05540_),
    .A2(net19054),
    .Z(_05884_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _29967_ (.A1(_05883_),
    .A2(net19559),
    .A3(_05884_),
    .ZN(_05885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29968_ (.A1(_05646_),
    .A2(_05363_),
    .ZN(_05886_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _29969_ (.A1(_16124_[0]),
    .A2(_16133_[0]),
    .Z(_05887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29970_ (.A1(net19054),
    .A2(_05887_),
    .B(net19546),
    .ZN(_05888_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29971_ (.A1(_05886_),
    .A2(_05888_),
    .Z(_05889_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29972_ (.A1(_05885_),
    .A2(_05889_),
    .B(_05514_),
    .ZN(_05890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29973_ (.A1(_05882_),
    .A2(_05890_),
    .ZN(_05891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29974_ (.A1(_05891_),
    .A2(_05457_),
    .ZN(_05892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29975_ (.A1(_05875_),
    .A2(_05892_),
    .ZN(_05893_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _29976_ (.A1(_05452_),
    .A2(net19027),
    .Z(_05894_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29977_ (.A1(_05894_),
    .A2(_05569_),
    .B(net18479),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29978_ (.A1(_05895_),
    .A2(net19553),
    .ZN(_05896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29979_ (.A1(net19051),
    .A2(net19019),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29980_ (.A1(_05699_),
    .A2(_05897_),
    .B(net20182),
    .ZN(_05898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29981_ (.A1(_05896_),
    .A2(_05898_),
    .ZN(_05899_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29982_ (.A1(_05736_),
    .A2(_05878_),
    .B(_05457_),
    .ZN(_05900_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29983_ (.A1(_05364_),
    .A2(net19555),
    .A3(net18039),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29984_ (.A1(_05900_),
    .A2(_05901_),
    .ZN(_05902_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29985_ (.A1(_05899_),
    .A2(_05902_),
    .A3(net20179),
    .ZN(_05903_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _29986_ (.A1(net17660),
    .A2(net17384),
    .B(_05582_),
    .ZN(_05904_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _29987_ (.I(_16125_[0]),
    .ZN(_05905_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29988_ (.A1(_05905_),
    .A2(net19023),
    .B(net19546),
    .ZN(_05906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29989_ (.A1(_05906_),
    .A2(_05835_),
    .B(net20182),
    .ZN(_05907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29990_ (.A1(_05904_),
    .A2(_05907_),
    .ZN(_05908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29991_ (.A1(_05604_),
    .A2(net19560),
    .ZN(_05909_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _29992_ (.A1(net17389),
    .A2(net19559),
    .ZN(_05910_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _29993_ (.A1(_05910_),
    .A2(_05800_),
    .B(_05457_),
    .ZN(_05911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29994_ (.A1(_05909_),
    .A2(_05911_),
    .ZN(_05912_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29995_ (.A1(_05908_),
    .A2(_05912_),
    .A3(net20397),
    .ZN(_05913_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _29996_ (.A1(_05903_),
    .A2(_05913_),
    .A3(net20181),
    .ZN(_05914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29997_ (.A1(_05893_),
    .A2(_05914_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _29998_ (.A1(_05440_),
    .A2(_05434_),
    .Z(_05915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _29999_ (.A1(_05915_),
    .A2(net19040),
    .ZN(_05916_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _30000_ (.A1(_05551_),
    .A2(net19040),
    .A3(net17666),
    .Z(_05917_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30001_ (.A1(_05916_),
    .A2(net19559),
    .A3(_05917_),
    .ZN(_05918_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30002_ (.A1(_05735_),
    .A2(net19017),
    .B(net19040),
    .ZN(_05919_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30003_ (.A1(_05919_),
    .A2(net19556),
    .A3(_05743_),
    .ZN(_05920_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30004_ (.A1(_05918_),
    .A2(_05920_),
    .A3(net19939),
    .ZN(_05921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30005_ (.A1(_05528_),
    .A2(_05778_),
    .ZN(_05922_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _30006_ (.A1(_05922_),
    .A2(net19559),
    .A3(_05434_),
    .Z(_05923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30007_ (.A1(net19040),
    .A2(net18373),
    .ZN(_05924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30008_ (.A1(_05886_),
    .A2(_05924_),
    .B(net19559),
    .ZN(_05925_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30009_ (.A1(_05923_),
    .A2(_05925_),
    .B(net20182),
    .ZN(_05926_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30010_ (.A1(_05921_),
    .A2(_05926_),
    .A3(_05514_),
    .ZN(_05927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30011_ (.A1(_05794_),
    .A2(net19028),
    .B(net19556),
    .ZN(_05928_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30012_ (.A1(_05928_),
    .A2(_05465_),
    .B(net20182),
    .ZN(_05929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30013_ (.A1(_05863_),
    .A2(net19040),
    .ZN(_05930_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30014_ (.A1(_05585_),
    .A2(net19549),
    .A3(_05930_),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30015_ (.A1(_05929_),
    .A2(_05931_),
    .B(_05514_),
    .ZN(_05932_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30016_ (.A1(_05425_),
    .A2(net18048),
    .ZN(_05933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30017_ (.A1(_05574_),
    .A2(net18467),
    .ZN(_05934_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30018_ (.A1(_05933_),
    .A2(_05934_),
    .A3(net19551),
    .ZN(_05935_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30019_ (.A1(net17383),
    .A2(net17657),
    .B(net19045),
    .ZN(_05936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30020_ (.A1(net18370),
    .A2(net19024),
    .B(net19546),
    .ZN(_05937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30021_ (.A1(_05936_),
    .A2(_05937_),
    .B(_05457_),
    .ZN(_05938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30022_ (.A1(_05935_),
    .A2(_05938_),
    .ZN(_05939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30023_ (.A1(_05932_),
    .A2(_05939_),
    .B(net20180),
    .ZN(_05940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30024_ (.A1(_05927_),
    .A2(_05940_),
    .ZN(_05941_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30025_ (.I(_05799_),
    .ZN(_05942_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30026_ (.A1(_05942_),
    .A2(_05581_),
    .ZN(_05943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30027_ (.A1(_05915_),
    .A2(net19031),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30028_ (.A1(_05943_),
    .A2(_05944_),
    .ZN(_05945_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30029_ (.A1(_05569_),
    .A2(net19547),
    .ZN(_05946_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30030_ (.A1(_05946_),
    .A2(_05800_),
    .B(net20397),
    .ZN(_05947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30031_ (.A1(_05945_),
    .A2(_05947_),
    .B(net20183),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30032_ (.A1(net18036),
    .A2(net19053),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30033_ (.A1(_05654_),
    .A2(_05765_),
    .A3(_05949_),
    .ZN(_05950_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30034_ (.A1(net19051),
    .A2(net19566),
    .ZN(_05951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30035_ (.A1(_05769_),
    .A2(_05951_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30036_ (.A1(_05952_),
    .A2(net19555),
    .B(_05514_),
    .ZN(_05953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30037_ (.A1(_05950_),
    .A2(_05953_),
    .ZN(_05954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30038_ (.A1(_05948_),
    .A2(_05954_),
    .ZN(_05955_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30039_ (.A1(_05720_),
    .A2(net19559),
    .Z(_05956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30040_ (.A1(_05561_),
    .A2(net19032),
    .ZN(_05957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30041_ (.A1(_05956_),
    .A2(_05957_),
    .B(_05514_),
    .ZN(_05958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30042_ (.A1(_05467_),
    .A2(net19032),
    .ZN(_05959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30043_ (.A1(_05689_),
    .A2(net18472),
    .ZN(_05960_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30044_ (.A1(_05959_),
    .A2(_05960_),
    .A3(net19547),
    .ZN(_05961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30045_ (.A1(_05958_),
    .A2(_05961_),
    .B(_05457_),
    .ZN(_05962_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30046_ (.A1(_05533_),
    .A2(_05724_),
    .A3(net19549),
    .ZN(_05963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30047_ (.A1(_05867_),
    .A2(_05647_),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30048_ (.A1(_05963_),
    .A2(_05964_),
    .A3(_05514_),
    .ZN(_05965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30049_ (.A1(_05962_),
    .A2(_05965_),
    .ZN(_05966_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30050_ (.A1(_05955_),
    .A2(_05966_),
    .A3(net20180),
    .ZN(_05967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30051_ (.A1(_05941_),
    .A2(_05967_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30052_ (.A1(_03026_),
    .A2(_03018_),
    .ZN(_05968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30053_ (.A1(_12024_),
    .A2(_03022_),
    .ZN(_05969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30054_ (.A1(_05968_),
    .A2(_05969_),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30055_ (.I(_05970_),
    .ZN(_05971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30056_ (.A1(_11973_),
    .A2(net21343),
    .ZN(_05972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30057_ (.A1(_11969_),
    .A2(net21032),
    .ZN(_05973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30058_ (.A1(_05973_),
    .A2(_05972_),
    .ZN(_05974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30059_ (.A1(_05971_),
    .A2(net20627),
    .ZN(_05975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30060_ (.I(_05974_),
    .ZN(_05976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30061_ (.A1(_05976_),
    .A2(net20628),
    .ZN(_05977_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30062_ (.A1(_05977_),
    .A2(_05975_),
    .A3(_10378_),
    .ZN(_05978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30063_ (.I(net21172),
    .ZN(_05979_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _30064_ (.A1(_10378_),
    .A2(\text_in_r[33] ),
    .Z(_05980_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30065_ (.A1(_05979_),
    .A2(_05978_),
    .A3(_05980_),
    .ZN(_05981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30066_ (.A1(_05976_),
    .A2(_05971_),
    .ZN(_05982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30067_ (.A1(_05970_),
    .A2(net20627),
    .ZN(_05983_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30068_ (.A1(_05983_),
    .A2(_10378_),
    .A3(_05982_),
    .ZN(_05984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30069_ (.A1(net21508),
    .A2(\text_in_r[33] ),
    .ZN(_05985_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30070_ (.A1(_05985_),
    .A2(net21172),
    .A3(_05984_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30071_ (.A1(_05986_),
    .A2(_05981_),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input94 (.I(key[69]),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30073_ (.A1(_12005_),
    .A2(_12007_),
    .A3(net21275),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30074_ (.A1(net21024),
    .A2(net21021),
    .ZN(_05989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30075_ (.A1(net21398),
    .A2(net21345),
    .ZN(_05990_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30076_ (.A1(_05989_),
    .A2(net20967),
    .A3(_05990_),
    .ZN(_05991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30077_ (.A1(_05988_),
    .A2(_05991_),
    .ZN(_05992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30078_ (.A1(_05992_),
    .A2(net20901),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30079_ (.A1(_05988_),
    .A2(_05991_),
    .A3(net20902),
    .ZN(_05994_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30080_ (.A1(_05993_),
    .A2(_05994_),
    .B(net21501),
    .ZN(_05995_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30081_ (.I(\text_in_r[32] ),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30082_ (.A1(_05996_),
    .A2(net21501),
    .Z(_05997_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30083_ (.A1(net20396),
    .A2(_05997_),
    .B(net21181),
    .ZN(_05998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30084_ (.A1(_05993_),
    .A2(_05994_),
    .ZN(_05999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30085_ (.A1(_05999_),
    .A2(net21083),
    .ZN(_06000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30086_ (.I(net21181),
    .ZN(_06001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30087_ (.I(_05997_),
    .ZN(_06002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30088_ (.A1(net20178),
    .A2(_06001_),
    .A3(_06002_),
    .ZN(_06003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30089_ (.A1(_05998_),
    .A2(_06003_),
    .ZN(_16146_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30090_ (.A1(net21283),
    .A2(\sa20_sub[2] ),
    .Z(_06004_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30091_ (.A1(net21283),
    .A2(net21340),
    .ZN(_06005_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30092_ (.A1(_06004_),
    .A2(_06005_),
    .B(net21452),
    .ZN(_06006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30093_ (.A1(net21031),
    .A2(_12025_),
    .ZN(_06007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30094_ (.A1(net21283),
    .A2(\sa20_sub[2] ),
    .ZN(_06008_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30095_ (.A1(_06007_),
    .A2(_12057_),
    .A3(_06008_),
    .ZN(_06009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30096_ (.A1(_06006_),
    .A2(_06009_),
    .ZN(_06010_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _30097_ (.A1(net21453),
    .A2(\sa12_sr[2] ),
    .ZN(_06011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30098_ (.I(_06011_),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30099_ (.A1(_06010_),
    .A2(_06012_),
    .ZN(_06013_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30100_ (.A1(_06006_),
    .A2(_06009_),
    .A3(_06011_),
    .ZN(_06014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30101_ (.A1(_06013_),
    .A2(_06014_),
    .B(net21501),
    .ZN(_06015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30102_ (.I(\text_in_r[34] ),
    .ZN(_06016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30103_ (.A1(_06016_),
    .A2(net21508),
    .Z(_06017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30104_ (.I(net21163),
    .ZN(_06018_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30105_ (.A1(_06015_),
    .A2(_06017_),
    .B(_06018_),
    .ZN(_06019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30106_ (.A1(_06013_),
    .A2(_06014_),
    .ZN(_06020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30107_ (.A1(_06020_),
    .A2(net21083),
    .ZN(_06021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30108_ (.I(_06017_),
    .ZN(_06022_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30109_ (.A1(_06021_),
    .A2(net21163),
    .A3(_06022_),
    .ZN(_06023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30110_ (.A1(_06023_),
    .A2(_06019_),
    .ZN(_06024_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input93 (.I(key[68]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input92 (.I(key[67]),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30113_ (.A1(_05995_),
    .A2(_05997_),
    .B(_06001_),
    .ZN(_06026_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30114_ (.A1(_06000_),
    .A2(net21181),
    .A3(_06002_),
    .ZN(_06027_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30115_ (.A1(_06026_),
    .A2(_06027_),
    .ZN(_16137_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30116_ (.A1(_06015_),
    .A2(net20926),
    .B(net21163),
    .ZN(_06028_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30117_ (.A1(_06021_),
    .A2(_06018_),
    .A3(_06022_),
    .ZN(_06029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30118_ (.A1(_06028_),
    .A2(_06029_),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input91 (.I(key[66]),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input90 (.I(key[65]),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30121_ (.A1(_06024_),
    .A2(net19534),
    .ZN(_06032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30122_ (.A1(_12064_),
    .A2(net21338),
    .ZN(_06033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30123_ (.A1(_12060_),
    .A2(net21015),
    .ZN(_06034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30124_ (.A1(_06033_),
    .A2(_06034_),
    .ZN(_06035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30125_ (.A1(_03108_),
    .A2(_06035_),
    .ZN(_06036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30126_ (.A1(_12060_),
    .A2(net21338),
    .ZN(_06037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30127_ (.A1(_12064_),
    .A2(net21015),
    .ZN(_06038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30128_ (.A1(_06037_),
    .A2(_06038_),
    .ZN(_06039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30129_ (.A1(_03116_),
    .A2(_06039_),
    .ZN(_06040_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30130_ (.A1(_06036_),
    .A2(_06040_),
    .A3(net21088),
    .ZN(_06041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30131_ (.I(net21160),
    .ZN(_06042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30132_ (.A1(net21508),
    .A2(\text_in_r[35] ),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30133_ (.A1(_06041_),
    .A2(_06042_),
    .A3(_06043_),
    .ZN(_06044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30134_ (.A1(_03108_),
    .A2(_06039_),
    .ZN(_06045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30135_ (.A1(_03116_),
    .A2(_06035_),
    .ZN(_06046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30136_ (.A1(_06045_),
    .A2(_06046_),
    .A3(net21088),
    .ZN(_06047_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _30137_ (.A1(net21081),
    .A2(\text_in_r[35] ),
    .Z(_06048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30138_ (.A1(_06047_),
    .A2(net21160),
    .A3(_06048_),
    .ZN(_06049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30139_ (.A1(_06044_),
    .A2(_06049_),
    .ZN(_06050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30140_ (.A1(_06032_),
    .A2(net19515),
    .Z(_06051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30141_ (.I(_16144_[0]),
    .ZN(_06052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30142_ (.A1(net20177),
    .A2(_06052_),
    .A3(net19931),
    .ZN(_06053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30143_ (.A1(_06047_),
    .A2(_06042_),
    .A3(_06048_),
    .ZN(_06054_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30144_ (.A1(_06041_),
    .A2(net21160),
    .A3(_06043_),
    .ZN(_06055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30145_ (.A1(_06054_),
    .A2(_06055_),
    .ZN(_06056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30146_ (.A1(_06053_),
    .A2(net19503),
    .ZN(_06057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30147_ (.I(_06057_),
    .ZN(_06058_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30148_ (.A1(_05978_),
    .A2(net21172),
    .A3(_05980_),
    .ZN(_06059_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30149_ (.A1(_05979_),
    .A2(_05984_),
    .A3(_05985_),
    .ZN(_06060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30150_ (.A1(_06059_),
    .A2(_06060_),
    .ZN(_16138_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _30151_ (.A1(_06032_),
    .A2(net19010),
    .Z(_06061_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30152_ (.A1(net18465),
    .A2(_06058_),
    .B(_06061_),
    .ZN(_06062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30153_ (.A1(_03130_),
    .A2(_12112_),
    .ZN(_06063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30154_ (.A1(_12109_),
    .A2(_03135_),
    .ZN(_06064_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30155_ (.A1(_06063_),
    .A2(_06064_),
    .A3(net21081),
    .ZN(_06065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30156_ (.A1(net21508),
    .A2(\text_in_r[36] ),
    .ZN(_06066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30157_ (.A1(_06065_),
    .A2(_06066_),
    .ZN(_06067_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30158_ (.A1(_06067_),
    .A2(net21159),
    .ZN(_06068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30159_ (.I(net21159),
    .ZN(_06069_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30160_ (.A1(_06065_),
    .A2(_06069_),
    .A3(_06066_),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30161_ (.A1(_06068_),
    .A2(_06070_),
    .ZN(_06071_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input89 (.I(key[64]),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input88 (.I(net551),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30164_ (.A1(_06062_),
    .A2(net19491),
    .ZN(_06074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30165_ (.A1(net19530),
    .A2(net19534),
    .ZN(_06075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input87 (.I(net586),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30167_ (.A1(_06075_),
    .A2(net19515),
    .Z(_06077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30168_ (.A1(_06061_),
    .A2(_06077_),
    .ZN(_06078_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30169_ (.I(_16153_[0]),
    .ZN(_06079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30170_ (.A1(net19541),
    .A2(_06079_),
    .ZN(_06080_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input86 (.I(key[61]),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30172_ (.A1(_06080_),
    .A2(net19510),
    .ZN(_06082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30173_ (.I(_06082_),
    .ZN(_06083_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30174_ (.I(_16140_[0]),
    .ZN(_06084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30175_ (.A1(net19530),
    .A2(_06084_),
    .ZN(_06085_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input85 (.I(net541),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30177_ (.A1(_06083_),
    .A2(net17651),
    .ZN(_06087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30178_ (.A1(_06067_),
    .A2(_06069_),
    .ZN(_06088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30179_ (.A1(_06065_),
    .A2(net21159),
    .A3(_06066_),
    .ZN(_06089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30180_ (.A1(_06088_),
    .A2(_06089_),
    .ZN(_06090_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input84 (.I(key[5]),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input83 (.I(net549),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30183_ (.A1(_06078_),
    .A2(_06087_),
    .A3(net19480),
    .ZN(_06093_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30184_ (.A1(net21278),
    .A2(net21336),
    .Z(_06094_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30185_ (.A1(_06094_),
    .A2(_15180_),
    .Z(_06095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30186_ (.A1(_06094_),
    .A2(_15180_),
    .ZN(_06096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30187_ (.A1(_06095_),
    .A2(_06096_),
    .ZN(_06097_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _30188_ (.A1(net21448),
    .A2(\sa12_sr[5] ),
    .ZN(_06098_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30189_ (.I(_06098_),
    .ZN(_06099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30190_ (.A1(_06097_),
    .A2(_06099_),
    .ZN(_06100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30191_ (.A1(_06095_),
    .A2(_06098_),
    .A3(_06096_),
    .ZN(_06101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30192_ (.A1(_06100_),
    .A2(_06101_),
    .A3(net21081),
    .ZN(_06102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30193_ (.A1(net21508),
    .A2(\text_in_r[37] ),
    .ZN(_06103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30194_ (.A1(_06102_),
    .A2(_06103_),
    .ZN(_06104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30195_ (.A1(_06104_),
    .A2(net21158),
    .ZN(_06105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30196_ (.I(net21158),
    .ZN(_06106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30197_ (.A1(_06102_),
    .A2(_06106_),
    .A3(_06103_),
    .ZN(_06107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30198_ (.A1(_06105_),
    .A2(_06107_),
    .ZN(_06108_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _30199_ (.I(_06108_),
    .ZN(_06109_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input82 (.I(key[58]),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30201_ (.A1(_06074_),
    .A2(_06093_),
    .A3(net19470),
    .ZN(_06111_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input81 (.I(net545),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30203_ (.A1(net19010),
    .A2(net19531),
    .B(net19497),
    .ZN(_06113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30204_ (.A1(_06113_),
    .A2(_06061_),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30205_ (.A1(_06032_),
    .A2(net19497),
    .Z(_06115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30206_ (.A1(_06079_),
    .A2(net19530),
    .ZN(_06116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30207_ (.A1(_06115_),
    .A2(net17647),
    .ZN(_06117_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input80 (.I(net547),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30209_ (.A1(_06114_),
    .A2(_06117_),
    .A3(net19485),
    .ZN(_06119_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30210_ (.A1(net19014),
    .A2(net19544),
    .A3(net19530),
    .ZN(_06120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30211_ (.A1(_06115_),
    .A2(_06120_),
    .ZN(_06121_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30212_ (.I(_16141_[0]),
    .ZN(_06122_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _30213_ (.A1(_06122_),
    .A2(net19535),
    .ZN(_06123_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input79 (.I(net582),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _30215_ (.A1(_06123_),
    .A2(net19516),
    .B(net19483),
    .ZN(_06125_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _30216_ (.A1(net19013),
    .A2(net19532),
    .ZN(_06126_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input78 (.I(net572),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30218_ (.A1(_06126_),
    .A2(net19520),
    .ZN(_06128_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30219_ (.A1(_06121_),
    .A2(_06125_),
    .A3(_06128_),
    .ZN(_06129_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input77 (.I(net568),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30221_ (.A1(_06119_),
    .A2(_06129_),
    .A3(net19928),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _30222_ (.A1(net21277),
    .A2(\sa20_sub[6] ),
    .A3(net21447),
    .Z(_06132_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30223_ (.A1(\sa02_sr[5] ),
    .A2(net21388),
    .Z(_06133_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30224_ (.A1(_06132_),
    .A2(_06133_),
    .Z(_06134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30225_ (.A1(_06132_),
    .A2(_06133_),
    .ZN(_06135_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30226_ (.A1(_06134_),
    .A2(net21081),
    .A3(_06135_),
    .ZN(_06136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30227_ (.A1(net21507),
    .A2(\text_in_r[38] ),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30228_ (.A1(_06136_),
    .A2(_06137_),
    .ZN(_06138_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30229_ (.I(\u0.w[2][6] ),
    .ZN(_06139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30230_ (.A1(_06138_),
    .A2(_06139_),
    .ZN(_06140_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30231_ (.A1(_06136_),
    .A2(\u0.w[2][6] ),
    .A3(_06137_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30232_ (.A1(_06140_),
    .A2(_06141_),
    .ZN(_06142_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input76 (.I(key[52]),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30234_ (.A1(_06111_),
    .A2(_06131_),
    .A3(net20395),
    .ZN(_06144_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30235_ (.I(_16139_[0]),
    .ZN(_06145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30236_ (.A1(net19538),
    .A2(_06145_),
    .ZN(_06146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30237_ (.I(_06146_),
    .ZN(_06147_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30238_ (.I(_16147_[0]),
    .ZN(_06148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30239_ (.A1(net19531),
    .A2(_06148_),
    .ZN(_06149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30240_ (.I(_06149_),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input75 (.I(key[51]),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30242_ (.A1(_06147_),
    .A2(_06150_),
    .B(net19507),
    .ZN(_06152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30243_ (.A1(net490),
    .A2(net19515),
    .Z(_06153_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30244_ (.A1(net19014),
    .A2(net19544),
    .A3(net19541),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30245_ (.A1(_06153_),
    .A2(_06154_),
    .ZN(_06155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30246_ (.A1(_06152_),
    .A2(_06155_),
    .A3(net19495),
    .ZN(_06156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30247_ (.A1(net19530),
    .A2(net19543),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30248_ (.A1(_06157_),
    .A2(net19515),
    .Z(_06158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30249_ (.A1(net19010),
    .A2(net19534),
    .ZN(_06159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30250_ (.A1(_06158_),
    .A2(_06159_),
    .ZN(_06160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30251_ (.A1(net19014),
    .A2(net19534),
    .ZN(_06161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30252_ (.A1(net19541),
    .A2(net19543),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30253_ (.A1(_06161_),
    .A2(net19505),
    .A3(_06162_),
    .ZN(_06163_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30254_ (.A1(_06160_),
    .A2(_06163_),
    .A3(net19481),
    .ZN(_06164_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30255_ (.A1(_06156_),
    .A2(_06164_),
    .A3(net19468),
    .ZN(_06165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30256_ (.A1(net19013),
    .A2(net19538),
    .ZN(_06166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30257_ (.A1(net19530),
    .A2(net18368),
    .ZN(_06167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30258_ (.A1(_06166_),
    .A2(net18033),
    .ZN(_06168_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input74 (.I(net584),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30260_ (.A1(_06168_),
    .A2(net19523),
    .ZN(_06170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30261_ (.A1(_06084_),
    .A2(net19540),
    .ZN(_06171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30262_ (.I(_06171_),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30263_ (.A1(_06172_),
    .A2(net19512),
    .Z(_06173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30264_ (.I(_06173_),
    .ZN(_06174_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30265_ (.A1(_06170_),
    .A2(_06174_),
    .A3(net19480),
    .ZN(_06175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30266_ (.A1(net19532),
    .A2(_06145_),
    .ZN(_06176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30267_ (.A1(net19538),
    .A2(_06148_),
    .ZN(_06177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30268_ (.A1(net17645),
    .A2(net17643),
    .ZN(_06178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30269_ (.A1(_06178_),
    .A2(net19524),
    .ZN(_06179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30270_ (.A1(net19537),
    .A2(net18369),
    .ZN(_06180_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input73 (.I(key[4]),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30272_ (.A1(net17651),
    .A2(_06180_),
    .A3(net19511),
    .ZN(_06182_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input72 (.I(net587),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30274_ (.A1(_06179_),
    .A2(_06182_),
    .A3(net19490),
    .ZN(_06184_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input71 (.I(net569),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30276_ (.A1(_06175_),
    .A2(_06184_),
    .A3(net19928),
    .ZN(_06186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _30277_ (.I(_06142_),
    .ZN(_06187_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input70 (.I(net542),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30279_ (.A1(_06165_),
    .A2(_06186_),
    .A3(_06187_),
    .ZN(_06189_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30280_ (.A1(net21276),
    .A2(net20900),
    .Z(_06190_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _30281_ (.A1(_15233_),
    .A2(net21332),
    .A3(_06190_),
    .Z(_06191_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30282_ (.A1(net21507),
    .A2(\text_in_r[39] ),
    .Z(_06192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30283_ (.A1(_06191_),
    .A2(net21081),
    .B(_06192_),
    .ZN(_06193_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30284_ (.A1(\u0.w[2][7] ),
    .A2(_06193_),
    .Z(_06194_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input69 (.I(net550),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30286_ (.A1(_06144_),
    .A2(_06189_),
    .A3(net20175),
    .ZN(_06196_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30287_ (.A1(net19538),
    .A2(net18366),
    .ZN(_06197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30288_ (.A1(_06157_),
    .A2(_06197_),
    .ZN(_06198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30289_ (.A1(net19530),
    .A2(net19010),
    .ZN(_06199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30290_ (.I(_06199_),
    .ZN(_06200_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30291_ (.A1(_06198_),
    .A2(_06200_),
    .B(net19521),
    .ZN(_06201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30292_ (.A1(net19536),
    .A2(net18367),
    .ZN(_06202_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30293_ (.I(_06202_),
    .ZN(_06203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30294_ (.A1(_06203_),
    .A2(net19515),
    .ZN(_06204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30295_ (.A1(_06162_),
    .A2(_06176_),
    .ZN(_06205_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input68 (.I(key[45]),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30297_ (.A1(_06205_),
    .A2(net19505),
    .ZN(_06207_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30298_ (.A1(_06201_),
    .A2(net17377),
    .A3(_06207_),
    .ZN(_06208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30299_ (.A1(net19540),
    .A2(net18368),
    .ZN(_06209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30300_ (.A1(_06209_),
    .A2(net19515),
    .Z(_06210_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input67 (.I(net570),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30302_ (.A1(net19515),
    .A2(_16160_[0]),
    .ZN(_06212_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30303_ (.A1(_06210_),
    .A2(_06212_),
    .Z(_06213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30304_ (.A1(_06213_),
    .A2(net19482),
    .ZN(_06214_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30305_ (.A1(_06208_),
    .A2(net19480),
    .B(net19928),
    .C(_06214_),
    .ZN(_06215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30306_ (.A1(net19535),
    .A2(_16147_[0]),
    .ZN(_06216_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30307_ (.A1(_06216_),
    .A2(net19515),
    .Z(_06217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30308_ (.A1(net19013),
    .A2(net19534),
    .A3(net19532),
    .ZN(_06218_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30309_ (.A1(_06217_),
    .A2(_06218_),
    .Z(_06219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30310_ (.A1(_06123_),
    .A2(net19512),
    .ZN(_06220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30311_ (.A1(_06220_),
    .A2(net19476),
    .ZN(_06221_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30312_ (.A1(_06219_),
    .A2(_06221_),
    .Z(_06222_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30313_ (.I(_16149_[0]),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30314_ (.A1(net19540),
    .A2(_06223_),
    .ZN(_06224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30315_ (.A1(_06224_),
    .A2(net19514),
    .Z(_06225_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30316_ (.A1(_06225_),
    .A2(_06218_),
    .ZN(_06226_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input66 (.I(net580),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30318_ (.A1(_06226_),
    .A2(_06125_),
    .B(net19930),
    .ZN(_06228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30319_ (.A1(_06222_),
    .A2(_06228_),
    .B(net20395),
    .ZN(_06229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30320_ (.A1(_06215_),
    .A2(_06229_),
    .ZN(_06230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30321_ (.A1(_06085_),
    .A2(net19510),
    .ZN(_06231_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input65 (.I(key[42]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30323_ (.A1(_06231_),
    .A2(net19476),
    .Z(_06233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30324_ (.A1(net19530),
    .A2(net18365),
    .ZN(_06234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30325_ (.A1(_06197_),
    .A2(_06234_),
    .ZN(_06235_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30326_ (.A1(_06235_),
    .A2(net19515),
    .ZN(_06236_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input64 (.I(net576),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30328_ (.A1(_06233_),
    .A2(_06236_),
    .B(_06109_),
    .ZN(_06238_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30329_ (.I(_06197_),
    .ZN(_06239_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input63 (.I(key[40]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30331_ (.A1(_06239_),
    .A2(net19522),
    .ZN(_06241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30332_ (.A1(_06121_),
    .A2(net19489),
    .A3(_06241_),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input62 (.I(key[3]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30334_ (.A1(_06238_),
    .A2(_06242_),
    .B(_06187_),
    .ZN(_06244_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input61 (.I(key[39]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30336_ (.A1(_06147_),
    .A2(net489),
    .B(net19522),
    .ZN(_06246_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input60 (.I(key[38]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30338_ (.A1(_06246_),
    .A2(net19479),
    .A3(net17381),
    .ZN(_06248_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30339_ (.A1(net19014),
    .A2(net19530),
    .ZN(_06249_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30340_ (.A1(_06249_),
    .A2(net19529),
    .A3(net18028),
    .ZN(_06250_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30341_ (.A1(net19007),
    .A2(net18027),
    .A3(net19513),
    .ZN(_06251_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30342_ (.A1(_06250_),
    .A2(_06251_),
    .A3(net19492),
    .ZN(_06252_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input59 (.I(key[37]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30344_ (.A1(_06248_),
    .A2(_06252_),
    .A3(net19471),
    .ZN(_06254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30345_ (.A1(_06244_),
    .A2(_06254_),
    .B(_06194_),
    .ZN(_06255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30346_ (.A1(_06230_),
    .A2(_06255_),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30347_ (.A1(_06196_),
    .A2(_06256_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30348_ (.I(_06085_),
    .ZN(_06257_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input58 (.I(key[36]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30350_ (.A1(net17374),
    .A2(_06239_),
    .B(net19506),
    .ZN(_06259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30351_ (.A1(net17376),
    .A2(net19528),
    .ZN(_06260_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30352_ (.A1(_06259_),
    .A2(net19481),
    .A3(_06260_),
    .ZN(_06261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30353_ (.A1(net19014),
    .A2(net19544),
    .ZN(_06262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30354_ (.A1(_06262_),
    .A2(_06075_),
    .ZN(_06263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30355_ (.A1(_06263_),
    .A2(net19505),
    .ZN(_06264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30356_ (.A1(_06075_),
    .A2(net18029),
    .A3(net19515),
    .ZN(_06265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30357_ (.A1(_06264_),
    .A2(net19495),
    .A3(_06265_),
    .ZN(_06266_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30358_ (.A1(_06261_),
    .A2(_06266_),
    .A3(net19928),
    .ZN(_06267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30359_ (.A1(_06199_),
    .A2(_06075_),
    .ZN(_06268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30360_ (.A1(_06268_),
    .A2(net19528),
    .ZN(_06269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30361_ (.A1(net18455),
    .A2(net19505),
    .A3(_06080_),
    .ZN(_06270_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30362_ (.A1(_06269_),
    .A2(_06270_),
    .A3(net19482),
    .ZN(_06271_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30363_ (.A1(_06154_),
    .A2(net19497),
    .A3(_06167_),
    .ZN(_06272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30364_ (.A1(net19530),
    .A2(net18366),
    .ZN(_06273_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30365_ (.I(_06273_),
    .ZN(_06274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30366_ (.A1(_06274_),
    .A2(net19515),
    .B(net19483),
    .ZN(_06275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30367_ (.A1(_06272_),
    .A2(_06275_),
    .ZN(_06276_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30368_ (.A1(_06271_),
    .A2(_06276_),
    .A3(net19473),
    .ZN(_06277_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30369_ (.A1(_06267_),
    .A2(_06277_),
    .A3(net20395),
    .ZN(_06278_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30370_ (.A1(_06249_),
    .A2(_06159_),
    .A3(net19525),
    .ZN(_06279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30371_ (.A1(_06161_),
    .A2(net19539),
    .A3(net19504),
    .ZN(_06280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30372_ (.A1(_06279_),
    .A2(_06280_),
    .A3(net19495),
    .ZN(_06281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30373_ (.A1(net19011),
    .A2(net17650),
    .A3(net19500),
    .ZN(_06282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30374_ (.A1(net19003),
    .A2(net19519),
    .A3(net17654),
    .ZN(_06283_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30375_ (.A1(_06282_),
    .A2(_06283_),
    .A3(net19483),
    .ZN(_06284_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30376_ (.A1(_06281_),
    .A2(_06284_),
    .A3(net19473),
    .ZN(_06285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _30377_ (.A1(net19013),
    .A2(net19539),
    .B(net19515),
    .ZN(_06286_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30378_ (.A1(_06286_),
    .A2(net18031),
    .ZN(_06287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30379_ (.A1(_06239_),
    .A2(net19523),
    .B(net19487),
    .ZN(_06288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30380_ (.A1(_06287_),
    .A2(_06288_),
    .B(_06109_),
    .ZN(_06289_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30381_ (.A1(_06171_),
    .A2(net19512),
    .Z(_06290_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input57 (.I(net544),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30383_ (.A1(_06290_),
    .A2(net17647),
    .B(net19480),
    .ZN(_06292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30384_ (.A1(_06292_),
    .A2(_06201_),
    .ZN(_06293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30385_ (.A1(_06289_),
    .A2(_06293_),
    .ZN(_06294_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30386_ (.A1(_06285_),
    .A2(_06294_),
    .A3(_06187_),
    .ZN(_06295_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30387_ (.A1(_06278_),
    .A2(_06295_),
    .B(net20174),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30388_ (.A1(_06077_),
    .A2(_06180_),
    .ZN(_06297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30389_ (.A1(_06109_),
    .A2(net19476),
    .Z(_06298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30390_ (.A1(net19509),
    .A2(net19533),
    .ZN(_06299_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30391_ (.I(_06299_),
    .ZN(_06300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30392_ (.A1(_06300_),
    .A2(_06262_),
    .ZN(_06301_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _30393_ (.A1(_06280_),
    .A2(_06297_),
    .A3(_06298_),
    .A4(_06301_),
    .ZN(_06302_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30394_ (.I(_16163_[0]),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _30395_ (.A1(_06108_),
    .A2(_06303_),
    .A3(net19512),
    .Z(_06304_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30396_ (.A1(_06304_),
    .A2(net19476),
    .ZN(_06305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30397_ (.A1(_06217_),
    .A2(_06120_),
    .ZN(_06306_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30398_ (.A1(_06305_),
    .A2(_06306_),
    .B(_06142_),
    .ZN(_06307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30399_ (.A1(_06302_),
    .A2(_06307_),
    .ZN(_06308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30400_ (.A1(_06158_),
    .A2(_06166_),
    .ZN(_06309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30401_ (.A1(net19010),
    .A2(net19541),
    .ZN(_06310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30402_ (.A1(_06058_),
    .A2(net18450),
    .ZN(_06311_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _30403_ (.A1(_06309_),
    .A2(net19478),
    .A3(_06311_),
    .A4(net19928),
    .Z(_06312_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30404_ (.A1(_06308_),
    .A2(_06312_),
    .B(net20175),
    .ZN(_06313_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30405_ (.I(_06176_),
    .ZN(_06314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30406_ (.A1(_06314_),
    .A2(net19512),
    .ZN(_06315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30407_ (.A1(_06123_),
    .A2(net19517),
    .ZN(_06316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30408_ (.A1(net17234),
    .A2(_06316_),
    .Z(_06317_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _30409_ (.I(_06162_),
    .ZN(_06318_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30410_ (.A1(_06318_),
    .A2(net19522),
    .B(net19487),
    .ZN(_06319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30411_ (.I(_06209_),
    .ZN(_06320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30412_ (.A1(_06320_),
    .A2(net19497),
    .Z(_06321_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30413_ (.I(_06321_),
    .ZN(_06322_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30414_ (.A1(_06317_),
    .A2(_06319_),
    .A3(_06322_),
    .ZN(_06323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30415_ (.A1(net18458),
    .A2(_06180_),
    .ZN(_06324_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30416_ (.A1(_06324_),
    .A2(net19491),
    .A3(_06311_),
    .ZN(_06325_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30417_ (.A1(_06323_),
    .A2(_06325_),
    .A3(net19471),
    .ZN(_06326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30418_ (.A1(net18464),
    .A2(net18461),
    .ZN(_06327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30419_ (.A1(_06231_),
    .A2(net19487),
    .Z(_06328_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30420_ (.A1(_06327_),
    .A2(_06328_),
    .B(net19472),
    .ZN(_06329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30421_ (.A1(_06116_),
    .A2(net19515),
    .Z(_06330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30422_ (.A1(net19535),
    .A2(net18034),
    .ZN(_06331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30423_ (.A1(_06330_),
    .A2(_06331_),
    .ZN(_06332_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30424_ (.A1(_06272_),
    .A2(net19477),
    .A3(_06332_),
    .ZN(_06333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30425_ (.A1(_06329_),
    .A2(_06333_),
    .ZN(_06334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30426_ (.A1(_06326_),
    .A2(_06334_),
    .B(net20176),
    .ZN(_06335_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30427_ (.A1(_06313_),
    .A2(_06335_),
    .ZN(_06336_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30428_ (.A1(_06336_),
    .A2(_06296_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30429_ (.A1(_06161_),
    .A2(_06249_),
    .A3(net19502),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30430_ (.A1(_06053_),
    .A2(net19515),
    .Z(_06338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30431_ (.A1(_06338_),
    .A2(_06080_),
    .ZN(_06339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30432_ (.A1(_06337_),
    .A2(_06339_),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input56 (.I(key[34]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30434_ (.A1(_06340_),
    .A2(net19480),
    .ZN(_06342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30435_ (.A1(_06161_),
    .A2(net19533),
    .ZN(_06343_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30436_ (.A1(_06197_),
    .A2(net19505),
    .Z(_06344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30437_ (.A1(_06343_),
    .A2(_06344_),
    .ZN(_06345_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input55 (.I(key[33]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30439_ (.A1(_06345_),
    .A2(net19489),
    .A3(_06250_),
    .ZN(_06347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30440_ (.A1(_06342_),
    .A2(_06347_),
    .ZN(_06348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30441_ (.A1(_06348_),
    .A2(net19929),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30442_ (.A1(_06154_),
    .A2(net19508),
    .A3(net17648),
    .ZN(_06350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30443_ (.A1(_06061_),
    .A2(net19515),
    .ZN(_06351_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30444_ (.A1(_06350_),
    .A2(net18024),
    .A3(net19495),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30445_ (.A1(net18456),
    .A2(net19524),
    .A3(net490),
    .ZN(_06353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30446_ (.A1(net19006),
    .A2(net18030),
    .ZN(_06354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30447_ (.A1(_06354_),
    .A2(net19507),
    .ZN(_06355_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30448_ (.A1(_06353_),
    .A2(_06355_),
    .A3(net19481),
    .ZN(_06356_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30449_ (.A1(_06352_),
    .A2(net19467),
    .A3(_06356_),
    .ZN(_06357_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30450_ (.A1(_06349_),
    .A2(_06357_),
    .A3(_06187_),
    .ZN(_06358_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30451_ (.A1(_06075_),
    .A2(net17636),
    .A3(net19518),
    .ZN(_06359_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30452_ (.A1(net17649),
    .A2(net18028),
    .A3(net19497),
    .ZN(_06360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30453_ (.A1(_06360_),
    .A2(_06359_),
    .ZN(_06361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30454_ (.A1(_06361_),
    .A2(net19493),
    .ZN(_06362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30455_ (.A1(net18448),
    .A2(net19500),
    .A3(net18026),
    .ZN(_06363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30456_ (.A1(net19541),
    .A2(_16153_[0]),
    .ZN(_06364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30457_ (.A1(_06157_),
    .A2(_06364_),
    .A3(net19519),
    .ZN(_06365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30458_ (.A1(_06363_),
    .A2(_06365_),
    .A3(net19485),
    .ZN(_06366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30459_ (.A1(_06362_),
    .A2(_06366_),
    .ZN(_06367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30460_ (.A1(_06367_),
    .A2(net19473),
    .ZN(_06368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30461_ (.A1(net17642),
    .A2(net19506),
    .ZN(_06369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30462_ (.A1(_06364_),
    .A2(net18026),
    .ZN(_06370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30463_ (.A1(_06370_),
    .A2(net19526),
    .ZN(_06371_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30464_ (.A1(_06369_),
    .A2(_06371_),
    .A3(net19480),
    .ZN(_06372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30465_ (.A1(net19536),
    .A2(net18035),
    .ZN(_06373_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30466_ (.A1(_06199_),
    .A2(net19505),
    .A3(_06373_),
    .ZN(_06374_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30467_ (.A1(_06374_),
    .A2(_06236_),
    .A3(net19488),
    .ZN(_06375_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30468_ (.A1(_06372_),
    .A2(_06375_),
    .A3(net19929),
    .ZN(_06376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30469_ (.A1(_06368_),
    .A2(_06376_),
    .A3(net20395),
    .ZN(_06377_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30470_ (.A1(_06358_),
    .A2(_06377_),
    .A3(net20175),
    .ZN(_06378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30471_ (.A1(_06310_),
    .A2(_06032_),
    .ZN(_06379_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30472_ (.A1(_06122_),
    .A2(_06052_),
    .Z(_06380_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30473_ (.A1(net19535),
    .A2(net17635),
    .ZN(_06381_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30474_ (.A1(_06379_),
    .A2(_06381_),
    .B(net19512),
    .ZN(_06382_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30475_ (.A1(_06382_),
    .A2(net19476),
    .A3(_06306_),
    .ZN(_06383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30476_ (.A1(_06314_),
    .A2(net19520),
    .ZN(_06384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input54 (.I(net552),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30478_ (.A1(_06384_),
    .A2(net19493),
    .Z(_06386_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30479_ (.I(_06231_),
    .ZN(_06387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30480_ (.A1(_06387_),
    .A2(_06373_),
    .ZN(_06388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30481_ (.A1(_06386_),
    .A2(_06388_),
    .B(net19928),
    .ZN(_06389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30482_ (.A1(_06383_),
    .A2(_06389_),
    .ZN(_06390_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30483_ (.A1(net19515),
    .A2(_16158_[0]),
    .Z(_06391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30484_ (.A1(_06351_),
    .A2(_06391_),
    .ZN(_06392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30485_ (.A1(_06392_),
    .A2(net19482),
    .Z(_06393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30486_ (.A1(_16167_[0]),
    .A2(net19515),
    .B(net19493),
    .ZN(_06394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30487_ (.A1(_06337_),
    .A2(_06394_),
    .B(_06109_),
    .ZN(_06395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30488_ (.A1(_06393_),
    .A2(_06395_),
    .ZN(_06396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30489_ (.A1(_06390_),
    .A2(_06396_),
    .A3(_06187_),
    .ZN(_06397_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30490_ (.A1(_06149_),
    .A2(net19502),
    .Z(_06398_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30491_ (.A1(_06398_),
    .A2(net18029),
    .Z(_06399_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _30492_ (.A1(_06249_),
    .A2(net19525),
    .A3(_06146_),
    .Z(_06400_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30493_ (.A1(_06399_),
    .A2(_06400_),
    .B(net19481),
    .ZN(_06401_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30494_ (.A1(_06249_),
    .A2(_06159_),
    .A3(net19501),
    .ZN(_06402_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30495_ (.A1(_06402_),
    .A2(net19494),
    .Z(_06403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30496_ (.A1(net19519),
    .A2(net18025),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30497_ (.A1(_06403_),
    .A2(_06404_),
    .ZN(_06405_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30498_ (.A1(_06401_),
    .A2(_06405_),
    .A3(net19928),
    .ZN(_06406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30499_ (.A1(_06290_),
    .A2(net18453),
    .ZN(_06407_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30500_ (.A1(net18363),
    .A2(net19515),
    .B(net19476),
    .ZN(_06408_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30501_ (.A1(_06407_),
    .A2(_06408_),
    .B(net19928),
    .ZN(_06409_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30502_ (.A1(net18449),
    .A2(net19504),
    .A3(_06075_),
    .ZN(_06410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30503_ (.A1(_06250_),
    .A2(_06410_),
    .A3(net19480),
    .ZN(_06411_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30504_ (.A1(_06409_),
    .A2(_06411_),
    .B(_06187_),
    .ZN(_06412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30505_ (.A1(_06406_),
    .A2(_06412_),
    .ZN(_06413_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30506_ (.I(_06194_),
    .ZN(_06414_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30507_ (.A1(_06397_),
    .A2(_06413_),
    .A3(net19927),
    .ZN(_06415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30508_ (.A1(_06378_),
    .A2(_06415_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30509_ (.A1(_06217_),
    .A2(net18452),
    .Z(_06416_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30510_ (.A1(_06416_),
    .A2(net17235),
    .B(net19930),
    .ZN(_06417_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30511_ (.A1(net19527),
    .A2(_06257_),
    .ZN(_06418_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30512_ (.I(_06418_),
    .ZN(_06419_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30513_ (.A1(_06419_),
    .A2(net19466),
    .B(_06221_),
    .ZN(_06420_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30514_ (.A1(_06417_),
    .A2(_06420_),
    .B(net20395),
    .ZN(_06421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30515_ (.A1(_06380_),
    .A2(net19532),
    .B(net19515),
    .ZN(_06422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30516_ (.A1(net17369),
    .A2(net17652),
    .ZN(_06423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30517_ (.A1(_06051_),
    .A2(net17649),
    .ZN(_06424_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30518_ (.A1(_06423_),
    .A2(_06424_),
    .A3(net19928),
    .ZN(_06425_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _30519_ (.A1(_06234_),
    .A2(net19515),
    .Z(_06426_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30520_ (.A1(_06359_),
    .A2(_06109_),
    .A3(_06426_),
    .ZN(_06427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30521_ (.A1(_06425_),
    .A2(_06427_),
    .ZN(_06428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30522_ (.A1(_06428_),
    .A2(net19487),
    .ZN(_06429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30523_ (.A1(_06429_),
    .A2(_06421_),
    .ZN(_06430_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30524_ (.A1(_06279_),
    .A2(_06207_),
    .A3(net19495),
    .ZN(_06431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30525_ (.A1(_06032_),
    .A2(_06234_),
    .ZN(_06432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30526_ (.A1(_06432_),
    .A2(net19505),
    .ZN(_06433_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30527_ (.A1(_06080_),
    .A2(net17650),
    .A3(net19527),
    .ZN(_06434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30528_ (.A1(_06433_),
    .A2(_06434_),
    .A3(net19481),
    .ZN(_06435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30529_ (.A1(_06431_),
    .A2(_06435_),
    .ZN(_06436_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30530_ (.A1(_06436_),
    .A2(_06109_),
    .ZN(_06437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30531_ (.A1(_06422_),
    .A2(net17638),
    .ZN(_06438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30532_ (.A1(_06438_),
    .A2(_06306_),
    .ZN(_06439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30533_ (.A1(_06439_),
    .A2(net19487),
    .ZN(_06440_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30534_ (.A1(_06365_),
    .A2(net19476),
    .B(_06109_),
    .ZN(_06441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30535_ (.A1(_06440_),
    .A2(_06441_),
    .ZN(_06442_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30536_ (.A1(_06437_),
    .A2(net20395),
    .A3(_06442_),
    .ZN(_06443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30537_ (.A1(_06430_),
    .A2(_06443_),
    .ZN(_06444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30538_ (.A1(_06444_),
    .A2(net20174),
    .ZN(_06445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30539_ (.A1(_06309_),
    .A2(_06174_),
    .ZN(_06446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30540_ (.A1(_06446_),
    .A2(net19478),
    .ZN(_06447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30541_ (.A1(net18458),
    .A2(net18457),
    .ZN(_06448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30542_ (.A1(_06168_),
    .A2(net19511),
    .ZN(_06449_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30543_ (.A1(_06448_),
    .A2(_06449_),
    .A3(net19491),
    .ZN(_06450_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30544_ (.A1(_06447_),
    .A2(_06450_),
    .A3(net19928),
    .ZN(_06451_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30545_ (.A1(net17373),
    .A2(net17379),
    .B(net19513),
    .ZN(_06452_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30546_ (.A1(_06318_),
    .A2(_06150_),
    .B(net19524),
    .ZN(_06453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30547_ (.A1(_06452_),
    .A2(_06453_),
    .A3(net19478),
    .ZN(_06454_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30548_ (.A1(_06167_),
    .A2(net19515),
    .Z(_06455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30549_ (.A1(_06455_),
    .A2(net18450),
    .ZN(_06456_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30550_ (.A1(net17647),
    .A2(_06373_),
    .A3(net19505),
    .ZN(_06457_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30551_ (.A1(_06456_),
    .A2(net19488),
    .A3(_06457_),
    .ZN(_06458_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30552_ (.A1(_06454_),
    .A2(_06458_),
    .A3(net19470),
    .ZN(_06459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30553_ (.A1(_06451_),
    .A2(_06459_),
    .A3(net20176),
    .ZN(_06460_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30554_ (.A1(_06398_),
    .A2(net18448),
    .A3(net19004),
    .ZN(_06461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30555_ (.I(_06268_),
    .ZN(_06462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30556_ (.A1(_06462_),
    .A2(net17639),
    .ZN(_06463_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30557_ (.A1(_06461_),
    .A2(_06463_),
    .A3(net19495),
    .ZN(_06464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30558_ (.A1(_06153_),
    .A2(net17643),
    .ZN(_06465_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30559_ (.A1(_06465_),
    .A2(_06163_),
    .A3(net19481),
    .ZN(_06466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30560_ (.A1(_06464_),
    .A2(_06466_),
    .ZN(_06467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30561_ (.A1(_06467_),
    .A2(net19469),
    .ZN(_06468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30562_ (.A1(_06455_),
    .A2(net17637),
    .ZN(_06469_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30563_ (.A1(_06469_),
    .A2(_06270_),
    .A3(net19482),
    .ZN(_06470_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30564_ (.A1(net19002),
    .A2(net19495),
    .Z(_06471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30565_ (.A1(_06161_),
    .A2(net19005),
    .ZN(_06472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30566_ (.A1(_06471_),
    .A2(_06472_),
    .B(net19469),
    .ZN(_06473_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30567_ (.A1(_06470_),
    .A2(_06473_),
    .B(_06187_),
    .ZN(_06474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30568_ (.A1(_06468_),
    .A2(_06474_),
    .ZN(_06475_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30569_ (.A1(_06460_),
    .A2(_06475_),
    .A3(net19926),
    .ZN(_06476_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30570_ (.A1(_06445_),
    .A2(_06476_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _30571_ (.A1(net17375),
    .A2(net19492),
    .A3(_06123_),
    .ZN(_06477_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30572_ (.A1(_06477_),
    .A2(net19930),
    .ZN(_06478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30573_ (.A1(_06286_),
    .A2(net19007),
    .ZN(_06479_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30574_ (.A1(_06479_),
    .A2(_06297_),
    .A3(net19491),
    .ZN(_06480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30575_ (.A1(_06478_),
    .A2(_06480_),
    .B(_06187_),
    .ZN(_06481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30576_ (.A1(_06403_),
    .A2(_06309_),
    .ZN(_06482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30577_ (.A1(net18455),
    .A2(net19505),
    .Z(_06483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30578_ (.A1(_06483_),
    .A2(net18032),
    .ZN(_06484_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30579_ (.A1(_06199_),
    .A2(_06262_),
    .A3(net19521),
    .ZN(_06485_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30580_ (.A1(_06484_),
    .A2(net19480),
    .A3(_06485_),
    .ZN(_06486_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30581_ (.A1(_06482_),
    .A2(_06486_),
    .A3(net19929),
    .ZN(_06487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30582_ (.A1(_06481_),
    .A2(_06487_),
    .B(net20174),
    .ZN(_06488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30583_ (.A1(_06218_),
    .A2(net19504),
    .ZN(_06489_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30584_ (.A1(net18460),
    .A2(net18023),
    .B(_06339_),
    .C(net19476),
    .ZN(_06490_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30585_ (.A1(_06315_),
    .A2(net19487),
    .Z(_06491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30586_ (.A1(net19013),
    .A2(net19505),
    .ZN(_06492_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30587_ (.A1(_06492_),
    .A2(net19533),
    .Z(_06493_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30588_ (.A1(net17378),
    .A2(net17203),
    .A3(_06493_),
    .ZN(_06494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30589_ (.A1(_06490_),
    .A2(_06494_),
    .A3(net19930),
    .ZN(_06495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30590_ (.A1(_06426_),
    .A2(net19484),
    .Z(_06496_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30591_ (.A1(_06496_),
    .A2(_06236_),
    .A3(_06322_),
    .ZN(_06497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30592_ (.A1(net17371),
    .A2(_06171_),
    .ZN(_06498_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30593_ (.A1(_06226_),
    .A2(_06498_),
    .A3(net19487),
    .ZN(_06499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30594_ (.A1(_06497_),
    .A2(_06499_),
    .A3(_06109_),
    .ZN(_06500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30595_ (.A1(_06495_),
    .A2(_06500_),
    .A3(_06187_),
    .ZN(_06501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30596_ (.A1(_06488_),
    .A2(_06501_),
    .ZN(_06502_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30597_ (.A1(net17375),
    .A2(net19006),
    .ZN(_06503_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30598_ (.A1(net18457),
    .A2(net18450),
    .A3(net19521),
    .ZN(_06504_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30599_ (.A1(_06503_),
    .A2(_06504_),
    .A3(net19480),
    .ZN(_06505_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30600_ (.A1(_06246_),
    .A2(_06163_),
    .A3(net19490),
    .ZN(_06506_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30601_ (.A1(_06505_),
    .A2(_06506_),
    .A3(net19928),
    .ZN(_06507_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30602_ (.I(net18364),
    .ZN(_06508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30603_ (.A1(net19515),
    .A2(_06508_),
    .ZN(_06509_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30604_ (.A1(net19516),
    .A2(_06320_),
    .B(_06509_),
    .C(net19487),
    .ZN(_06510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30605_ (.A1(_06510_),
    .A2(_06109_),
    .ZN(_06511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30606_ (.I(_06511_),
    .ZN(_06512_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30607_ (.A1(_06343_),
    .A2(net19513),
    .Z(_06513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30608_ (.A1(_06225_),
    .A2(net491),
    .ZN(_06514_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30609_ (.A1(_06513_),
    .A2(net17233),
    .A3(net19479),
    .ZN(_06515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30610_ (.A1(_06512_),
    .A2(_06515_),
    .ZN(_06516_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30611_ (.A1(_06507_),
    .A2(_06516_),
    .A3(_06187_),
    .ZN(_06517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30612_ (.A1(_06121_),
    .A2(net19489),
    .Z(_06518_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30613_ (.A1(_06338_),
    .A2(net18028),
    .Z(_06519_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30614_ (.I(_06519_),
    .ZN(_06520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30615_ (.A1(_06518_),
    .A2(_06520_),
    .ZN(_06521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30616_ (.A1(_06331_),
    .A2(net19517),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30617_ (.A1(_06522_),
    .A2(net19477),
    .Z(_06523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30618_ (.A1(net18459),
    .A2(net19504),
    .ZN(_06524_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30619_ (.A1(_06523_),
    .A2(_06524_),
    .B(net19930),
    .ZN(_06525_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30620_ (.A1(_06521_),
    .A2(_06525_),
    .ZN(_06526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30621_ (.A1(_06158_),
    .A2(_06080_),
    .ZN(_06527_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30622_ (.A1(net19538),
    .A2(net19497),
    .B(net19483),
    .ZN(_06528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30623_ (.A1(_06527_),
    .A2(_06528_),
    .B(_06109_),
    .ZN(_06529_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30624_ (.A1(_06057_),
    .A2(_06126_),
    .B(net19476),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30625_ (.A1(_06128_),
    .A2(_06384_),
    .ZN(_06531_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30626_ (.A1(_06530_),
    .A2(_06531_),
    .Z(_06532_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30627_ (.A1(_06529_),
    .A2(_06532_),
    .ZN(_06533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30628_ (.A1(_06526_),
    .A2(_06533_),
    .A3(net20395),
    .ZN(_06534_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30629_ (.A1(_06517_),
    .A2(_06534_),
    .A3(net20174),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30630_ (.A1(_06502_),
    .A2(_06535_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30631_ (.I(_06249_),
    .ZN(_06536_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30632_ (.A1(_06522_),
    .A2(_06536_),
    .ZN(_06537_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30633_ (.A1(_06537_),
    .A2(_06321_),
    .B(net19477),
    .ZN(_06538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30634_ (.A1(_06387_),
    .A2(_06146_),
    .ZN(_06539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30635_ (.A1(net19519),
    .A2(_06364_),
    .B(net19483),
    .ZN(_06540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30636_ (.A1(_06539_),
    .A2(_06540_),
    .ZN(_06541_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30637_ (.A1(_06538_),
    .A2(net19928),
    .A3(_06541_),
    .ZN(_06542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30638_ (.A1(_06542_),
    .A2(_06187_),
    .ZN(_06543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30639_ (.A1(net18464),
    .A2(net18451),
    .ZN(_06544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30640_ (.A1(_06544_),
    .A2(net19476),
    .ZN(_06545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30641_ (.A1(net18461),
    .A2(net18027),
    .B(net19517),
    .ZN(_06546_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30642_ (.A1(_06545_),
    .A2(_06546_),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30643_ (.A1(_06485_),
    .A2(_06492_),
    .B(net19478),
    .ZN(_06548_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _30644_ (.A1(_06547_),
    .A2(_06548_),
    .A3(net19930),
    .ZN(_06549_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30645_ (.A1(_06543_),
    .A2(_06549_),
    .ZN(_06550_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30646_ (.A1(net17638),
    .A2(net19518),
    .Z(_06551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30647_ (.A1(_06551_),
    .A2(net18453),
    .ZN(_06552_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30648_ (.A1(net17646),
    .A2(net18366),
    .B(net19499),
    .ZN(_06553_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30649_ (.A1(_06552_),
    .A2(net19485),
    .A3(_06553_),
    .ZN(_06554_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30650_ (.A1(net17652),
    .A2(net17654),
    .A3(net19498),
    .ZN(_06555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30651_ (.A1(_06125_),
    .A2(_06128_),
    .A3(_06555_),
    .ZN(_06556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30652_ (.A1(_06554_),
    .A2(_06556_),
    .A3(net19475),
    .ZN(_06557_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30653_ (.A1(_06153_),
    .A2(net19481),
    .ZN(_06558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30654_ (.A1(_06433_),
    .A2(_06558_),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30655_ (.A1(net17370),
    .A2(net19488),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30656_ (.A1(_06560_),
    .A2(_06280_),
    .ZN(_06561_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30657_ (.A1(_06559_),
    .A2(_06561_),
    .A3(net19930),
    .ZN(_06562_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30658_ (.A1(_06562_),
    .A2(_06557_),
    .B(_06187_),
    .ZN(_06563_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30659_ (.A1(_06563_),
    .A2(_06550_),
    .B(net19926),
    .ZN(_06564_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30660_ (.A1(net19545),
    .A2(net19502),
    .B(net19476),
    .ZN(_06565_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30661_ (.A1(_06160_),
    .A2(_06565_),
    .B(net19928),
    .ZN(_06566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30662_ (.A1(net18463),
    .A2(_06387_),
    .ZN(_06567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30663_ (.A1(_06551_),
    .A2(_06199_),
    .ZN(_06568_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30664_ (.A1(_06567_),
    .A2(_06568_),
    .A3(net19481),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30665_ (.A1(_06566_),
    .A2(_06569_),
    .B(_06187_),
    .ZN(_06570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30666_ (.A1(net17642),
    .A2(net19524),
    .ZN(_06571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30667_ (.A1(_06518_),
    .A2(_06571_),
    .ZN(_06572_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30668_ (.A1(net18462),
    .A2(net19524),
    .A3(net17653),
    .ZN(_06573_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30669_ (.I(_06177_),
    .ZN(_06574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30670_ (.A1(net17368),
    .A2(net19511),
    .B(net19490),
    .ZN(_06575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30671_ (.A1(_06573_),
    .A2(_06575_),
    .B(net19470),
    .ZN(_06576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30672_ (.A1(_06572_),
    .A2(_06576_),
    .ZN(_06577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30673_ (.A1(_06570_),
    .A2(_06577_),
    .ZN(_06578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30674_ (.A1(net17634),
    .A2(net17653),
    .ZN(_06579_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30675_ (.A1(_06387_),
    .A2(net18027),
    .ZN(_06580_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30676_ (.A1(_06579_),
    .A2(_06580_),
    .A3(net19480),
    .ZN(_06581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30677_ (.A1(_06148_),
    .A2(net19507),
    .B(net19481),
    .ZN(_06582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30678_ (.A1(net18462),
    .A2(net19524),
    .ZN(_06583_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30679_ (.A1(_06582_),
    .A2(_06583_),
    .B(net19468),
    .ZN(_06584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30680_ (.A1(_06581_),
    .A2(_06584_),
    .ZN(_06585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30681_ (.A1(_06288_),
    .A2(net17380),
    .B(net19928),
    .ZN(_06586_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30682_ (.A1(_06061_),
    .A2(net18462),
    .A3(net19524),
    .ZN(_06587_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30683_ (.A1(net17369),
    .A2(net19484),
    .ZN(_06588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30684_ (.A1(_06587_),
    .A2(_06588_),
    .ZN(_06589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30685_ (.A1(_06586_),
    .A2(_06589_),
    .ZN(_06590_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30686_ (.A1(_06585_),
    .A2(_06590_),
    .A3(_06187_),
    .ZN(_06591_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30687_ (.A1(_06578_),
    .A2(_06591_),
    .A3(net20175),
    .ZN(_06592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30688_ (.A1(_06564_),
    .A2(_06592_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30689_ (.I(_06217_),
    .ZN(_06593_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30690_ (.A1(_06514_),
    .A2(_06593_),
    .ZN(_06594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30691_ (.A1(_06594_),
    .A2(net19476),
    .ZN(_06595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30692_ (.A1(_06345_),
    .A2(net19491),
    .ZN(_06596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30693_ (.A1(_06595_),
    .A2(_06596_),
    .ZN(_06597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30694_ (.A1(_06597_),
    .A2(net19928),
    .ZN(_06598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30695_ (.A1(_06083_),
    .A2(net18033),
    .ZN(_06599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30696_ (.A1(_06319_),
    .A2(_06599_),
    .ZN(_06600_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30697_ (.I(_16157_[0]),
    .ZN(_06601_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30698_ (.A1(_06601_),
    .A2(net19497),
    .B(net19486),
    .ZN(_06602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30699_ (.A1(_06568_),
    .A2(_06602_),
    .ZN(_06603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30700_ (.A1(_06600_),
    .A2(_06603_),
    .A3(net19470),
    .ZN(_06604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30701_ (.A1(_06598_),
    .A2(net20176),
    .A3(_06604_),
    .ZN(_06605_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30702_ (.A1(net19013),
    .A2(net19508),
    .B(_06472_),
    .C(net19495),
    .ZN(_06606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30703_ (.A1(_06472_),
    .A2(net19508),
    .ZN(_06607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30704_ (.A1(_06330_),
    .A2(net19004),
    .ZN(_06608_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30705_ (.A1(_06607_),
    .A2(_06608_),
    .A3(net19481),
    .ZN(_06609_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30706_ (.A1(_06606_),
    .A2(_06609_),
    .A3(net19469),
    .ZN(_06610_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30707_ (.A1(net18033),
    .A2(net19511),
    .Z(_06611_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30708_ (.A1(_06433_),
    .A2(net19490),
    .A3(_06611_),
    .ZN(_06612_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30709_ (.A1(_06286_),
    .A2(net19490),
    .ZN(_06613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30710_ (.A1(_06613_),
    .A2(_06078_),
    .ZN(_06614_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30711_ (.A1(_06612_),
    .A2(_06614_),
    .A3(net19928),
    .ZN(_06615_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30712_ (.A1(_06610_),
    .A2(net20395),
    .A3(_06615_),
    .ZN(_06616_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30713_ (.A1(_06605_),
    .A2(_06616_),
    .A3(net20175),
    .ZN(_06617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30714_ (.A1(net17640),
    .A2(net19498),
    .ZN(_06618_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30715_ (.A1(_06384_),
    .A2(_06618_),
    .Z(_06619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30716_ (.A1(_06496_),
    .A2(_06619_),
    .B(net19928),
    .ZN(_06620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30717_ (.A1(_06310_),
    .A2(net19497),
    .Z(_06621_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30718_ (.A1(_06621_),
    .A2(_06161_),
    .ZN(_06622_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30719_ (.A1(_16156_[0]),
    .A2(net18362),
    .B(net19515),
    .ZN(_06623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30720_ (.A1(net17633),
    .A2(net19493),
    .A3(_06623_),
    .ZN(_06624_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30721_ (.A1(_06620_),
    .A2(_06624_),
    .B(_06187_),
    .ZN(_06625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30722_ (.A1(_06379_),
    .A2(net19512),
    .ZN(_06626_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30723_ (.A1(_06626_),
    .A2(_06220_),
    .Z(_06627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30724_ (.A1(_06330_),
    .A2(net17638),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30725_ (.A1(_06628_),
    .A2(net19487),
    .Z(_06629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30726_ (.A1(_06627_),
    .A2(_06629_),
    .ZN(_06630_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30727_ (.A1(_06235_),
    .A2(net17641),
    .B(net19504),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30728_ (.A1(net17639),
    .A2(net19005),
    .ZN(_06632_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30729_ (.A1(_06631_),
    .A2(net19480),
    .A3(_06632_),
    .ZN(_06633_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30730_ (.A1(_06630_),
    .A2(_06633_),
    .A3(net19928),
    .ZN(_06634_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30731_ (.A1(_06625_),
    .A2(_06634_),
    .ZN(_06635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30732_ (.A1(_06316_),
    .A2(net19492),
    .ZN(_06636_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30733_ (.A1(_06519_),
    .A2(_06636_),
    .ZN(_06637_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30734_ (.A1(_06489_),
    .A2(_06318_),
    .Z(_06638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30735_ (.A1(_06637_),
    .A2(_06638_),
    .ZN(_06639_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30736_ (.A1(net17368),
    .A2(net19517),
    .B(net19492),
    .ZN(_06640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30737_ (.A1(_06157_),
    .A2(net19013),
    .ZN(_06641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30738_ (.A1(net18447),
    .A2(net19513),
    .ZN(_06642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30739_ (.A1(_06640_),
    .A2(_06642_),
    .B(net19471),
    .ZN(_06643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30740_ (.A1(_06639_),
    .A2(_06643_),
    .B(net20395),
    .ZN(_06644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30741_ (.A1(_06392_),
    .A2(_06418_),
    .ZN(_06645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30742_ (.A1(net19481),
    .A2(_06645_),
    .ZN(_06646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30743_ (.A1(net17650),
    .A2(net18030),
    .ZN(_06647_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30744_ (.A1(_06647_),
    .A2(net19528),
    .B(net19481),
    .ZN(_06648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30745_ (.A1(_06483_),
    .A2(_06061_),
    .ZN(_06649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30746_ (.A1(_06648_),
    .A2(_06649_),
    .B(net19928),
    .ZN(_06650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30747_ (.A1(_06650_),
    .A2(_06646_),
    .ZN(_06651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30748_ (.A1(_06651_),
    .A2(_06644_),
    .ZN(_06652_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30749_ (.A1(_06652_),
    .A2(_06635_),
    .A3(net19926),
    .ZN(_06653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30750_ (.A1(_06653_),
    .A2(_06617_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30751_ (.A1(_06199_),
    .A2(net19011),
    .A3(net19515),
    .ZN(_06654_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30752_ (.A1(_06167_),
    .A2(_06171_),
    .A3(net19497),
    .ZN(_06655_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30753_ (.A1(_06654_),
    .A2(_06655_),
    .ZN(_06656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30754_ (.A1(_06656_),
    .A2(net19486),
    .ZN(_06657_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30755_ (.A1(_06171_),
    .A2(_06234_),
    .A3(net19515),
    .ZN(_06658_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30756_ (.A1(net19515),
    .A2(_16165_[0]),
    .Z(_06659_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30757_ (.A1(_06658_),
    .A2(net19493),
    .A3(_06659_),
    .ZN(_06660_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30758_ (.A1(_06657_),
    .A2(net19928),
    .A3(_06660_),
    .ZN(_06661_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30759_ (.A1(_06641_),
    .A2(net19515),
    .Z(_06662_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30760_ (.A1(net19515),
    .A2(_16151_[0]),
    .ZN(_06663_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30761_ (.A1(_06663_),
    .A2(net19483),
    .ZN(_06664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30762_ (.A1(_06664_),
    .A2(_06204_),
    .ZN(_06665_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30763_ (.A1(_06530_),
    .A2(_06662_),
    .B(_06665_),
    .ZN(_06666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30764_ (.A1(_06666_),
    .A2(net19475),
    .ZN(_06667_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30765_ (.A1(_06661_),
    .A2(_06667_),
    .A3(_06187_),
    .ZN(_06668_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30766_ (.A1(_06668_),
    .A2(_06414_),
    .ZN(_06669_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30767_ (.A1(_06249_),
    .A2(_06262_),
    .A3(net19516),
    .ZN(_06670_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30768_ (.A1(_06438_),
    .A2(_06670_),
    .B(net19487),
    .ZN(_06671_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30769_ (.A1(_06231_),
    .A2(_06574_),
    .B(net19487),
    .ZN(_06672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30770_ (.A1(net17644),
    .A2(net19529),
    .ZN(_06673_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30771_ (.A1(_06379_),
    .A2(_06673_),
    .ZN(_06674_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30772_ (.A1(_06672_),
    .A2(_06674_),
    .ZN(_06675_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30773_ (.A1(_06671_),
    .A2(_06675_),
    .B(net19466),
    .ZN(_06676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30774_ (.A1(net18366),
    .A2(net19515),
    .B(net19496),
    .ZN(_06677_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30775_ (.A1(_06622_),
    .A2(_06677_),
    .B(_06109_),
    .ZN(_06678_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30776_ (.A1(net19520),
    .A2(_06126_),
    .B(_06673_),
    .ZN(_06679_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30777_ (.A1(_06679_),
    .A2(_06491_),
    .A3(_06204_),
    .ZN(_06680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30778_ (.A1(_06678_),
    .A2(_06680_),
    .ZN(_06681_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30779_ (.A1(_06676_),
    .A2(_06681_),
    .B(_06187_),
    .ZN(_06682_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30780_ (.A1(_06669_),
    .A2(_06682_),
    .ZN(_06683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30781_ (.A1(_06113_),
    .A2(_06154_),
    .ZN(_06684_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30782_ (.A1(_06684_),
    .A2(_06402_),
    .A3(net19494),
    .ZN(_06685_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30783_ (.A1(net18448),
    .A2(net19502),
    .A3(net19005),
    .ZN(_06686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30784_ (.A1(net19515),
    .A2(net19545),
    .ZN(_06687_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30785_ (.A1(_06686_),
    .A2(net19476),
    .A3(_06687_),
    .ZN(_06688_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30786_ (.A1(_06685_),
    .A2(net19474),
    .A3(_06688_),
    .ZN(_06689_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30787_ (.A1(_06455_),
    .A2(_06154_),
    .ZN(_06690_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30788_ (.A1(_06690_),
    .A2(_06489_),
    .A3(net19476),
    .ZN(_06691_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30789_ (.A1(_06418_),
    .A2(net19488),
    .A3(_06301_),
    .ZN(_06692_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30790_ (.A1(_06692_),
    .A2(net19930),
    .A3(_06691_),
    .ZN(_06693_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30791_ (.A1(_06689_),
    .A2(_06187_),
    .A3(_06693_),
    .ZN(_06694_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30792_ (.A1(net17647),
    .A2(net19517),
    .B(_06108_),
    .ZN(_06695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30793_ (.A1(_06514_),
    .A2(_06695_),
    .B(net19476),
    .ZN(_06696_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30794_ (.A1(_06628_),
    .A2(_06410_),
    .A3(net19930),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30795_ (.A1(_06696_),
    .A2(_06697_),
    .B(_06187_),
    .ZN(_06698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30796_ (.A1(_06051_),
    .A2(net18454),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30797_ (.A1(net17372),
    .A2(net19512),
    .B(_06108_),
    .ZN(_06700_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30798_ (.A1(_06626_),
    .A2(_06699_),
    .A3(_06700_),
    .ZN(_06701_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30799_ (.A1(_06290_),
    .A2(net17647),
    .ZN(_06702_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30800_ (.A1(_06424_),
    .A2(_06702_),
    .A3(net19930),
    .ZN(_06703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30801_ (.A1(_06701_),
    .A2(_06703_),
    .A3(net19476),
    .ZN(_06704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30802_ (.A1(_06698_),
    .A2(_06704_),
    .ZN(_06705_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30803_ (.A1(_06705_),
    .A2(_06694_),
    .B(_06414_),
    .ZN(_06706_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30804_ (.A1(_06706_),
    .A2(_06683_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30805_ (.A1(_03780_),
    .A2(_03769_),
    .ZN(_06707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30806_ (.A1(_12833_),
    .A2(_03776_),
    .ZN(_06708_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30807_ (.A1(_06708_),
    .A2(_06707_),
    .ZN(_06709_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _30808_ (.I(_06709_),
    .ZN(_06710_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30809_ (.A1(net21328),
    .A2(_12774_),
    .ZN(_06711_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30810_ (.A1(_12765_),
    .A2(net21008),
    .ZN(_06712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30811_ (.A1(_06712_),
    .A2(_06711_),
    .ZN(_06713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30812_ (.A1(_06710_),
    .A2(net20626),
    .ZN(_06714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30813_ (.I(_06713_),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30814_ (.A1(_06715_),
    .A2(net463),
    .ZN(_06716_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30815_ (.A1(_06716_),
    .A2(_06714_),
    .A3(net21089),
    .ZN(_06717_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30816_ (.I(net21147),
    .ZN(_06718_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30817_ (.A1(net21089),
    .A2(\text_in_r[1] ),
    .Z(_06719_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30818_ (.A1(_06718_),
    .A2(net19925),
    .A3(net20925),
    .ZN(_06720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30819_ (.A1(_06710_),
    .A2(_06715_),
    .ZN(_06721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30820_ (.A1(_06709_),
    .A2(net20626),
    .ZN(_06722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30821_ (.A1(_06722_),
    .A2(net21089),
    .A3(_06721_),
    .ZN(_06723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30822_ (.A1(net21486),
    .A2(\text_in_r[1] ),
    .ZN(_06724_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30823_ (.A1(net19924),
    .A2(net21147),
    .A3(_06724_),
    .ZN(_06725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30824_ (.A1(_06725_),
    .A2(_06720_),
    .ZN(_06726_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input53 (.I(key[31]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30826_ (.A1(net21258),
    .A2(_12816_),
    .A3(_12814_),
    .ZN(_06727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30827_ (.A1(net21007),
    .A2(net21001),
    .ZN(_06728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30828_ (.A1(net21383),
    .A2(net21331),
    .ZN(_06729_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30829_ (.A1(_06728_),
    .A2(net20966),
    .A3(_06729_),
    .ZN(_06730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30830_ (.A1(_06730_),
    .A2(_06727_),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30831_ (.A1(net20894),
    .A2(_06731_),
    .ZN(_06732_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30832_ (.A1(_06727_),
    .A2(_06730_),
    .A3(net20896),
    .ZN(_06733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30833_ (.A1(_06732_),
    .A2(_06733_),
    .B(net21486),
    .ZN(_06734_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30834_ (.I(\text_in_r[0] ),
    .ZN(_06735_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30835_ (.A1(_06735_),
    .A2(net21486),
    .Z(_06736_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30836_ (.A1(net20394),
    .A2(net20924),
    .B(net21155),
    .ZN(_06737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30837_ (.A1(_06732_),
    .A2(_06733_),
    .ZN(_06738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30838_ (.A1(_06738_),
    .A2(net21089),
    .ZN(_06739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30839_ (.I(net21155),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30840_ (.I(_06736_),
    .ZN(_06741_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30841_ (.A1(net20173),
    .A2(_06740_),
    .A3(_06741_),
    .ZN(_06742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30842_ (.A1(_06742_),
    .A2(_06737_),
    .ZN(_16178_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30843_ (.A1(net21269),
    .A2(net21325),
    .Z(_06743_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _30844_ (.A1(net21269),
    .A2(net21325),
    .ZN(_06744_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30845_ (.A1(_06743_),
    .A2(_06744_),
    .B(net21440),
    .ZN(_06745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30846_ (.A1(net21009),
    .A2(_12834_),
    .ZN(_06746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30847_ (.A1(net21270),
    .A2(net21325),
    .ZN(_06747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30848_ (.A1(_06746_),
    .A2(net20995),
    .A3(_06747_),
    .ZN(_06748_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30849_ (.A1(_06745_),
    .A2(_06748_),
    .ZN(_06749_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _30850_ (.A1(net21441),
    .A2(net21381),
    .ZN(_06750_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30851_ (.I(_06750_),
    .ZN(_06751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30852_ (.A1(_06749_),
    .A2(_06751_),
    .ZN(_06752_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30853_ (.A1(_06745_),
    .A2(_06748_),
    .A3(_06750_),
    .ZN(_06753_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30854_ (.A1(_06752_),
    .A2(_06753_),
    .B(net21486),
    .ZN(_06754_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30855_ (.I(\text_in_r[2] ),
    .ZN(_06755_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30856_ (.A1(_06755_),
    .A2(net21486),
    .Z(_06756_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30857_ (.A1(_06754_),
    .A2(_06756_),
    .B(net21139),
    .ZN(_06757_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30858_ (.A1(_06752_),
    .A2(_06753_),
    .ZN(_06758_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30859_ (.A1(_06758_),
    .A2(net21089),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30860_ (.I(_06756_),
    .ZN(_06760_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30861_ (.A1(_06759_),
    .A2(net21124),
    .A3(_06760_),
    .ZN(_06761_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30862_ (.A1(_06757_),
    .A2(_06761_),
    .ZN(_06762_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _30863_ (.I(_06762_),
    .ZN(_06763_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input52 (.I(key[30]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30865_ (.A1(_06736_),
    .A2(_06734_),
    .B(_06740_),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30866_ (.A1(_06739_),
    .A2(net21155),
    .A3(_06741_),
    .ZN(_06765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30867_ (.A1(_06765_),
    .A2(_06764_),
    .ZN(_16169_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input51 (.I(key[2]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30869_ (.A1(_06763_),
    .A2(net19457),
    .ZN(_06766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30870_ (.A1(net20890),
    .A2(net21323),
    .ZN(_06767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30871_ (.A1(net20889),
    .A2(net20992),
    .ZN(_06768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30872_ (.A1(_06767_),
    .A2(_06768_),
    .ZN(_06769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30873_ (.A1(net20405),
    .A2(_06769_),
    .ZN(_06770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30874_ (.A1(_06767_),
    .A2(_06768_),
    .Z(_06771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30875_ (.A1(net20404),
    .A2(_06771_),
    .ZN(_06772_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30876_ (.A1(_06770_),
    .A2(net21090),
    .A3(_06772_),
    .ZN(_06773_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30877_ (.I(net21138),
    .ZN(_06774_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _30878_ (.A1(net21090),
    .A2(\text_in_r[3] ),
    .Z(_06775_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30879_ (.A1(_06773_),
    .A2(_06774_),
    .A3(_06775_),
    .ZN(_06776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30880_ (.A1(net20405),
    .A2(_06771_),
    .ZN(_06777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30881_ (.A1(net20404),
    .A2(_06769_),
    .ZN(_06778_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30882_ (.A1(_06777_),
    .A2(net21090),
    .A3(_06778_),
    .ZN(_06779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30883_ (.A1(net21486),
    .A2(\text_in_r[3] ),
    .ZN(_06780_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30884_ (.A1(_06779_),
    .A2(net21138),
    .A3(_06780_),
    .ZN(_06781_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30885_ (.A1(_06776_),
    .A2(_06781_),
    .ZN(_06782_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input50 (.I(key[29]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30887_ (.A1(_06766_),
    .A2(net18985),
    .Z(_06784_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input49 (.I(key[28]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30889_ (.A1(net18999),
    .A2(net19465),
    .A3(net19458),
    .ZN(_06786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30890_ (.A1(_06784_),
    .A2(net18445),
    .ZN(_06787_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input48 (.I(key[27]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input47 (.I(key[26]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30893_ (.A1(net20170),
    .A2(net19922),
    .A3(net18358),
    .ZN(_06790_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _30894_ (.A1(net18988),
    .A2(_06790_),
    .Z(_06791_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30895_ (.A1(_12931_),
    .A2(_03869_),
    .B(net21090),
    .ZN(_06792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30896_ (.A1(_12931_),
    .A2(_03869_),
    .ZN(_06793_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30897_ (.I(_06793_),
    .ZN(_06794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30898_ (.A1(net21486),
    .A2(\text_in_r[4] ),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _30899_ (.A1(_06792_),
    .A2(_06794_),
    .B(_06795_),
    .ZN(_06796_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30900_ (.A1(_06796_),
    .A2(\u0.tmp_w[4] ),
    .ZN(_06797_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30901_ (.I(\u0.tmp_w[4] ),
    .ZN(_06798_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _30902_ (.A1(_06792_),
    .A2(_06794_),
    .B(_06798_),
    .C(_06795_),
    .ZN(_06799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30903_ (.A1(_06797_),
    .A2(_06799_),
    .ZN(_06800_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30904_ (.A1(_06791_),
    .A2(net19454),
    .Z(_06801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30905_ (.A1(_06787_),
    .A2(_06801_),
    .ZN(_06802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30906_ (.I(\u0.tmp_w[5] ),
    .ZN(_06803_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30907_ (.A1(net21263),
    .A2(\sa21_sub[5] ),
    .Z(_06804_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30908_ (.A1(_06804_),
    .A2(_00956_),
    .Z(_06805_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30909_ (.A1(_06804_),
    .A2(_00956_),
    .ZN(_06806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30910_ (.A1(_06805_),
    .A2(_06806_),
    .ZN(_06807_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _30911_ (.A1(net21437),
    .A2(\sa10_sub[5] ),
    .ZN(_06808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30912_ (.I(_06808_),
    .ZN(_06809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30913_ (.A1(_06807_),
    .A2(_06809_),
    .ZN(_06810_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30914_ (.A1(_06805_),
    .A2(_06808_),
    .A3(_06806_),
    .ZN(_06811_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30915_ (.A1(_06810_),
    .A2(_06811_),
    .A3(net21091),
    .ZN(_06812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30916_ (.A1(net21483),
    .A2(\text_in_r[5] ),
    .ZN(_06813_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30917_ (.A1(_06812_),
    .A2(_06813_),
    .ZN(_06814_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30918_ (.A1(_06803_),
    .A2(_06814_),
    .Z(_06815_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input46 (.I(key[25]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _30920_ (.I(_16172_[0]),
    .ZN(_06817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30921_ (.A1(net19459),
    .A2(_06817_),
    .ZN(_06818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30922_ (.A1(_06782_),
    .A2(_06818_),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30923_ (.I(_06800_),
    .ZN(_06820_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input45 (.I(key[24]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30925_ (.A1(_06819_),
    .A2(net18978),
    .Z(_06822_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30926_ (.A1(net19458),
    .A2(net18356),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30927_ (.A1(_06823_),
    .A2(_06790_),
    .ZN(_06824_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30928_ (.A1(_06779_),
    .A2(_06774_),
    .A3(_06780_),
    .ZN(_06825_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30929_ (.A1(_06773_),
    .A2(net21138),
    .A3(_06775_),
    .ZN(_06826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30930_ (.A1(_06825_),
    .A2(_06826_),
    .ZN(_06827_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input44 (.I(key[23]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30932_ (.A1(_06824_),
    .A2(net18966),
    .ZN(_06829_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30933_ (.A1(_06822_),
    .A2(_06829_),
    .ZN(_06830_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30934_ (.A1(_06802_),
    .A2(net20164),
    .A3(_06830_),
    .ZN(_06831_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _30935_ (.I(net415),
    .ZN(_06832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30936_ (.A1(_06832_),
    .A2(net19459),
    .ZN(_06833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30937_ (.A1(net18988),
    .A2(_06833_),
    .ZN(_06834_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30938_ (.A1(_06834_),
    .A2(net18978),
    .Z(_06835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30939_ (.A1(net19458),
    .A2(_16173_[0]),
    .ZN(_06836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30940_ (.I(_16171_[0]),
    .ZN(_06837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30941_ (.A1(net20170),
    .A2(net19923),
    .A3(_06837_),
    .ZN(_06838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30942_ (.A1(_06836_),
    .A2(_06838_),
    .ZN(_06839_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input43 (.I(key[22]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input42 (.I(key[21]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30945_ (.A1(_06839_),
    .A2(net18963),
    .ZN(_06842_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input41 (.I(key[20]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30947_ (.A1(_06835_),
    .A2(_06842_),
    .B(net20163),
    .ZN(_06844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30948_ (.A1(net19000),
    .A2(net19462),
    .ZN(_06845_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input40 (.I(key[1]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30950_ (.A1(net461),
    .A2(net19921),
    .A3(net20170),
    .ZN(_06847_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30951_ (.A1(_06845_),
    .A2(net18971),
    .A3(net18018),
    .ZN(_06848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30952_ (.A1(_06763_),
    .A2(_16179_[0]),
    .ZN(_06849_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input39 (.I(key[19]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30954_ (.A1(net19463),
    .A2(net19457),
    .ZN(_06851_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30955_ (.A1(net18017),
    .A2(net18991),
    .A3(_06851_),
    .ZN(_06852_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input38 (.I(key[18]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30957_ (.A1(_06848_),
    .A2(_06852_),
    .A3(net19448),
    .ZN(_06854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30958_ (.A1(_06844_),
    .A2(_06854_),
    .ZN(_06855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30959_ (.A1(_06831_),
    .A2(_06855_),
    .ZN(_06856_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _30960_ (.A1(net21262),
    .A2(\sa21_sub[6] ),
    .A3(\sa03_sr[6] ),
    .Z(_06857_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30961_ (.A1(\sa03_sr[5] ),
    .A2(net21376),
    .Z(_06858_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30962_ (.A1(_06857_),
    .A2(_06858_),
    .Z(_06859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30963_ (.A1(_06857_),
    .A2(_06858_),
    .ZN(_06860_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30964_ (.A1(_06859_),
    .A2(net21092),
    .A3(_06860_),
    .ZN(_06861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30965_ (.A1(net21492),
    .A2(\text_in_r[6] ),
    .ZN(_06862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30966_ (.A1(_06861_),
    .A2(_06862_),
    .Z(_06863_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _30967_ (.A1(_06863_),
    .A2(\u0.tmp_w[6] ),
    .Z(_06864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30968_ (.A1(_06863_),
    .A2(\u0.tmp_w[6] ),
    .ZN(_06865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30969_ (.A1(_06864_),
    .A2(_06865_),
    .ZN(_06866_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input37 (.I(key[17]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30971_ (.A1(_06856_),
    .A2(net20391),
    .ZN(_06868_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _30972_ (.A1(net21261),
    .A2(net20892),
    .A3(net20988),
    .ZN(_06869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _30973_ (.A1(net21489),
    .A2(\text_in_r[7] ),
    .Z(_06870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _30974_ (.A1(_06869_),
    .A2(net21092),
    .B(_06870_),
    .ZN(_06871_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _30975_ (.A1(\u0.tmp_w[7] ),
    .A2(_06871_),
    .Z(_06872_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input36 (.I(key[16]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30977_ (.I(_06872_),
    .ZN(_06874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30978_ (.A1(_06868_),
    .A2(_06874_),
    .ZN(_06875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30979_ (.A1(_06849_),
    .A2(net18967),
    .ZN(_06876_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _30980_ (.I(_06876_),
    .ZN(_06877_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30981_ (.A1(net18999),
    .A2(net19457),
    .A3(net19463),
    .ZN(_06878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30982_ (.A1(_06877_),
    .A2(net18443),
    .ZN(_06879_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input35 (.I(key[15]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _30984_ (.I(_06836_),
    .ZN(_06881_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input34 (.I(key[14]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30986_ (.A1(_06881_),
    .A2(net18986),
    .ZN(_06883_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30987_ (.A1(_06879_),
    .A2(net18978),
    .A3(_06883_),
    .ZN(_06884_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30988_ (.A1(_06881_),
    .A2(net18969),
    .ZN(_06885_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30989_ (.A1(_06885_),
    .A2(net19447),
    .Z(_06886_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _30990_ (.I(_16181_[0]),
    .ZN(_06887_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _30991_ (.A1(_06887_),
    .A2(net19923),
    .A3(net20172),
    .ZN(_06888_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _30992_ (.A1(net18985),
    .A2(_06888_),
    .Z(_06889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30993_ (.A1(net18443),
    .A2(_06889_),
    .ZN(_06890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _30994_ (.A1(_06886_),
    .A2(_06890_),
    .ZN(_06891_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _30995_ (.I(_06815_),
    .ZN(_06892_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input33 (.I(key[13]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input32 (.I(key[12]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _30998_ (.A1(_06884_),
    .A2(_06891_),
    .A3(net19918),
    .ZN(_06895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _30999_ (.A1(net19458),
    .A2(_06837_),
    .ZN(_06896_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31000_ (.A1(_06896_),
    .A2(net18971),
    .B(net19450),
    .ZN(_06897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31001_ (.A1(_06763_),
    .A2(net19465),
    .ZN(_06898_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31002_ (.A1(_06898_),
    .A2(net18971),
    .ZN(_06899_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31003_ (.A1(_06897_),
    .A2(_06899_),
    .ZN(_06900_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input31 (.I(net585),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31005_ (.A1(net20171),
    .A2(net19922),
    .A3(_06832_),
    .ZN(_06902_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31006_ (.A1(_06878_),
    .A2(net18971),
    .A3(_06902_),
    .ZN(_06903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31007_ (.A1(net18995),
    .A2(net18359),
    .Z(_06904_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input30 (.I(net546),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31009_ (.A1(_06904_),
    .A2(net18963),
    .ZN(_06906_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31010_ (.A1(_06900_),
    .A2(_06903_),
    .A3(_06906_),
    .ZN(_06907_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31011_ (.A1(_06847_),
    .A2(_06827_),
    .Z(_06908_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31012_ (.A1(net18970),
    .A2(_16192_[0]),
    .ZN(_06909_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31013_ (.A1(_06908_),
    .A2(_06909_),
    .Z(_06910_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input29 (.I(net565),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input28 (.I(net588),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31016_ (.A1(net18981),
    .A2(_06910_),
    .B(net19914),
    .ZN(_06913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31017_ (.A1(_06907_),
    .A2(_06913_),
    .ZN(_06914_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31018_ (.A1(_06914_),
    .A2(_06895_),
    .B(net20391),
    .ZN(_06915_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31019_ (.A1(_06875_),
    .A2(_06915_),
    .ZN(_06916_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31020_ (.A1(_06717_),
    .A2(net21147),
    .A3(_06719_),
    .ZN(_06917_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31021_ (.A1(_06723_),
    .A2(_06718_),
    .A3(_06724_),
    .ZN(_06918_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31022_ (.A1(_06918_),
    .A2(_06917_),
    .ZN(_16170_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31023_ (.A1(net519),
    .A2(net18995),
    .Z(_06919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31024_ (.A1(_06919_),
    .A2(_06881_),
    .B(net18961),
    .ZN(_06920_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input27 (.I(net536),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31026_ (.A1(_06787_),
    .A2(_06920_),
    .A3(net19454),
    .ZN(_06922_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31027_ (.A1(net19462),
    .A2(net18355),
    .ZN(_06923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31028_ (.A1(_06898_),
    .A2(_06923_),
    .ZN(_06924_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input26 (.I(net539),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input25 (.I(net538),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31031_ (.A1(_06924_),
    .A2(net18994),
    .B(net19448),
    .ZN(_06927_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31032_ (.A1(_06762_),
    .A2(net19465),
    .ZN(_06928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31033_ (.A1(_06928_),
    .A2(net18999),
    .ZN(_06929_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input24 (.I(net537),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31035_ (.A1(net19462),
    .A2(net519),
    .ZN(_06931_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input23 (.I(key[11]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31037_ (.A1(net18439),
    .A2(net18977),
    .A3(_06931_),
    .ZN(_06933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31038_ (.A1(_06927_),
    .A2(_06933_),
    .ZN(_06934_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input22 (.I(key[119]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31040_ (.A1(_06922_),
    .A2(_06934_),
    .A3(net20167),
    .ZN(_06936_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _31041_ (.I(_06834_),
    .ZN(_06937_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31042_ (.A1(_06937_),
    .A2(net18438),
    .ZN(_06938_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31043_ (.A1(_06766_),
    .A2(net18971),
    .Z(_06939_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31044_ (.I(_06939_),
    .ZN(_06940_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input21 (.I(key[118]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31046_ (.A1(_06938_),
    .A2(_06940_),
    .A3(net19448),
    .ZN(_06942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31047_ (.A1(net18360),
    .A2(net19460),
    .ZN(_06943_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31048_ (.A1(net20172),
    .A2(net19923),
    .A3(net18355),
    .ZN(_06944_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31049_ (.A1(_06943_),
    .A2(_06944_),
    .ZN(_06945_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input20 (.I(net540),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31051_ (.A1(net17620),
    .A2(net18991),
    .B(net19448),
    .ZN(_06947_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31052_ (.A1(_06929_),
    .A2(net18970),
    .A3(_06851_),
    .ZN(_06948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31053_ (.A1(_06947_),
    .A2(_06948_),
    .ZN(_06949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31054_ (.A1(_06942_),
    .A2(_06949_),
    .A3(net19915),
    .ZN(_06950_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _31055_ (.I(_06866_),
    .ZN(_06951_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input19 (.I(key[116]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31057_ (.A1(_06936_),
    .A2(_06950_),
    .B(_06951_),
    .ZN(_06953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _31058_ (.I(_06819_),
    .ZN(_06954_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31059_ (.A1(net20172),
    .A2(net19923),
    .A3(net18361),
    .ZN(_06955_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31060_ (.A1(_06954_),
    .A2(net18014),
    .ZN(_06956_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _31061_ (.I(_06896_),
    .ZN(_06957_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31062_ (.A1(net19458),
    .A2(_16179_[0]),
    .ZN(_06958_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31063_ (.A1(net17363),
    .A2(net18012),
    .B(net18972),
    .ZN(_06959_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input18 (.I(key[115]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31065_ (.A1(_06956_),
    .A2(_06959_),
    .B(net18981),
    .ZN(_06961_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31066_ (.A1(net20171),
    .A2(net439),
    .A3(net19922),
    .ZN(_06962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31067_ (.A1(net18985),
    .A2(_06962_),
    .Z(_06963_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31068_ (.A1(_06963_),
    .A2(net19448),
    .ZN(_06964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31069_ (.A1(net19001),
    .A2(net18996),
    .ZN(_06965_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31070_ (.A1(_06965_),
    .A2(net18970),
    .A3(_06943_),
    .ZN(_06966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31071_ (.A1(_06964_),
    .A2(_06966_),
    .ZN(_06967_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input17 (.I(key[114]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31073_ (.A1(_06967_),
    .A2(net20167),
    .ZN(_06969_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31074_ (.A1(_06969_),
    .A2(_06961_),
    .B(_06951_),
    .ZN(_06970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31075_ (.A1(net19462),
    .A2(net19465),
    .ZN(_06971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31076_ (.A1(_06971_),
    .A2(net18961),
    .Z(_06972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31077_ (.A1(net519),
    .A2(net19457),
    .ZN(_06973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31078_ (.A1(_06972_),
    .A2(_06973_),
    .ZN(_06974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31079_ (.A1(net18999),
    .A2(net19457),
    .ZN(_06975_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31080_ (.A1(_06975_),
    .A2(_06898_),
    .A3(net18994),
    .ZN(_06976_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31081_ (.A1(_06974_),
    .A2(_06976_),
    .A3(net18982),
    .ZN(_06977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31082_ (.A1(net17631),
    .A2(net18961),
    .ZN(_06978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31083_ (.I(_06978_),
    .ZN(_06979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31084_ (.A1(net19000),
    .A2(_06763_),
    .A3(net19465),
    .ZN(_06980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31085_ (.A1(_06979_),
    .A2(net18432),
    .ZN(_06981_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input16 (.I(key[113]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31087_ (.I(_16179_[0]),
    .ZN(_06983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31088_ (.A1(net19462),
    .A2(_06983_),
    .ZN(_06984_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31089_ (.A1(_06984_),
    .A2(net17627),
    .ZN(_06985_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input15 (.I(key[112]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31091_ (.A1(_06985_),
    .A2(net18994),
    .ZN(_06987_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31092_ (.A1(_06981_),
    .A2(net19449),
    .A3(_06987_),
    .ZN(_06988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31093_ (.A1(_06977_),
    .A2(_06988_),
    .B(net20169),
    .ZN(_06989_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31094_ (.A1(_06970_),
    .A2(_06989_),
    .B(net20389),
    .ZN(_06990_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31095_ (.A1(_06990_),
    .A2(_06953_),
    .ZN(_06991_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _31096_ (.A1(_06916_),
    .A2(_06991_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31097_ (.A1(_06975_),
    .A2(net18997),
    .ZN(_06992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31098_ (.A1(net18999),
    .A2(net19465),
    .ZN(_06993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31099_ (.A1(_06993_),
    .A2(net19462),
    .ZN(_06994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31100_ (.A1(_06992_),
    .A2(_06994_),
    .Z(_06995_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31101_ (.A1(_06851_),
    .A2(net18970),
    .A3(_06955_),
    .ZN(_06996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31102_ (.A1(_06996_),
    .A2(_06892_),
    .Z(_06997_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31103_ (.A1(net18977),
    .A2(_06995_),
    .B(_06997_),
    .ZN(_06998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31104_ (.A1(_06972_),
    .A2(_06965_),
    .ZN(_06999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31105_ (.A1(_06763_),
    .A2(net519),
    .ZN(_07000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31106_ (.A1(_06937_),
    .A2(_07000_),
    .ZN(_07001_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31107_ (.A1(_06999_),
    .A2(_07001_),
    .A3(net20163),
    .ZN(_07002_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31108_ (.A1(_06998_),
    .A2(net18983),
    .A3(_07002_),
    .ZN(_07003_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31109_ (.A1(_06892_),
    .A2(_16195_[0]),
    .A3(net18971),
    .Z(_07004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31110_ (.A1(_06877_),
    .A2(net476),
    .ZN(_07005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31111_ (.A1(_07004_),
    .A2(_07005_),
    .ZN(_07006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31112_ (.A1(_07006_),
    .A2(net19451),
    .B(net20391),
    .ZN(_07007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31113_ (.A1(_07007_),
    .A2(_07003_),
    .B(_06874_),
    .ZN(_07008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31114_ (.A1(_06786_),
    .A2(net18961),
    .ZN(_07009_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31115_ (.A1(_07009_),
    .A2(net18957),
    .B(net19454),
    .C(net17367),
    .ZN(_07010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31116_ (.A1(_06980_),
    .A2(net18991),
    .ZN(_07011_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _31117_ (.I(_06943_),
    .ZN(_07012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _31118_ (.A1(_07011_),
    .A2(_07012_),
    .Z(_07013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _31119_ (.I(_16185_[0]),
    .ZN(_07014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31120_ (.A1(net19458),
    .A2(_07014_),
    .ZN(_07015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31121_ (.A1(_07015_),
    .A2(net18961),
    .Z(_07016_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _31122_ (.I(_16173_[0]),
    .ZN(_07017_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31123_ (.A1(net20171),
    .A2(_07017_),
    .A3(net19922),
    .ZN(_07018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31124_ (.A1(net17362),
    .A2(net17615),
    .B(net19454),
    .ZN(_07019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31125_ (.A1(_07013_),
    .A2(_07019_),
    .ZN(_07020_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31126_ (.A1(_07010_),
    .A2(_07020_),
    .A3(net20168),
    .ZN(_07021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31127_ (.A1(_06957_),
    .A2(net18987),
    .ZN(_07022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31128_ (.A1(_06885_),
    .A2(_07022_),
    .Z(_07023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31129_ (.I(_06898_),
    .ZN(_07024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31130_ (.A1(_07024_),
    .A2(net18969),
    .B(net19447),
    .ZN(_07025_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31131_ (.I(_06847_),
    .ZN(_07026_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31132_ (.A1(_07026_),
    .A2(net18989),
    .ZN(_07027_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31133_ (.A1(_07023_),
    .A2(_07025_),
    .A3(net17361),
    .ZN(_07028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31134_ (.A1(_06972_),
    .A2(net18014),
    .ZN(_07029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31135_ (.A1(_07029_),
    .A2(_07001_),
    .A3(net19451),
    .ZN(_07030_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31136_ (.A1(_07028_),
    .A2(net19919),
    .A3(_07030_),
    .ZN(_07031_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31137_ (.A1(_07021_),
    .A2(_07031_),
    .A3(net20392),
    .ZN(_07032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31138_ (.A1(_07008_),
    .A2(_07032_),
    .ZN(_07033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31139_ (.A1(net18992),
    .A2(net19462),
    .ZN(_07034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31140_ (.A1(net18992),
    .A2(net519),
    .ZN(_07035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31141_ (.A1(_07034_),
    .A2(_07035_),
    .ZN(_07036_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31142_ (.A1(_07036_),
    .A2(net19454),
    .ZN(_07037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31143_ (.A1(_06791_),
    .A2(net521),
    .Z(_07038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31144_ (.A1(_07037_),
    .A2(_07038_),
    .B(net19918),
    .ZN(_07039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31145_ (.A1(_06963_),
    .A2(net17616),
    .ZN(_07040_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31146_ (.A1(_06903_),
    .A2(_07040_),
    .A3(net19450),
    .ZN(_07041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31147_ (.A1(_07039_),
    .A2(_07041_),
    .B(net20391),
    .ZN(_07042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31148_ (.A1(_06898_),
    .A2(net18968),
    .Z(_07043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31149_ (.A1(_07043_),
    .A2(net17628),
    .ZN(_07044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31150_ (.A1(net18022),
    .A2(net393),
    .ZN(_07045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31151_ (.A1(_07044_),
    .A2(_07045_),
    .A3(net18978),
    .ZN(_07046_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31152_ (.A1(_06845_),
    .A2(_06973_),
    .A3(net18970),
    .ZN(_07047_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31153_ (.A1(net18992),
    .A2(_06763_),
    .Z(_07048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31154_ (.A1(_07048_),
    .A2(_06975_),
    .ZN(_07049_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31155_ (.A1(_07047_),
    .A2(net19447),
    .A3(_07049_),
    .ZN(_07050_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31156_ (.A1(_07046_),
    .A2(_07050_),
    .A3(net19918),
    .ZN(_07051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31157_ (.A1(_07042_),
    .A2(_07051_),
    .B(net20390),
    .ZN(_07052_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _31158_ (.A1(_07014_),
    .A2(net20172),
    .A3(net19923),
    .ZN(_07053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31159_ (.A1(_07053_),
    .A2(net18985),
    .Z(_07054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31160_ (.A1(_07054_),
    .A2(_06931_),
    .ZN(_07055_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31161_ (.A1(net18991),
    .A2(net18010),
    .B(_07055_),
    .C(net18981),
    .ZN(_07056_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31162_ (.A1(net18962),
    .A2(net18357),
    .Z(_07057_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input14 (.I(net581),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31164_ (.A1(_07057_),
    .A2(net19461),
    .B(net18978),
    .ZN(_07059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31165_ (.A1(_07013_),
    .A2(_07059_),
    .ZN(_07060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31166_ (.A1(_07056_),
    .A2(_07060_),
    .A3(net19913),
    .ZN(_07061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31167_ (.A1(_07043_),
    .A2(net17623),
    .ZN(_07062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31168_ (.A1(_06954_),
    .A2(net18021),
    .ZN(_07063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31169_ (.A1(_07062_),
    .A2(_07063_),
    .ZN(_07064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31170_ (.A1(_07064_),
    .A2(net18978),
    .ZN(_07065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31171_ (.I(_06993_),
    .ZN(_07066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31172_ (.I(_06851_),
    .ZN(_07067_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31173_ (.A1(_07066_),
    .A2(_07067_),
    .B(net18993),
    .ZN(_07068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31174_ (.A1(net17621),
    .A2(_06851_),
    .ZN(_07069_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31175_ (.A1(_07068_),
    .A2(net19448),
    .A3(_07069_),
    .ZN(_07070_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31176_ (.A1(_07065_),
    .A2(_07070_),
    .A3(net20165),
    .ZN(_07071_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31177_ (.A1(_07061_),
    .A2(_07071_),
    .A3(net20391),
    .ZN(_07072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31178_ (.A1(_07072_),
    .A2(_07052_),
    .ZN(_07073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31179_ (.A1(_07033_),
    .A2(_07073_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31180_ (.A1(net18439),
    .A2(net18975),
    .B(net18981),
    .ZN(_07074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31181_ (.A1(net18432),
    .A2(net18994),
    .A3(net17616),
    .ZN(_07075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31182_ (.A1(_07074_),
    .A2(_07075_),
    .B(net20167),
    .ZN(_07076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31183_ (.A1(net19464),
    .A2(net19465),
    .Z(_07077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31184_ (.A1(_06904_),
    .A2(_07077_),
    .B(net18990),
    .ZN(_07078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31185_ (.A1(net18434),
    .A2(net18977),
    .A3(net17632),
    .ZN(_07079_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31186_ (.A1(_07078_),
    .A2(_07079_),
    .A3(net18982),
    .ZN(_07080_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31187_ (.A1(_07076_),
    .A2(_07080_),
    .B(net20391),
    .ZN(_07081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31188_ (.A1(_06845_),
    .A2(_06975_),
    .A3(net18994),
    .ZN(_07082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31189_ (.I(_07082_),
    .ZN(_07083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31190_ (.A1(_06833_),
    .A2(net18967),
    .ZN(_07084_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31191_ (.I(_07053_),
    .ZN(_07085_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31192_ (.A1(_07085_),
    .A2(_07084_),
    .ZN(_07086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31193_ (.A1(_07083_),
    .A2(_07086_),
    .B(net18981),
    .ZN(_07087_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31194_ (.A1(_06851_),
    .A2(_06902_),
    .ZN(_07088_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31195_ (.A1(_07088_),
    .A2(net18991),
    .A3(net521),
    .ZN(_07089_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31196_ (.A1(_07089_),
    .A2(net19452),
    .A3(_06848_),
    .ZN(_07090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31197_ (.A1(_07087_),
    .A2(_07090_),
    .ZN(_07091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31198_ (.A1(_07091_),
    .A2(net20166),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31199_ (.A1(_07081_),
    .A2(_07092_),
    .ZN(_07093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31200_ (.A1(net18429),
    .A2(net18991),
    .A3(net18020),
    .ZN(_07094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31201_ (.A1(net18956),
    .A2(net18973),
    .A3(_06944_),
    .ZN(_07095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31202_ (.A1(_07094_),
    .A2(net18981),
    .A3(_07095_),
    .ZN(_07096_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31203_ (.A1(_06851_),
    .A2(net18971),
    .A3(net17625),
    .ZN(_07097_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31204_ (.A1(net17632),
    .A2(net18018),
    .A3(net18991),
    .ZN(_07098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31205_ (.A1(_07097_),
    .A2(_07098_),
    .ZN(_07099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31206_ (.A1(_07099_),
    .A2(net19452),
    .ZN(_07100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31207_ (.A1(_07096_),
    .A2(_07100_),
    .ZN(_07101_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31208_ (.A1(_07101_),
    .A2(net19918),
    .ZN(_07102_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31209_ (.A1(net18436),
    .A2(net18991),
    .A3(net17622),
    .ZN(_07103_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31210_ (.A1(_07103_),
    .A2(net17366),
    .A3(net19453),
    .ZN(_07104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31211_ (.A1(net18020),
    .A2(net18015),
    .ZN(_07105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31212_ (.A1(_07105_),
    .A2(net18974),
    .ZN(_07106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31213_ (.A1(net18960),
    .A2(net18991),
    .A3(net17622),
    .ZN(_07107_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31214_ (.A1(_07106_),
    .A2(_07107_),
    .A3(net18983),
    .ZN(_07108_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31215_ (.A1(_07104_),
    .A2(_07108_),
    .A3(net20166),
    .ZN(_07109_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31216_ (.A1(_07102_),
    .A2(_07109_),
    .A3(net20391),
    .ZN(_07110_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31217_ (.A1(_07093_),
    .A2(net20390),
    .A3(_07110_),
    .ZN(_07111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31218_ (.A1(_06984_),
    .A2(net18994),
    .Z(_07112_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31219_ (.A1(_07112_),
    .A2(net18018),
    .Z(_07113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31220_ (.A1(_06845_),
    .A2(net18970),
    .ZN(_07114_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31221_ (.I(_06838_),
    .ZN(_07115_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31222_ (.A1(_07114_),
    .A2(_07115_),
    .ZN(_07116_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31223_ (.A1(_07113_),
    .A2(_07116_),
    .B(net18982),
    .ZN(_07117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31224_ (.A1(_06845_),
    .A2(_06973_),
    .A3(net18994),
    .ZN(_07118_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31225_ (.A1(_07118_),
    .A2(net19448),
    .Z(_07119_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31226_ (.A1(net18994),
    .A2(_16195_[0]),
    .Z(_07120_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31227_ (.A1(_07119_),
    .A2(_07120_),
    .ZN(_07121_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31228_ (.A1(_07117_),
    .A2(_07121_),
    .A3(net20167),
    .ZN(_07122_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31229_ (.A1(_07000_),
    .A2(net18991),
    .Z(_07123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31230_ (.A1(_07123_),
    .A2(net18960),
    .ZN(_07124_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31231_ (.A1(_07124_),
    .A2(net18981),
    .A3(_06848_),
    .ZN(_07125_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input13 (.I(net553),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31233_ (.A1(net18354),
    .A2(net18975),
    .B(net18981),
    .ZN(_07127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31234_ (.A1(net18444),
    .A2(net474),
    .ZN(_07128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31235_ (.A1(_07128_),
    .A2(_07127_),
    .B(net20166),
    .ZN(_07129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31236_ (.A1(_07125_),
    .A2(_07129_),
    .B(_06951_),
    .ZN(_07130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31237_ (.A1(_07130_),
    .A2(_07122_),
    .ZN(_07131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31238_ (.A1(_07000_),
    .A2(_06766_),
    .ZN(_07132_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31239_ (.I(_07132_),
    .ZN(_07133_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31240_ (.A1(_07017_),
    .A2(_06832_),
    .ZN(_07134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31241_ (.A1(net19461),
    .A2(net17613),
    .ZN(_07135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31242_ (.A1(_07133_),
    .A2(_07135_),
    .ZN(_07136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31243_ (.A1(_07136_),
    .A2(net18991),
    .ZN(_07137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31244_ (.A1(net17365),
    .A2(net18446),
    .B(net19451),
    .ZN(_07138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31245_ (.A1(_07137_),
    .A2(_07138_),
    .ZN(_07139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31246_ (.A1(_06957_),
    .A2(net18971),
    .ZN(_07140_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31247_ (.A1(_07140_),
    .A2(net19453),
    .Z(_07141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31248_ (.A1(_06954_),
    .A2(net17622),
    .ZN(_07142_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31249_ (.A1(_07142_),
    .A2(_07141_),
    .B(net20166),
    .ZN(_07143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31250_ (.A1(_07139_),
    .A2(_07143_),
    .ZN(_07144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31251_ (.A1(net392),
    .A2(net18971),
    .ZN(_07145_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31252_ (.A1(net18971),
    .A2(_16190_[0]),
    .Z(_07146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31253_ (.A1(_07145_),
    .A2(_07146_),
    .ZN(_07147_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31254_ (.A1(_07147_),
    .A2(net18981),
    .Z(_07148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31255_ (.A1(_16199_[0]),
    .A2(net18977),
    .B(net19448),
    .ZN(_07149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31256_ (.A1(_07082_),
    .A2(_07149_),
    .B(net19916),
    .ZN(_07150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31257_ (.A1(_07148_),
    .A2(_07150_),
    .ZN(_07151_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31258_ (.A1(_07144_),
    .A2(_07151_),
    .A3(_06951_),
    .ZN(_07152_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31259_ (.A1(net20162),
    .A2(_07152_),
    .A3(_07131_),
    .ZN(_07153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31260_ (.A1(_07153_),
    .A2(_07111_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31261_ (.A1(_06900_),
    .A2(_07047_),
    .ZN(_07154_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _31262_ (.I(_06823_),
    .ZN(_07155_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _31263_ (.A1(_07155_),
    .A2(net18957),
    .B(net18988),
    .ZN(_07156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31264_ (.A1(_06945_),
    .A2(net18972),
    .ZN(_07157_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31265_ (.A1(_07156_),
    .A2(net18978),
    .A3(_07157_),
    .ZN(_07158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31266_ (.A1(_07154_),
    .A2(_07158_),
    .ZN(_07159_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31267_ (.A1(_07159_),
    .A2(net19920),
    .ZN(_07160_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _31268_ (.A1(net18996),
    .A2(_07134_),
    .B(_06888_),
    .C(net18991),
    .ZN(_07161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31269_ (.A1(_07005_),
    .A2(_07161_),
    .ZN(_07162_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31270_ (.A1(_07162_),
    .A2(net19451),
    .ZN(_07163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31271_ (.A1(_07095_),
    .A2(net18983),
    .B(net19920),
    .ZN(_07164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31272_ (.A1(_07163_),
    .A2(_07164_),
    .ZN(_07165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31273_ (.A1(_07160_),
    .A2(_07165_),
    .A3(net20391),
    .ZN(_07166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31274_ (.A1(_06939_),
    .A2(net393),
    .ZN(_07167_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31275_ (.A1(net18996),
    .A2(_07134_),
    .B(net17614),
    .C(net18991),
    .ZN(_07168_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31276_ (.A1(_07167_),
    .A2(_07168_),
    .A3(net20163),
    .ZN(_07169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31277_ (.A1(_07155_),
    .A2(net18986),
    .ZN(_07170_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31278_ (.A1(_07097_),
    .A2(_07170_),
    .A3(net19920),
    .ZN(_07171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31279_ (.A1(_07169_),
    .A2(_07171_),
    .ZN(_07172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31280_ (.A1(_07172_),
    .A2(net19451),
    .ZN(_07173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _31281_ (.I(net17632),
    .ZN(_07174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31282_ (.A1(net18975),
    .A2(_07174_),
    .ZN(_07175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31283_ (.I(_07175_),
    .ZN(_07176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31284_ (.A1(_06883_),
    .A2(net18978),
    .ZN(_07177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31285_ (.A1(_07176_),
    .A2(net19919),
    .B(_07177_),
    .ZN(_07178_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31286_ (.I(_06845_),
    .ZN(_07179_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31287_ (.A1(_06876_),
    .A2(_07179_),
    .ZN(_07180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _31288_ (.I(_06962_),
    .ZN(_07181_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31289_ (.A1(_07181_),
    .A2(net18986),
    .Z(_07182_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31290_ (.A1(_07180_),
    .A2(_07182_),
    .B(net20163),
    .ZN(_07183_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31291_ (.A1(_07178_),
    .A2(_07183_),
    .B(net20391),
    .ZN(_07184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31292_ (.A1(_07184_),
    .A2(_07173_),
    .ZN(_07185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31293_ (.A1(_07166_),
    .A2(_07185_),
    .ZN(_07186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31294_ (.A1(_07186_),
    .A2(net20390),
    .ZN(_07187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31295_ (.I(_07182_),
    .ZN(_07188_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31296_ (.A1(_07188_),
    .A2(net20163),
    .A3(_06999_),
    .ZN(_07189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31297_ (.A1(net473),
    .A2(net17624),
    .ZN(_07190_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31298_ (.A1(net18442),
    .A2(net18976),
    .A3(net17618),
    .ZN(_07191_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31299_ (.A1(_07190_),
    .A2(_07191_),
    .A3(net19918),
    .ZN(_07192_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31300_ (.A1(_07189_),
    .A2(_07192_),
    .ZN(_07193_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31301_ (.A1(net18983),
    .A2(_07193_),
    .ZN(_07194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31302_ (.A1(_06972_),
    .A2(net18433),
    .ZN(_07195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31303_ (.A1(_06954_),
    .A2(net18429),
    .ZN(_07196_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31304_ (.A1(_07195_),
    .A2(_07196_),
    .A3(net20166),
    .ZN(_07197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31305_ (.A1(_06943_),
    .A2(net18970),
    .Z(_07198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31306_ (.A1(_07198_),
    .A2(net18429),
    .ZN(_07199_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31307_ (.A1(net17616),
    .A2(net17622),
    .A3(net18991),
    .ZN(_07200_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31308_ (.A1(_07199_),
    .A2(net19918),
    .A3(_07200_),
    .ZN(_07201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31309_ (.A1(_07197_),
    .A2(_07201_),
    .A3(net19453),
    .ZN(_07202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31310_ (.A1(_06951_),
    .A2(_07194_),
    .A3(_07202_),
    .ZN(_07203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31311_ (.A1(_07198_),
    .A2(net17625),
    .ZN(_07204_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31312_ (.A1(_07204_),
    .A2(_07055_),
    .A3(net18981),
    .ZN(_07205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31313_ (.A1(net18428),
    .A2(net19448),
    .Z(_07206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31314_ (.A1(_06975_),
    .A2(_06971_),
    .ZN(_07207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31315_ (.A1(_07206_),
    .A2(net18005),
    .B(net19916),
    .ZN(_07208_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31316_ (.A1(_07205_),
    .A2(_07208_),
    .B(_06951_),
    .ZN(_07209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31317_ (.A1(_06992_),
    .A2(_07112_),
    .ZN(_07210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31318_ (.A1(_06994_),
    .A2(net477),
    .ZN(_07211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31319_ (.A1(_07210_),
    .A2(_07211_),
    .A3(net19448),
    .ZN(_07212_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31320_ (.A1(_06978_),
    .A2(net18013),
    .Z(_07213_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31321_ (.A1(_07213_),
    .A2(_06976_),
    .A3(net18982),
    .ZN(_07214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31322_ (.A1(_07212_),
    .A2(_07214_),
    .ZN(_07215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31323_ (.A1(_07215_),
    .A2(net19918),
    .ZN(_07216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31324_ (.A1(_07209_),
    .A2(_07216_),
    .ZN(_07217_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31325_ (.A1(net20162),
    .A2(_07217_),
    .A3(_07203_),
    .ZN(_07218_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31326_ (.A1(_07218_),
    .A2(_07187_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31327_ (.A1(_07048_),
    .A2(net19000),
    .Z(_07219_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31328_ (.A1(_07219_),
    .A2(_06897_),
    .ZN(_07220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31329_ (.A1(_07220_),
    .A2(_06903_),
    .ZN(_07221_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31330_ (.A1(_07086_),
    .A2(net19452),
    .ZN(_07222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31331_ (.A1(net18008),
    .A2(net18444),
    .ZN(_07223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31332_ (.A1(_07222_),
    .A2(_07223_),
    .ZN(_07224_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31333_ (.A1(_07221_),
    .A2(net20166),
    .A3(_07224_),
    .ZN(_07225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31334_ (.A1(_07027_),
    .A2(net18978),
    .Z(_07226_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31335_ (.A1(_07226_),
    .A2(_06829_),
    .A3(_07170_),
    .ZN(_07227_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31336_ (.A1(net17362),
    .A2(net17619),
    .ZN(_07228_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31337_ (.A1(_07228_),
    .A2(_06890_),
    .A3(net19447),
    .ZN(_07229_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31338_ (.A1(_07227_),
    .A2(_07229_),
    .A3(net19919),
    .ZN(_07230_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31339_ (.A1(_07225_),
    .A2(_07230_),
    .A3(_06951_),
    .ZN(_07231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31340_ (.A1(_06999_),
    .A2(_07118_),
    .A3(net19448),
    .ZN(_07233_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31341_ (.A1(net521),
    .A2(net18431),
    .A3(net18977),
    .ZN(_07234_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31342_ (.A1(net18437),
    .A2(net18994),
    .A3(net18014),
    .ZN(_07235_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31343_ (.A1(_07234_),
    .A2(_07235_),
    .A3(net18981),
    .ZN(_07236_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31344_ (.A1(_07233_),
    .A2(_07236_),
    .A3(net20167),
    .ZN(_07237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31345_ (.A1(_07036_),
    .A2(_06851_),
    .ZN(_07238_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31346_ (.A1(_07238_),
    .A2(net19449),
    .A3(net17617),
    .ZN(_07239_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31347_ (.A1(net18978),
    .A2(net18019),
    .Z(_07240_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31348_ (.I(net17364),
    .ZN(_07241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31349_ (.A1(_07240_),
    .A2(_07241_),
    .B(net20163),
    .ZN(_07242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31350_ (.A1(_07239_),
    .A2(_07242_),
    .ZN(_07244_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31351_ (.A1(_07244_),
    .A2(net20391),
    .A3(_07237_),
    .ZN(_07245_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31352_ (.A1(_07231_),
    .A2(_07245_),
    .A3(net20162),
    .ZN(_07246_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31353_ (.A1(net18433),
    .A2(net19461),
    .A3(net18976),
    .ZN(_07247_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31354_ (.A1(_06889_),
    .A2(_06931_),
    .ZN(_07248_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31355_ (.A1(_07247_),
    .A2(_07248_),
    .B(net19447),
    .ZN(_07249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31356_ (.A1(net18961),
    .A2(_16183_[0]),
    .ZN(_07250_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31357_ (.A1(_07027_),
    .A2(net19454),
    .A3(_07250_),
    .Z(_07251_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31358_ (.A1(_07249_),
    .A2(_07251_),
    .B(net19918),
    .ZN(_07252_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31359_ (.A1(_07000_),
    .A2(_06975_),
    .A3(net18965),
    .ZN(_07253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31360_ (.A1(_06889_),
    .A2(net18956),
    .ZN(_07255_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31361_ (.A1(_07253_),
    .A2(_07255_),
    .A3(net18980),
    .ZN(_07256_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31362_ (.A1(_06976_),
    .A2(net19454),
    .A3(_06842_),
    .ZN(_07257_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31363_ (.A1(_07256_),
    .A2(_07257_),
    .A3(net20169),
    .ZN(_07258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31364_ (.A1(_07252_),
    .A2(_07258_),
    .A3(_06951_),
    .ZN(_07259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31365_ (.A1(net18429),
    .A2(net17624),
    .ZN(_07260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31366_ (.A1(_07260_),
    .A2(net18971),
    .ZN(_07261_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31367_ (.A1(_07261_),
    .A2(_07001_),
    .A3(net18983),
    .ZN(_07262_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31368_ (.A1(_06972_),
    .A2(net17614),
    .ZN(_07263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31369_ (.I(net18426),
    .ZN(_07264_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31370_ (.A1(_07263_),
    .A2(net19448),
    .A3(_07264_),
    .ZN(_07266_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31371_ (.A1(_07262_),
    .A2(_07266_),
    .A3(net20166),
    .ZN(_07267_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31372_ (.A1(net17621),
    .A2(net17628),
    .ZN(_07268_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31373_ (.A1(_06787_),
    .A2(net19447),
    .A3(_07268_),
    .ZN(_07269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31374_ (.A1(_07018_),
    .A2(net18970),
    .ZN(_07270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31375_ (.A1(_07270_),
    .A2(net18978),
    .Z(_07271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31376_ (.A1(_07271_),
    .A2(_07011_),
    .B(net20168),
    .ZN(_07272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31377_ (.A1(_07269_),
    .A2(_07272_),
    .ZN(_07273_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31378_ (.A1(_07267_),
    .A2(net20391),
    .A3(_07273_),
    .ZN(_07274_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31379_ (.A1(_07259_),
    .A2(_07274_),
    .A3(net20390),
    .ZN(_07275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31380_ (.A1(_07246_),
    .A2(_07275_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31381_ (.A1(net519),
    .A2(net19464),
    .B(net18961),
    .ZN(_07277_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31382_ (.A1(_07067_),
    .A2(net18013),
    .ZN(_07278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31383_ (.A1(_07277_),
    .A2(_07278_),
    .ZN(_07279_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31384_ (.A1(net18430),
    .A2(_06766_),
    .A3(net18964),
    .ZN(_07280_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31385_ (.A1(_07279_),
    .A2(net18978),
    .A3(_07280_),
    .ZN(_07281_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31386_ (.A1(_07253_),
    .A2(net19454),
    .A3(net18427),
    .ZN(_07282_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31387_ (.A1(_07281_),
    .A2(_07282_),
    .A3(net19913),
    .ZN(_07283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31388_ (.A1(_07179_),
    .A2(_07270_),
    .ZN(_07284_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31389_ (.I(_07027_),
    .ZN(_07285_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31390_ (.A1(_07284_),
    .A2(_07285_),
    .B(net18979),
    .ZN(_07287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31391_ (.A1(_06944_),
    .A2(net18970),
    .ZN(_07288_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31392_ (.A1(net17367),
    .A2(_07115_),
    .B(net19454),
    .C(_07288_),
    .ZN(_07289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31393_ (.A1(_07287_),
    .A2(_07289_),
    .A3(net20164),
    .ZN(_07290_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31394_ (.A1(_07283_),
    .A2(_06951_),
    .A3(_07290_),
    .ZN(_07291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31395_ (.A1(net18988),
    .A2(net18357),
    .ZN(_07292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31396_ (.A1(_07292_),
    .A2(net18978),
    .ZN(_07293_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31397_ (.A1(_06836_),
    .A2(net18961),
    .ZN(_07294_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31398_ (.A1(_07293_),
    .A2(_07294_),
    .ZN(_07295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31399_ (.A1(_06888_),
    .A2(net18967),
    .Z(_07296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31400_ (.A1(net18443),
    .A2(_07296_),
    .ZN(_07298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31401_ (.A1(_07295_),
    .A2(_07298_),
    .B(net20163),
    .ZN(_07299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31402_ (.A1(_07054_),
    .A2(net17628),
    .ZN(_07300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31403_ (.A1(_06920_),
    .A2(_07300_),
    .A3(net19454),
    .ZN(_07301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31404_ (.A1(_07299_),
    .A2(_07301_),
    .ZN(_07302_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31405_ (.A1(_07084_),
    .A2(net18978),
    .Z(_07303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31406_ (.A1(_07303_),
    .A2(_07049_),
    .B(_06892_),
    .ZN(_07304_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31407_ (.A1(_07156_),
    .A2(net19454),
    .A3(_06978_),
    .ZN(_07305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31408_ (.A1(_07304_),
    .A2(_07305_),
    .ZN(_07306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31409_ (.A1(_07302_),
    .A2(_07306_),
    .ZN(_07307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31410_ (.A1(_07307_),
    .A2(net20393),
    .ZN(_07309_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31411_ (.A1(_07291_),
    .A2(_07309_),
    .ZN(_07310_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31412_ (.A1(_07310_),
    .A2(net20161),
    .ZN(_07311_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31413_ (.A1(net18986),
    .A2(net17359),
    .B(_06787_),
    .C(net19454),
    .ZN(_07312_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31414_ (.A1(_07009_),
    .A2(_07085_),
    .Z(_07313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31415_ (.A1(net18012),
    .A2(net18986),
    .B(net19454),
    .ZN(_07314_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31416_ (.A1(_07313_),
    .A2(_07314_),
    .B(net19913),
    .ZN(_07315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31417_ (.A1(_07312_),
    .A2(_07315_),
    .ZN(_07316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31418_ (.A1(net19465),
    .A2(net18990),
    .B(net18978),
    .ZN(_07317_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31419_ (.A1(_07317_),
    .A2(_06974_),
    .B(net20169),
    .ZN(_07318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31420_ (.A1(_06954_),
    .A2(net18438),
    .ZN(_07320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31421_ (.A1(_07296_),
    .A2(net521),
    .ZN(_07321_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31422_ (.A1(_07320_),
    .A2(_07321_),
    .A3(net18984),
    .ZN(_07322_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31423_ (.A1(_07318_),
    .A2(_07322_),
    .B(_06951_),
    .ZN(_07323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31424_ (.A1(_07323_),
    .A2(_07316_),
    .ZN(_07324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31425_ (.A1(_06791_),
    .A2(net18978),
    .Z(_07325_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31426_ (.I(net17360),
    .ZN(_07326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31427_ (.A1(_07325_),
    .A2(_07326_),
    .B(net20164),
    .ZN(_07327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31428_ (.A1(net18990),
    .A2(net18359),
    .ZN(_07328_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31429_ (.A1(_06834_),
    .A2(net19454),
    .A3(_07328_),
    .Z(_07329_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31430_ (.A1(net18438),
    .A2(net18445),
    .A3(net18970),
    .ZN(_07331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31431_ (.A1(_07329_),
    .A2(_07331_),
    .ZN(_07332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31432_ (.A1(_07327_),
    .A2(_07332_),
    .ZN(_07333_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31433_ (.A1(net18011),
    .A2(net18988),
    .B(net18979),
    .ZN(_07334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31434_ (.A1(_07334_),
    .A2(net18009),
    .B(net19913),
    .ZN(_07335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31435_ (.A1(_07198_),
    .A2(net17614),
    .ZN(_07336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31436_ (.A1(net18017),
    .A2(_06954_),
    .ZN(_07337_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31437_ (.A1(_07337_),
    .A2(_07336_),
    .A3(net18978),
    .ZN(_07338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31438_ (.A1(_07335_),
    .A2(_07338_),
    .ZN(_07339_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31439_ (.A1(_07333_),
    .A2(_06951_),
    .A3(_07339_),
    .ZN(_07340_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31440_ (.A1(_07340_),
    .A2(_07324_),
    .A3(net20389),
    .ZN(_07342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31441_ (.A1(_07342_),
    .A2(_07311_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31442_ (.A1(_07054_),
    .A2(net18016),
    .ZN(_07343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31443_ (.A1(_07025_),
    .A2(_07343_),
    .ZN(_07344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31444_ (.I(_16189_[0]),
    .ZN(_07345_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31445_ (.A1(_07345_),
    .A2(net18990),
    .B(net18978),
    .ZN(_07346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31446_ (.A1(_07346_),
    .A2(_07321_),
    .ZN(_07347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31447_ (.A1(_07344_),
    .A2(_07347_),
    .ZN(_07348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31448_ (.A1(_07348_),
    .A2(net19919),
    .B(net20391),
    .ZN(_07349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31449_ (.A1(_07248_),
    .A2(net17626),
    .Z(_07350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31450_ (.A1(_07089_),
    .A2(net19451),
    .ZN(_07351_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31451_ (.A1(net19447),
    .A2(_07350_),
    .B(_07351_),
    .C(net20163),
    .ZN(_07352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31452_ (.A1(_07349_),
    .A2(_07352_),
    .ZN(_07353_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31453_ (.A1(_07037_),
    .A2(_06948_),
    .ZN(_07354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31454_ (.A1(_07012_),
    .A2(net18970),
    .B(net18978),
    .ZN(_07355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31455_ (.A1(_07355_),
    .A2(_07156_),
    .ZN(_07356_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31456_ (.A1(_07354_),
    .A2(_07356_),
    .A3(net20169),
    .ZN(_07357_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31457_ (.A1(net519),
    .A2(net18961),
    .B(net18978),
    .ZN(_07358_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31458_ (.A1(_07358_),
    .A2(_07207_),
    .B(net20163),
    .ZN(_07359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31459_ (.A1(_07207_),
    .A2(net18990),
    .ZN(_07360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31460_ (.A1(_07016_),
    .A2(net18441),
    .ZN(_07362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31461_ (.A1(_07360_),
    .A2(_07362_),
    .A3(net18978),
    .ZN(_07363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31462_ (.A1(_07359_),
    .A2(_07363_),
    .ZN(_07364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31463_ (.A1(_07357_),
    .A2(_07364_),
    .ZN(_07365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31464_ (.A1(_07365_),
    .A2(net20392),
    .ZN(_07366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31465_ (.A1(_07353_),
    .A2(_07366_),
    .ZN(_07367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31466_ (.A1(_07367_),
    .A2(net20390),
    .ZN(_07368_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31467_ (.A1(_16188_[0]),
    .A2(_16197_[0]),
    .Z(_07369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31468_ (.A1(net18961),
    .A2(_07369_),
    .B(net20163),
    .ZN(_07370_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31469_ (.A1(_07000_),
    .A2(_06975_),
    .A3(net18990),
    .ZN(_07371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31470_ (.A1(_07370_),
    .A2(_07371_),
    .B(net18980),
    .ZN(_07373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31471_ (.A1(net18006),
    .A2(net18986),
    .B(net17611),
    .ZN(_07374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31472_ (.A1(_07296_),
    .A2(net17616),
    .B(_06892_),
    .ZN(_07375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31473_ (.A1(_07374_),
    .A2(_07375_),
    .ZN(_07376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31474_ (.A1(_07373_),
    .A2(_07376_),
    .B(_06951_),
    .ZN(_07377_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31475_ (.A1(net17621),
    .A2(net18956),
    .A3(net20163),
    .ZN(_07378_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31476_ (.A1(net17629),
    .A2(net18986),
    .A3(net20163),
    .ZN(_07379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31477_ (.A1(_06904_),
    .A2(net18986),
    .ZN(_07380_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31478_ (.A1(_07378_),
    .A2(_07379_),
    .A3(_07380_),
    .ZN(_07381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31479_ (.A1(_07140_),
    .A2(_07170_),
    .B(net20165),
    .ZN(_07382_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31480_ (.A1(_07381_),
    .A2(_07382_),
    .B(net18978),
    .ZN(_07384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31481_ (.A1(_07377_),
    .A2(_07384_),
    .B(net20390),
    .ZN(_07385_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _31482_ (.A1(_07147_),
    .A2(net18981),
    .A3(_07175_),
    .Z(_07386_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31483_ (.A1(net18439),
    .A2(net18994),
    .A3(net521),
    .ZN(_07387_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31484_ (.A1(_07270_),
    .A2(_07012_),
    .Z(_07388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31485_ (.A1(_07387_),
    .A2(_07388_),
    .B(net18978),
    .ZN(_07389_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31486_ (.A1(_07386_),
    .A2(_07389_),
    .B(net19913),
    .ZN(_07390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31487_ (.A1(_06878_),
    .A2(net18991),
    .ZN(_07391_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31488_ (.A1(_07391_),
    .A2(_07024_),
    .Z(_07392_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31489_ (.A1(_07392_),
    .A2(_06886_),
    .A3(_07268_),
    .ZN(_07393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31490_ (.A1(net18012),
    .A2(net18966),
    .B(net19447),
    .ZN(_07395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31491_ (.A1(_06971_),
    .A2(net19001),
    .ZN(_07396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31492_ (.A1(_07396_),
    .A2(net18986),
    .ZN(_07397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31493_ (.A1(_07395_),
    .A2(_07397_),
    .B(net19917),
    .ZN(_07398_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31494_ (.A1(_07393_),
    .A2(_07398_),
    .B(net20391),
    .ZN(_07399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31495_ (.A1(_07390_),
    .A2(_07399_),
    .ZN(_07400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31496_ (.A1(_07385_),
    .A2(_07400_),
    .ZN(_07401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31497_ (.A1(_07368_),
    .A2(_07401_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31498_ (.A1(_07114_),
    .A2(_07066_),
    .B(_07161_),
    .ZN(_07402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31499_ (.A1(_07402_),
    .A2(net18978),
    .ZN(_07403_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31500_ (.A1(_07133_),
    .A2(net18971),
    .A3(net17623),
    .ZN(_07405_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31501_ (.A1(net18012),
    .A2(_06819_),
    .Z(_07406_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31502_ (.A1(_07405_),
    .A2(net19454),
    .A3(_07406_),
    .ZN(_07407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31503_ (.A1(_07403_),
    .A2(_07407_),
    .ZN(_07408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31504_ (.A1(_07408_),
    .A2(net19913),
    .ZN(_07409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31505_ (.A1(net18440),
    .A2(net18990),
    .ZN(_07410_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _31506_ (.A1(net19454),
    .A2(_07410_),
    .A3(_06906_),
    .A4(net17623),
    .ZN(_07411_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31507_ (.A1(_07057_),
    .A2(net19454),
    .ZN(_07412_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31508_ (.A1(_07371_),
    .A2(_07412_),
    .B(net19913),
    .ZN(_07413_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31509_ (.A1(_07411_),
    .A2(_07413_),
    .B(_06951_),
    .ZN(_07414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31510_ (.A1(_07409_),
    .A2(_07414_),
    .ZN(_07416_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31511_ (.I(_16183_[0]),
    .ZN(_07417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31512_ (.A1(_07417_),
    .A2(net18990),
    .B(net18978),
    .ZN(_07418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _31513_ (.A1(_07418_),
    .A2(_06906_),
    .B(net20163),
    .ZN(_07419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31514_ (.A1(_07396_),
    .A2(net18969),
    .ZN(_07420_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31515_ (.A1(_07001_),
    .A2(net18984),
    .A3(_07420_),
    .ZN(_07421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31516_ (.A1(_07419_),
    .A2(_07421_),
    .B(net20391),
    .ZN(_07422_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31517_ (.A1(_07181_),
    .A2(net18968),
    .A3(_07012_),
    .Z(_07423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31518_ (.A1(_06939_),
    .A2(net18435),
    .ZN(_07424_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31519_ (.A1(net18984),
    .A2(_07424_),
    .A3(_07423_),
    .ZN(_07425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31520_ (.A1(net18353),
    .A2(net18990),
    .B(net18978),
    .ZN(_07427_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31521_ (.A1(net17612),
    .A2(net440),
    .B(net18969),
    .ZN(_07428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31522_ (.A1(_07427_),
    .A2(_07428_),
    .B(net19918),
    .ZN(_07429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31523_ (.A1(_07429_),
    .A2(_07425_),
    .ZN(_07430_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31524_ (.A1(_07430_),
    .A2(_07422_),
    .B(net20389),
    .ZN(_07431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31525_ (.A1(_07431_),
    .A2(_07416_),
    .ZN(_07432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31526_ (.A1(_07375_),
    .A2(_07124_),
    .ZN(_07433_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31527_ (.A1(_07016_),
    .A2(net20163),
    .ZN(_07434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31528_ (.A1(_07434_),
    .A2(_07248_),
    .B(net18978),
    .ZN(_07435_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31529_ (.A1(_07433_),
    .A2(_07435_),
    .B(_06951_),
    .ZN(_07436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31530_ (.A1(_07022_),
    .A2(_06892_),
    .Z(_07438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31531_ (.A1(_06939_),
    .A2(net18443),
    .ZN(_07439_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31532_ (.A1(net18007),
    .A2(net18986),
    .ZN(_07440_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31533_ (.A1(_07438_),
    .A2(_07439_),
    .A3(_07440_),
    .ZN(_07441_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31534_ (.A1(_07040_),
    .A2(net20163),
    .A3(_07167_),
    .ZN(_07442_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31535_ (.A1(_07442_),
    .A2(_07441_),
    .A3(net18978),
    .ZN(_07443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31536_ (.A1(_07436_),
    .A2(_07443_),
    .B(_06874_),
    .ZN(_07444_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31537_ (.A1(net18432),
    .A2(net18975),
    .A3(net18437),
    .ZN(_07445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31538_ (.A1(_07119_),
    .A2(_07445_),
    .ZN(_07446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31539_ (.A1(net18965),
    .A2(net19457),
    .ZN(_07447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31540_ (.A1(_07238_),
    .A2(_07447_),
    .ZN(_07449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31541_ (.A1(_07449_),
    .A2(net18982),
    .ZN(_07450_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31542_ (.A1(_07446_),
    .A2(_07450_),
    .A3(net19916),
    .ZN(_07451_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _31543_ (.A1(net18010),
    .A2(net18975),
    .B(_07175_),
    .C(net19448),
    .ZN(_07452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31544_ (.A1(_07198_),
    .A2(net18432),
    .ZN(_07453_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31545_ (.A1(_07453_),
    .A2(_07391_),
    .A3(net18981),
    .ZN(_07454_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31546_ (.A1(_07452_),
    .A2(_07454_),
    .A3(net20167),
    .ZN(_07455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31547_ (.A1(_07451_),
    .A2(_07455_),
    .A3(_06951_),
    .ZN(_07456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31548_ (.A1(_07456_),
    .A2(_07444_),
    .ZN(_07457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31549_ (.A1(_07432_),
    .A2(_07457_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31550_ (.I(\dcnt[3] ),
    .ZN(_07459_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31551_ (.I(\dcnt[2] ),
    .ZN(_07460_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31552_ (.A1(_07459_),
    .A2(_07460_),
    .Z(_07461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31553_ (.I(\dcnt[1] ),
    .ZN(_07462_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _31554_ (.A1(_07461_),
    .A2(net21521),
    .A3(_07462_),
    .A4(\dcnt[0] ),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31555_ (.A1(net21223),
    .A2(net21480),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31556_ (.A1(net21222),
    .A2(net21478),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31557_ (.A1(net21221),
    .A2(net21475),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31558_ (.A1(net21220),
    .A2(net21474),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31559_ (.A1(net21219),
    .A2(net21473),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31560_ (.A1(net21218),
    .A2(\sa00_sr[5] ),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31561_ (.A1(net21216),
    .A2(\sa00_sr[6] ),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31562_ (.A1(net21215),
    .A2(net21470),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31563_ (.A1(net21195),
    .A2(net21467),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31564_ (.A1(net21194),
    .A2(net21466),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31565_ (.A1(net21193),
    .A2(net21463),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31566_ (.A1(net21192),
    .A2(net21462),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31567_ (.A1(net21191),
    .A2(net21461),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31568_ (.A1(net21190),
    .A2(net21460),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31569_ (.A1(\u0.w[1][30] ),
    .A2(\sa01_sr[6] ),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31570_ (.A1(\u0.w[1][31] ),
    .A2(net21459),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31571_ (.A1(net21169),
    .A2(net21455),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31572_ (.A1(net21168),
    .A2(net21453),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31573_ (.A1(net21167),
    .A2(net21451),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31574_ (.A1(net21166),
    .A2(net21450),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31575_ (.A1(net21165),
    .A2(net21448),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31576_ (.A1(net21164),
    .A2(\sa02_sr[5] ),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31577_ (.A1(net21162),
    .A2(net21447),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31578_ (.A1(net21161),
    .A2(net21445),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31579_ (.A1(net21145),
    .A2(net21443),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31580_ (.A1(net21144),
    .A2(net21441),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31581_ (.A1(net21143),
    .A2(net21440),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31582_ (.A1(net21142),
    .A2(net21439),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31583_ (.A1(net21141),
    .A2(net21437),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31584_ (.A1(net21140),
    .A2(\sa03_sr[5] ),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31585_ (.A1(\u0.tmp_w[30] ),
    .A2(\sa03_sr[6] ),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31586_ (.A1(\u0.tmp_w[31] ),
    .A2(net21435),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31587_ (.A1(net21230),
    .A2(net21431),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31588_ (.A1(net21229),
    .A2(net21426),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31589_ (.A1(net21228),
    .A2(net21422),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31590_ (.A1(net21227),
    .A2(net21419),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31591_ (.A1(net21225),
    .A2(net21418),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31592_ (.A1(net21224),
    .A2(net21417),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31593_ (.A1(\u0.w[0][22] ),
    .A2(\sa10_sr[6] ),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31594_ (.A1(\u0.w[0][23] ),
    .A2(net21414),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31595_ (.A1(net21203),
    .A2(net21412),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31596_ (.A1(net21202),
    .A2(net21409),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31597_ (.A1(net21201),
    .A2(net21408),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31598_ (.A1(net21200),
    .A2(net21407),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31599_ (.A1(net21198),
    .A2(net21406),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31600_ (.A1(net21197),
    .A2(net21405),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31601_ (.A1(net21196),
    .A2(net21404),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31602_ (.A1(\u0.w[1][23] ),
    .A2(net21403),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31603_ (.A1(net21176),
    .A2(net21399),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31604_ (.A1(net21175),
    .A2(net21397),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31605_ (.A1(net21174),
    .A2(net21394),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31606_ (.A1(net21173),
    .A2(net21391),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31607_ (.A1(net21171),
    .A2(net21390),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31608_ (.A1(net21170),
    .A2(\sa12_sr[5] ),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31609_ (.A1(\u0.w[2][22] ),
    .A2(net21389),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31610_ (.A1(\u0.w[2][23] ),
    .A2(net21385),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31611_ (.A1(net21151),
    .A2(\sa10_sub[0] ),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31612_ (.A1(net21150),
    .A2(net21382),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31613_ (.A1(net21149),
    .A2(net21381),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31614_ (.A1(net21148),
    .A2(\sa10_sub[3] ),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31615_ (.A1(net21146),
    .A2(net21378),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31616_ (.A1(\u0.tmp_w[21] ),
    .A2(net21377),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31617_ (.A1(\u0.tmp_w[22] ),
    .A2(net21376),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31618_ (.A1(\u0.tmp_w[23] ),
    .A2(net21373),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31619_ (.A1(net21211),
    .A2(net21369),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31620_ (.A1(net21209),
    .A2(net21368),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31621_ (.A1(net21235),
    .A2(net21367),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31622_ (.A1(net21234),
    .A2(net21366),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31623_ (.A1(net21233),
    .A2(net21364),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31624_ (.A1(net21232),
    .A2(\sa20_sr[5] ),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31625_ (.A1(net21231),
    .A2(\sa20_sr[6] ),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31626_ (.A1(\u0.w[0][15] ),
    .A2(net21362),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31627_ (.A1(net21183),
    .A2(\sa21_sr[0] ),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31628_ (.A1(net21182),
    .A2(net21357),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31629_ (.A1(net21207),
    .A2(net21354),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31630_ (.A1(net21206),
    .A2(net21352),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31631_ (.A1(net21205),
    .A2(net21351),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31632_ (.A1(net21204),
    .A2(net21350),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31633_ (.A1(\u0.w[1][14] ),
    .A2(net21349),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31634_ (.A1(\u0.w[1][15] ),
    .A2(net443),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31635_ (.A1(net21157),
    .A2(net21344),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31636_ (.A1(net21156),
    .A2(net21342),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31637_ (.A1(net21180),
    .A2(\sa20_sub[2] ),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31638_ (.A1(net21179),
    .A2(net21338),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31639_ (.A1(net21178),
    .A2(net21337),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31640_ (.A1(net21177),
    .A2(net21336),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31641_ (.A1(\u0.w[2][14] ),
    .A2(net21335),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31642_ (.A1(\u0.w[2][15] ),
    .A2(net21332),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31643_ (.A1(net21137),
    .A2(net21329),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31644_ (.A1(net21136),
    .A2(net21326),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31645_ (.A1(net21154),
    .A2(net21324),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31646_ (.A1(net21153),
    .A2(net21321),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31647_ (.A1(net21152),
    .A2(net21320),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31648_ (.A1(\u0.tmp_w[13] ),
    .A2(net21317),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31649_ (.A1(\u0.tmp_w[14] ),
    .A2(\sa21_sub[6] ),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31650_ (.A1(\u0.tmp_w[15] ),
    .A2(net21315),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31651_ (.A1(net21236),
    .A2(net21313),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31652_ (.A1(net21226),
    .A2(net21311),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31653_ (.A1(net21217),
    .A2(net21308),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31654_ (.A1(net21214),
    .A2(net21306),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31655_ (.A1(net21213),
    .A2(net21303),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31656_ (.A1(net21212),
    .A2(net21301),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31657_ (.A1(\u0.w[0][6] ),
    .A2(\sa30_sr[6] ),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31658_ (.A1(\u0.w[0][7] ),
    .A2(net21298),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31659_ (.A1(net21208),
    .A2(net21297),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31660_ (.A1(net21199),
    .A2(net21296),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31661_ (.A1(net21189),
    .A2(net21294),
    .Z(_00251_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31662_ (.A1(net21188),
    .A2(net21291),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31663_ (.A1(net21187),
    .A2(net21290),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31664_ (.A1(net21186),
    .A2(net21289),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31665_ (.A1(net21185),
    .A2(net21288),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31666_ (.A1(net21184),
    .A2(net21285),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31667_ (.A1(net21181),
    .A2(net21284),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31668_ (.A1(net21172),
    .A2(net21283),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31669_ (.A1(net21163),
    .A2(net21281),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31670_ (.A1(net21160),
    .A2(net21279),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31671_ (.A1(net21159),
    .A2(net21278),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31672_ (.A1(net21158),
    .A2(net21277),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31673_ (.A1(\u0.w[2][6] ),
    .A2(net21276),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31674_ (.A1(\u0.w[2][7] ),
    .A2(net21275),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31675_ (.A1(net21155),
    .A2(\sa32_sub[0] ),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31676_ (.A1(net21147),
    .A2(\sa32_sub[1] ),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31677_ (.A1(net21139),
    .A2(net21267),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31678_ (.A1(net21138),
    .A2(net21266),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31679_ (.A1(\u0.tmp_w[4] ),
    .A2(net21264),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31680_ (.A1(\u0.tmp_w[5] ),
    .A2(net21262),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31681_ (.A1(\u0.tmp_w[6] ),
    .A2(net21261),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31682_ (.A1(\u0.tmp_w[7] ),
    .A2(net21258),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31683_ (.I(\u0.r0.rcnt[0] ),
    .ZN(\u0.r0.rcnt_next[0] ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31684_ (.I(\u0.r0.rcnt[1] ),
    .ZN(_16201_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31685_ (.I0(\text_in_r[0] ),
    .I1(net131),
    .S(net21539),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(key[10]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31687_ (.I0(\text_in_r[100] ),
    .I1(net132),
    .S(net21537),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31688_ (.I0(\text_in_r[101] ),
    .I1(net133),
    .S(net21535),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31689_ (.I0(\text_in_r[102] ),
    .I1(net134),
    .S(net21539),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31690_ (.I0(\text_in_r[103] ),
    .I1(net135),
    .S(net21535),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31691_ (.I0(\text_in_r[104] ),
    .I1(net136),
    .S(net21537),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31692_ (.I0(\text_in_r[105] ),
    .I1(net137),
    .S(net21537),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31693_ (.I0(\text_in_r[106] ),
    .I1(net138),
    .S(net21537),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31694_ (.I0(\text_in_r[107] ),
    .I1(net139),
    .S(net21537),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31695_ (.I0(\text_in_r[108] ),
    .I1(net140),
    .S(net21535),
    .Z(_00418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31696_ (.I0(\text_in_r[109] ),
    .I1(net141),
    .S(net21539),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input11 (.I(net562),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31698_ (.I0(\text_in_r[10] ),
    .I1(net142),
    .S(net21532),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31699_ (.I0(\text_in_r[110] ),
    .I1(net143),
    .S(net21539),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31700_ (.I0(\text_in_r[111] ),
    .I1(net144),
    .S(net21535),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31701_ (.I0(\text_in_r[112] ),
    .I1(net145),
    .S(net21535),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31702_ (.I0(\text_in_r[113] ),
    .I1(net146),
    .S(net21540),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31703_ (.I0(\text_in_r[114] ),
    .I1(net147),
    .S(net21539),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31704_ (.I0(\text_in_r[115] ),
    .I1(net148),
    .S(net21540),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31705_ (.I0(\text_in_r[116] ),
    .I1(net149),
    .S(net21541),
    .Z(_00427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31706_ (.I0(\text_in_r[117] ),
    .I1(net150),
    .S(net21539),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31707_ (.I0(\text_in_r[118] ),
    .I1(net151),
    .S(net21539),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input10 (.I(key[108]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31709_ (.I0(\text_in_r[119] ),
    .I1(net152),
    .S(net21535),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31710_ (.I0(\text_in_r[11] ),
    .I1(net153),
    .S(net21539),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31711_ (.I0(\text_in_r[120] ),
    .I1(net154),
    .S(net21535),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31712_ (.I0(\text_in_r[121] ),
    .I1(net155),
    .S(net21535),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31713_ (.I0(\text_in_r[122] ),
    .I1(net156),
    .S(net21535),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31714_ (.I0(\text_in_r[123] ),
    .I1(net157),
    .S(net21535),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31715_ (.I0(\text_in_r[124] ),
    .I1(net158),
    .S(net21535),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31716_ (.I0(\text_in_r[125] ),
    .I1(net159),
    .S(net21539),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31717_ (.I0(\text_in_r[126] ),
    .I1(net160),
    .S(net21535),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31718_ (.I0(\text_in_r[127] ),
    .I1(net161),
    .S(net21535),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input9 (.I(key[107]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31720_ (.I0(\text_in_r[12] ),
    .I1(net162),
    .S(net21534),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31721_ (.I0(\text_in_r[13] ),
    .I1(net163),
    .S(net21543),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31722_ (.I0(\text_in_r[14] ),
    .I1(net164),
    .S(net21539),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31723_ (.I0(\text_in_r[15] ),
    .I1(net165),
    .S(net21539),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31724_ (.I0(\text_in_r[16] ),
    .I1(net166),
    .S(net21539),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31725_ (.I0(\text_in_r[17] ),
    .I1(net167),
    .S(net21539),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31726_ (.I0(\text_in_r[18] ),
    .I1(net168),
    .S(net21539),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31727_ (.I0(\text_in_r[19] ),
    .I1(net169),
    .S(net21539),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31728_ (.I0(\text_in_r[1] ),
    .I1(net170),
    .S(net21539),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31729_ (.I0(\text_in_r[20] ),
    .I1(net171),
    .S(net21539),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input8 (.I(key[106]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31731_ (.I0(\text_in_r[21] ),
    .I1(net172),
    .S(net21541),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31732_ (.I0(\text_in_r[22] ),
    .I1(net173),
    .S(net21541),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31733_ (.I0(\text_in_r[23] ),
    .I1(net174),
    .S(net21541),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31734_ (.I0(\text_in_r[24] ),
    .I1(net175),
    .S(net21539),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31735_ (.I0(\text_in_r[25] ),
    .I1(net176),
    .S(net21541),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31736_ (.I0(\text_in_r[26] ),
    .I1(net177),
    .S(net21541),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31737_ (.I0(\text_in_r[27] ),
    .I1(net178),
    .S(net21541),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31738_ (.I0(\text_in_r[28] ),
    .I1(net179),
    .S(net21541),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31739_ (.I0(\text_in_r[29] ),
    .I1(net180),
    .S(net21541),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31740_ (.I0(\text_in_r[2] ),
    .I1(net181),
    .S(net21539),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(key[105]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31742_ (.I0(\text_in_r[30] ),
    .I1(net182),
    .S(net21541),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31743_ (.I0(\text_in_r[31] ),
    .I1(net183),
    .S(net21541),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31744_ (.I0(\text_in_r[32] ),
    .I1(net184),
    .S(net21535),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31745_ (.I0(\text_in_r[33] ),
    .I1(net185),
    .S(net21535),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31746_ (.I0(\text_in_r[34] ),
    .I1(net186),
    .S(net21535),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31747_ (.I0(\text_in_r[35] ),
    .I1(net187),
    .S(net21535),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31748_ (.I0(\text_in_r[36] ),
    .I1(net188),
    .S(net21535),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31749_ (.I0(\text_in_r[37] ),
    .I1(net189),
    .S(net21535),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31750_ (.I0(\text_in_r[38] ),
    .I1(net190),
    .S(net21535),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31751_ (.I0(\text_in_r[39] ),
    .I1(net191),
    .S(net21535),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input6 (.I(key[104]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31753_ (.I0(\text_in_r[3] ),
    .I1(net192),
    .S(net21539),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31754_ (.I0(\text_in_r[40] ),
    .I1(net193),
    .S(net21535),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31755_ (.I0(\text_in_r[41] ),
    .I1(net194),
    .S(net21535),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31756_ (.I0(\text_in_r[42] ),
    .I1(net195),
    .S(net21535),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31757_ (.I0(\text_in_r[43] ),
    .I1(net196),
    .S(net21535),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31758_ (.I0(\text_in_r[44] ),
    .I1(net197),
    .S(net21535),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31759_ (.I0(\text_in_r[45] ),
    .I1(net198),
    .S(net21535),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31760_ (.I0(\text_in_r[46] ),
    .I1(net199),
    .S(net21535),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31761_ (.I0(\text_in_r[47] ),
    .I1(net200),
    .S(net21535),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31762_ (.I0(\text_in_r[48] ),
    .I1(net201),
    .S(net21535),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input5 (.I(net566),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31764_ (.I0(\text_in_r[49] ),
    .I1(net202),
    .S(net21537),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31765_ (.I0(\text_in_r[4] ),
    .I1(net203),
    .S(net21539),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31766_ (.I0(\text_in_r[50] ),
    .I1(net204),
    .S(net21537),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31767_ (.I0(\text_in_r[51] ),
    .I1(net205),
    .S(net21537),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31768_ (.I0(\text_in_r[52] ),
    .I1(net206),
    .S(net21537),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31769_ (.I0(\text_in_r[53] ),
    .I1(net207),
    .S(net21535),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31770_ (.I0(\text_in_r[54] ),
    .I1(net208),
    .S(net21535),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31771_ (.I0(\text_in_r[55] ),
    .I1(net209),
    .S(net21537),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31772_ (.I0(\text_in_r[56] ),
    .I1(net210),
    .S(net21535),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31773_ (.I0(\text_in_r[57] ),
    .I1(net211),
    .S(net21535),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input4 (.I(key[102]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31775_ (.I0(\text_in_r[58] ),
    .I1(net212),
    .S(net21535),
    .Z(_00490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31776_ (.I0(\text_in_r[59] ),
    .I1(net213),
    .S(net21535),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31777_ (.I0(\text_in_r[5] ),
    .I1(net214),
    .S(net21539),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31778_ (.I0(\text_in_r[60] ),
    .I1(net215),
    .S(net21535),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31779_ (.I0(\text_in_r[61] ),
    .I1(net216),
    .S(net21535),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31780_ (.I0(\text_in_r[62] ),
    .I1(net217),
    .S(net21535),
    .Z(_00495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31781_ (.I0(\text_in_r[63] ),
    .I1(net218),
    .S(net21535),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31782_ (.I0(\text_in_r[64] ),
    .I1(net219),
    .S(net21535),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31783_ (.I0(\text_in_r[65] ),
    .I1(net220),
    .S(net21535),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31784_ (.I0(\text_in_r[66] ),
    .I1(net221),
    .S(net21537),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input3 (.I(key[101]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31786_ (.I0(\text_in_r[67] ),
    .I1(net222),
    .S(net21535),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31787_ (.I0(\text_in_r[68] ),
    .I1(net223),
    .S(net21535),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31788_ (.I0(\text_in_r[69] ),
    .I1(net224),
    .S(net21537),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31789_ (.I0(\text_in_r[6] ),
    .I1(net225),
    .S(net21539),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31790_ (.I0(\text_in_r[70] ),
    .I1(net226),
    .S(net21535),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31791_ (.I0(\text_in_r[71] ),
    .I1(net227),
    .S(net21537),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31792_ (.I0(\text_in_r[72] ),
    .I1(net228),
    .S(net21534),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31793_ (.I0(\text_in_r[73] ),
    .I1(net229),
    .S(net21534),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31794_ (.I0(\text_in_r[74] ),
    .I1(net230),
    .S(net21534),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31795_ (.I0(\text_in_r[75] ),
    .I1(net231),
    .S(net21534),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input2 (.I(key[100]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31797_ (.I0(\text_in_r[76] ),
    .I1(net232),
    .S(net21534),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31798_ (.I0(\text_in_r[77] ),
    .I1(net233),
    .S(net21535),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31799_ (.I0(\text_in_r[78] ),
    .I1(net234),
    .S(net21535),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31800_ (.I0(\text_in_r[79] ),
    .I1(net235),
    .S(net21536),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31801_ (.I0(\text_in_r[7] ),
    .I1(net236),
    .S(net21539),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31802_ (.I0(\text_in_r[80] ),
    .I1(net237),
    .S(net21536),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31803_ (.I0(\text_in_r[81] ),
    .I1(net238),
    .S(net21536),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31804_ (.I0(\text_in_r[82] ),
    .I1(net239),
    .S(net21536),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31805_ (.I0(\text_in_r[83] ),
    .I1(net240),
    .S(net21536),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31806_ (.I0(\text_in_r[84] ),
    .I1(net241),
    .S(net21535),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(key[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31808_ (.I0(\text_in_r[85] ),
    .I1(net242),
    .S(net21535),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31809_ (.I0(\text_in_r[86] ),
    .I1(net243),
    .S(net21536),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31810_ (.I0(\text_in_r[87] ),
    .I1(net244),
    .S(net21536),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31811_ (.I0(\text_in_r[88] ),
    .I1(net245),
    .S(net21536),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31812_ (.I0(\text_in_r[89] ),
    .I1(net246),
    .S(net21536),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31813_ (.I0(\text_in_r[8] ),
    .I1(net247),
    .S(net21539),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31814_ (.I0(\text_in_r[90] ),
    .I1(net248),
    .S(net21536),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31815_ (.I0(\text_in_r[91] ),
    .I1(net249),
    .S(net21535),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31816_ (.I0(\text_in_r[92] ),
    .I1(net250),
    .S(net21536),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31817_ (.I0(\text_in_r[93] ),
    .I1(net251),
    .S(net21535),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31818_ (.I0(\text_in_r[94] ),
    .I1(net252),
    .S(net21537),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31819_ (.I0(\text_in_r[95] ),
    .I1(net253),
    .S(net21537),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31820_ (.I0(\text_in_r[96] ),
    .I1(net254),
    .S(net21537),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31821_ (.I0(\text_in_r[97] ),
    .I1(net255),
    .S(net21535),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31822_ (.I0(\text_in_r[98] ),
    .I1(net256),
    .S(net21535),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31823_ (.I0(\text_in_r[99] ),
    .I1(net257),
    .S(net21537),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _31824_ (.I0(\text_in_r[9] ),
    .I1(net258),
    .S(net21532),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31825_ (.A1(\dcnt[1] ),
    .A2(\dcnt[0] ),
    .ZN(_07499_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31826_ (.A1(_07461_),
    .A2(_07499_),
    .ZN(_07500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31827_ (.A1(_07500_),
    .A2(net130),
    .ZN(_07501_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31828_ (.A1(_07499_),
    .A2(_07460_),
    .Z(_07502_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31829_ (.A1(_07499_),
    .A2(_07460_),
    .ZN(_07503_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _31830_ (.A1(_07502_),
    .A2(_07503_),
    .ZN(_07505_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31831_ (.A1(_07501_),
    .A2(_07505_),
    .A3(net21535),
    .Z(_07506_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31832_ (.I(_07506_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31833_ (.A1(\u0.r0.rcnt[2] ),
    .A2(_16209_[0]),
    .Z(_07507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31834_ (.A1(\u0.r0.rcnt[2] ),
    .A2(_16209_[0]),
    .ZN(_07508_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _31835_ (.A1(_07507_),
    .A2(_07508_),
    .ZN(_07509_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31836_ (.A1(_07509_),
    .A2(_16207_[0]),
    .Z(_07510_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _31837_ (.A1(_07510_),
    .A2(net21535),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31838_ (.A1(\u0.r0.rcnt[2] ),
    .A2(\u0.r0.rcnt[1] ),
    .A3(\u0.r0.rcnt[0] ),
    .ZN(_07511_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _31839_ (.A1(\u0.r0.rcnt[3] ),
    .A2(_07511_),
    .Z(_07512_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31840_ (.I(_07512_),
    .ZN(_07514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31841_ (.I(_16202_[0]),
    .ZN(_07515_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _31842_ (.I(_07509_),
    .ZN(_07516_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31843_ (.A1(_07514_),
    .A2(_07515_),
    .A3(_07516_),
    .Z(_07517_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _31844_ (.A1(_07512_),
    .A2(\u0.r0.rcnt_next[1] ),
    .A3(_07516_),
    .Z(_07518_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31845_ (.A1(_07517_),
    .A2(_07518_),
    .B(net21535),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _31846_ (.A1(_07512_),
    .A2(_07515_),
    .A3(_07516_),
    .Z(_07519_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31847_ (.A1(_07512_),
    .A2(_16205_[0]),
    .A3(_07509_),
    .ZN(_07520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31848_ (.A1(_07519_),
    .A2(_07520_),
    .B(net21535),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _31849_ (.A1(_07512_),
    .A2(_16203_[0]),
    .A3(_07509_),
    .ZN(_07521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31850_ (.A1(_07514_),
    .A2(_07510_),
    .ZN(_07522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31851_ (.A1(_07521_),
    .A2(_07522_),
    .B(net21535),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _31852_ (.A1(_07512_),
    .A2(_07516_),
    .Z(_07523_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31853_ (.A1(_07523_),
    .A2(_16207_[0]),
    .ZN(_07524_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31854_ (.A1(_07518_),
    .A2(_07524_),
    .B(net21535),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31855_ (.A1(_07523_),
    .A2(_16202_[0]),
    .ZN(_07525_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31856_ (.A1(_07519_),
    .A2(_07525_),
    .B(net21535),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31857_ (.A1(_07523_),
    .A2(net21522),
    .A3(_16205_[0]),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _31858_ (.A1(_07523_),
    .A2(net21522),
    .A3(_16203_[0]),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31859_ (.A1(net21522),
    .A2(\u0.r0.rcnt_next[0] ),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31860_ (.A1(net21522),
    .A2(\u0.r0.rcnt_next[1] ),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31861_ (.A1(_07516_),
    .A2(net21522),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _31862_ (.A1(_07514_),
    .A2(net21522),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _31863_ (.A1(net21535),
    .A2(net130),
    .ZN(_07527_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _31864_ (.A1(_07501_),
    .A2(\dcnt[0] ),
    .B(_07527_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _31865_ (.A1(_07461_),
    .A2(\dcnt[1] ),
    .A3(\dcnt[0] ),
    .Z(_07528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31866_ (.A1(\dcnt[1] ),
    .A2(\dcnt[0] ),
    .B(net21535),
    .ZN(_07529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _31867_ (.I(net130),
    .ZN(_07530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _31868_ (.A1(_07528_),
    .A2(_07529_),
    .B(_07530_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _31869_ (.A1(_07502_),
    .A2(_07530_),
    .A3(_07459_),
    .B(_07527_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31870_ (.A(_15538_[0]),
    .B(_15537_[0]),
    .CO(_15539_[0]),
    .S(_15540_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31871_ (.A(net20834),
    .B(net20832),
    .CO(_15541_[0]),
    .S(_15542_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31872_ (.A(net20834),
    .B(_15543_[0]),
    .CO(_15544_[0]),
    .S(_15545_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31873_ (.A(net20834),
    .B(_15543_[0]),
    .CO(_15546_[0]),
    .S(_15547_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31874_ (.A(net20791),
    .B(net20832),
    .CO(_15549_[0]),
    .S(_15550_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31875_ (.A(_15538_[0]),
    .B(_15548_[0]),
    .CO(_15551_[0]),
    .S(_15552_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31876_ (.A(net20791),
    .B(_15543_[0]),
    .CO(_15553_[0]),
    .S(_15554_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31877_ (.A(net20791),
    .B(_15543_[0]),
    .CO(_15555_[0]),
    .S(_15556_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31878_ (.A(net20835),
    .B(_07976_),
    .CO(_15558_[0]),
    .S(_15559_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31879_ (.A(net20836),
    .B(net20554),
    .CO(_15560_[0]),
    .S(_15561_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31880_ (.A(net20835),
    .B(net20779),
    .CO(_15563_[0]),
    .S(_15564_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31881_ (.A(net20836),
    .B(net20777),
    .CO(_15565_[0]),
    .S(_15566_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31882_ (.A(net20792),
    .B(_07976_),
    .CO(_15567_[0]),
    .S(_15568_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31883_ (.A(net20792),
    .B(_07976_),
    .CO(_15569_[0]),
    .S(_15570_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31884_ (.A(_15572_[0]),
    .B(_15571_[0]),
    .CO(_15573_[0]),
    .S(_15574_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31885_ (.A(net20828),
    .B(net20820),
    .CO(_15575_[0]),
    .S(_15576_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31886_ (.A(net20828),
    .B(net20746),
    .CO(_15578_[0]),
    .S(_15579_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31887_ (.A(net20828),
    .B(_15577_[0]),
    .CO(_15580_[0]),
    .S(_15581_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31888_ (.A(net20741),
    .B(net20822),
    .CO(_15583_[0]),
    .S(_15584_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31889_ (.A(net20822),
    .B(_15582_[0]),
    .CO(_15585_[0]),
    .S(_15586_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31890_ (.A(net20741),
    .B(_15577_[0]),
    .CO(_15587_[0]),
    .S(_15588_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31891_ (.A(net20741),
    .B(_15577_[0]),
    .CO(_15589_[0]),
    .S(_15590_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31892_ (.A(net20830),
    .B(net20827),
    .CO(_15592_[0]),
    .S(_15593_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31893_ (.A(net20830),
    .B(net20823),
    .CO(_15594_[0]),
    .S(_15595_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31894_ (.A(net20831),
    .B(net20738),
    .CO(_15597_[0]),
    .S(_15598_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31895_ (.A(net20831),
    .B(net20738),
    .CO(_15599_[0]),
    .S(_15600_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31896_ (.A(net20744),
    .B(net20823),
    .CO(_15601_[0]),
    .S(_15602_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31897_ (.A(net20743),
    .B(net20823),
    .CO(_15603_[0]),
    .S(_15604_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31898_ (.A(_15606_[0]),
    .B(_15605_[0]),
    .CO(_15607_[0]),
    .S(_15608_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31899_ (.A(net20817),
    .B(net20812),
    .CO(_15609_[0]),
    .S(_15610_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31900_ (.A(net20817),
    .B(_15611_[0]),
    .CO(_15612_[0]),
    .S(_15613_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31901_ (.A(net20817),
    .B(_15611_[0]),
    .CO(_15614_[0]),
    .S(_15615_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31902_ (.A(_15616_[0]),
    .B(net20812),
    .CO(_15617_[0]),
    .S(_15618_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31903_ (.A(_15616_[0]),
    .B(net20812),
    .CO(_15619_[0]),
    .S(_15620_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31904_ (.A(net20774),
    .B(_15611_[0]),
    .CO(_15621_[0]),
    .S(_15622_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31905_ (.A(net20774),
    .B(_15611_[0]),
    .CO(_15623_[0]),
    .S(_15624_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31906_ (.A(net20818),
    .B(net20813),
    .CO(_15626_[0]),
    .S(_15627_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31907_ (.A(net20819),
    .B(net20814),
    .CO(_15628_[0]),
    .S(_15629_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31908_ (.A(net20818),
    .B(net20767),
    .CO(_15631_[0]),
    .S(_15632_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31909_ (.A(net20819),
    .B(net20768),
    .CO(_15633_[0]),
    .S(_15634_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31910_ (.A(net20773),
    .B(net20813),
    .CO(_15635_[0]),
    .S(_15636_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31911_ (.A(net20775),
    .B(net20814),
    .CO(_15637_[0]),
    .S(_15638_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31912_ (.A(_15639_[0]),
    .B(_15640_[0]),
    .CO(_15641_[0]),
    .S(_15642_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31913_ (.A(net20473),
    .B(net20471),
    .CO(_15643_[0]),
    .S(_15644_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31914_ (.A(net20473),
    .B(net20706),
    .CO(_15646_[0]),
    .S(_15647_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31915_ (.A(net20473),
    .B(_15645_[0]),
    .CO(_15648_[0]),
    .S(_15649_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31916_ (.A(net20703),
    .B(net20471),
    .CO(_15651_[0]),
    .S(_15652_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31917_ (.A(net20703),
    .B(net20471),
    .CO(_15653_[0]),
    .S(_15654_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31918_ (.A(net20703),
    .B(_15645_[0]),
    .CO(_15655_[0]),
    .S(_15656_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31919_ (.A(net20703),
    .B(net20707),
    .CO(_15657_[0]),
    .S(_15658_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31920_ (.A(net20810),
    .B(net20474),
    .CO(_15660_[0]),
    .S(_15661_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31921_ (.A(net20810),
    .B(net20474),
    .CO(_15662_[0]),
    .S(_15663_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31922_ (.A(net20697),
    .B(net20474),
    .CO(_15665_[0]),
    .S(_15666_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31923_ (.A(net20697),
    .B(net20474),
    .CO(_15667_[0]),
    .S(_15668_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31924_ (.A(net20697),
    .B(net20704),
    .CO(_15669_[0]),
    .S(_15670_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31925_ (.A(net20697),
    .B(net20704),
    .CO(_15671_[0]),
    .S(_15672_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31926_ (.A(_15674_[0]),
    .B(_15673_[0]),
    .CO(_15675_[0]),
    .S(_15676_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31927_ (.A(net19426),
    .B(net501),
    .CO(_15677_[0]),
    .S(_15678_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31928_ (.A(net19426),
    .B(_15679_[0]),
    .CO(_15680_[0]),
    .S(_15681_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31929_ (.A(net496),
    .B(net19398),
    .CO(_15683_[0]),
    .S(_15684_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31930_ (.A(_15682_[0]),
    .B(_15674_[0]),
    .CO(_15685_[0]),
    .S(_15686_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31931_ (.A(net19427),
    .B(net19431),
    .CO(_15687_[0]),
    .S(_15688_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31932_ (.A(net495),
    .B(_15679_[0]),
    .CO(_15689_[0]),
    .S(_15690_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31933_ (.A(net19868),
    .B(net19399),
    .CO(_15692_[0]),
    .S(_15693_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31934_ (.A(net19866),
    .B(net19431),
    .CO(_15694_[0]),
    .S(_15695_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31935_ (.A(net19866),
    .B(net19431),
    .CO(_15696_[0]),
    .S(_15697_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31936_ (.A(net19869),
    .B(net19399),
    .CO(_15699_[0]),
    .S(_15700_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31937_ (.A(net19869),
    .B(net19399),
    .CO(_15701_[0]),
    .S(_15702_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31938_ (.A(net19870),
    .B(net19429),
    .CO(_15703_[0]),
    .S(_15704_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31939_ (.A(_15705_[0]),
    .B(_15706_[0]),
    .CO(_15707_[0]),
    .S(_15708_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31940_ (.A(net19834),
    .B(net18915),
    .CO(_15709_[0]),
    .S(_15710_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31941_ (.A(net19834),
    .B(_11186_),
    .CO(_15712_[0]),
    .S(_15713_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31942_ (.A(_15714_[0]),
    .B(net18915),
    .CO(_15715_[0]),
    .S(_15716_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31943_ (.A(_15714_[0]),
    .B(net18915),
    .CO(_15717_[0]),
    .S(_15718_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31944_ (.A(net19837),
    .B(net18919),
    .CO(_15719_[0]),
    .S(_15720_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31945_ (.A(_15714_[0]),
    .B(_11186_),
    .CO(_15721_[0]),
    .S(_15722_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31946_ (.A(net19386),
    .B(net18918),
    .CO(_15724_[0]),
    .S(_15725_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31947_ (.A(net19386),
    .B(net18920),
    .CO(_15726_[0]),
    .S(_15727_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31948_ (.A(net19389),
    .B(net18920),
    .CO(_15728_[0]),
    .S(_15729_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31949_ (.A(net19396),
    .B(net18918),
    .CO(_15731_[0]),
    .S(_15732_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31950_ (.A(net19396),
    .B(net18918),
    .CO(_15733_[0]),
    .S(_15734_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31951_ (.A(net19396),
    .B(net18922),
    .CO(_15735_[0]),
    .S(_15736_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31952_ (.A(_15738_[0]),
    .B(_15737_[0]),
    .CO(_15739_[0]),
    .S(_15740_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31953_ (.A(net656),
    .B(net18314),
    .CO(_15741_[0]),
    .S(_15742_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31954_ (.A(_11997_),
    .B(_15737_[0]),
    .CO(_15744_[0]),
    .S(_15745_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31955_ (.A(net18315),
    .B(net19339),
    .CO(_15747_[0]),
    .S(_15748_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31956_ (.A(_15746_[0]),
    .B(net18314),
    .CO(_15749_[0]),
    .S(_15750_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31957_ (.A(net19340),
    .B(net435),
    .CO(_15751_[0]),
    .S(_15752_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31958_ (.A(_15746_[0]),
    .B(_11997_),
    .CO(_15753_[0]),
    .S(_15754_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31959_ (.A(net19330),
    .B(net18316),
    .CO(_15756_[0]),
    .S(_15757_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31960_ (.A(net19330),
    .B(net641),
    .CO(_15758_[0]),
    .S(_15759_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31961_ (.A(net19329),
    .B(net18320),
    .CO(_15760_[0]),
    .S(_15761_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31962_ (.A(net19336),
    .B(net18315),
    .CO(_15763_[0]),
    .S(_15764_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31963_ (.A(net19338),
    .B(net18316),
    .CO(_15765_[0]),
    .S(_15766_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31964_ (.A(net19338),
    .B(net641),
    .CO(_15767_[0]),
    .S(_15768_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31965_ (.A(_15770_[0]),
    .B(_15769_[0]),
    .CO(_15771_[0]),
    .S(_15772_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31966_ (.A(net19285),
    .B(net19273),
    .CO(_15773_[0]),
    .S(_15774_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31967_ (.A(net19284),
    .B(_15775_[0]),
    .CO(_15776_[0]),
    .S(_15777_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31968_ (.A(net19294),
    .B(net19273),
    .CO(_15779_[0]),
    .S(_15780_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31969_ (.A(_15778_[0]),
    .B(net19273),
    .CO(_15781_[0]),
    .S(_15782_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31970_ (.A(net19296),
    .B(net19299),
    .CO(_15783_[0]),
    .S(_15784_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31971_ (.A(_15778_[0]),
    .B(_15775_[0]),
    .CO(_15785_[0]),
    .S(_15786_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31972_ (.A(net19281),
    .B(net19276),
    .CO(_15788_[0]),
    .S(_15789_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31973_ (.A(_12861_),
    .B(net19298),
    .CO(_15790_[0]),
    .S(_15791_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31974_ (.A(net19283),
    .B(net19299),
    .CO(_15792_[0]),
    .S(_15793_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31975_ (.A(net19292),
    .B(net19275),
    .CO(_15795_[0]),
    .S(_15796_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31976_ (.A(net19290),
    .B(net19274),
    .CO(_15797_[0]),
    .S(_15798_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31977_ (.A(net19293),
    .B(net19298),
    .CO(_15799_[0]),
    .S(_15800_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31978_ (.A(_15801_[0]),
    .B(_15802_[0]),
    .CO(_15803_[0]),
    .S(_15804_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31979_ (.A(net604),
    .B(net19242),
    .CO(_15805_[0]),
    .S(_15806_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31980_ (.A(_15807_[0]),
    .B(net604),
    .CO(_15808_[0]),
    .S(_15809_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31981_ (.A(_15810_[0]),
    .B(net19242),
    .CO(_15811_[0]),
    .S(_15812_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _31982_ (.A(_15810_[0]),
    .B(net619),
    .CO(_15813_[0]),
    .S(_15814_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31983_ (.A(net19807),
    .B(net19259),
    .CO(_15815_[0]),
    .S(_15816_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31984_ (.A(_15810_[0]),
    .B(_15807_[0]),
    .CO(_15817_[0]),
    .S(_15818_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31985_ (.A(net19799),
    .B(net430),
    .CO(_15820_[0]),
    .S(_15821_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31986_ (.A(net19800),
    .B(net19261),
    .CO(_15822_[0]),
    .S(_15823_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31987_ (.A(net19800),
    .B(net19261),
    .CO(_15824_[0]),
    .S(_15825_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31988_ (.A(net395),
    .B(net19243),
    .CO(_15827_[0]),
    .S(_15828_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31989_ (.A(net395),
    .B(net19243),
    .CO(_15829_[0]),
    .S(_15830_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31990_ (.A(net19803),
    .B(net19261),
    .CO(_15831_[0]),
    .S(_15832_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31991_ (.A(_15834_[0]),
    .B(_15833_[0]),
    .CO(_15835_[0]),
    .S(_15836_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31992_ (.A(net19786),
    .B(net19224),
    .CO(_15837_[0]),
    .S(_15838_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31993_ (.A(_15839_[0]),
    .B(net19786),
    .CO(_15840_[0]),
    .S(_15841_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31994_ (.A(_15842_[0]),
    .B(net19227),
    .CO(_15843_[0]),
    .S(_15844_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31995_ (.A(_15842_[0]),
    .B(net19224),
    .CO(_15845_[0]),
    .S(_15846_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31996_ (.A(net19797),
    .B(net19230),
    .CO(_15847_[0]),
    .S(_15848_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31997_ (.A(_15842_[0]),
    .B(_15839_[0]),
    .CO(_15849_[0]),
    .S(_15850_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31998_ (.A(net19780),
    .B(net19225),
    .CO(_15852_[0]),
    .S(_15853_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _31999_ (.A(net19784),
    .B(net19230),
    .CO(_15854_[0]),
    .S(_15855_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32000_ (.A(net19785),
    .B(net19230),
    .CO(_15856_[0]),
    .S(_15857_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32001_ (.A(_14379_),
    .B(net19225),
    .CO(_15859_[0]),
    .S(_15860_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32002_ (.A(net19793),
    .B(net19225),
    .CO(_15861_[0]),
    .S(_15862_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32003_ (.A(net19789),
    .B(net19229),
    .CO(_15863_[0]),
    .S(_15864_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32004_ (.A(_15865_[0]),
    .B(_15866_[0]),
    .CO(_15867_[0]),
    .S(_15868_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32005_ (.A(net19207),
    .B(net18200),
    .CO(_15869_[0]),
    .S(_15870_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32006_ (.A(_15871_[0]),
    .B(_15865_[0]),
    .CO(_15872_[0]),
    .S(_15873_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32007_ (.A(net19210),
    .B(net401),
    .CO(_15875_[0]),
    .S(_15876_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32008_ (.A(_15874_[0]),
    .B(net399),
    .CO(_15877_[0]),
    .S(_15878_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32009_ (.A(net19209),
    .B(net18204),
    .CO(_15879_[0]),
    .S(_15880_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32010_ (.A(_15874_[0]),
    .B(net406),
    .CO(_15881_[0]),
    .S(_15882_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32011_ (.A(net19768),
    .B(net18201),
    .CO(_15884_[0]),
    .S(_15885_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32012_ (.A(net19768),
    .B(net18207),
    .CO(_15886_[0]),
    .S(_15887_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32013_ (.A(net19768),
    .B(net18207),
    .CO(_15888_[0]),
    .S(_15889_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32014_ (.A(net19772),
    .B(net18203),
    .CO(_15891_[0]),
    .S(_15892_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32015_ (.A(net19769),
    .B(net18202),
    .CO(_15893_[0]),
    .S(_15894_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32016_ (.A(net19772),
    .B(net18207),
    .CO(_15895_[0]),
    .S(_15896_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32017_ (.A(_15898_[0]),
    .B(_15897_[0]),
    .CO(_15899_[0]),
    .S(_15900_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32018_ (.A(net19735),
    .B(net19196),
    .CO(_15901_[0]),
    .S(_15902_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32019_ (.A(_15903_[0]),
    .B(net19735),
    .CO(_15904_[0]),
    .S(_15905_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32020_ (.A(_15906_[0]),
    .B(net19197),
    .CO(_15907_[0]),
    .S(_15908_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32021_ (.A(_15906_[0]),
    .B(net19196),
    .CO(_15909_[0]),
    .S(_15910_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32022_ (.A(net19741),
    .B(net427),
    .CO(_15911_[0]),
    .S(_15912_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32023_ (.A(_15903_[0]),
    .B(_15906_[0]),
    .CO(_15913_[0]),
    .S(_15914_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32024_ (.A(net19731),
    .B(net19198),
    .CO(_15916_[0]),
    .S(_15917_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32025_ (.A(net19731),
    .B(net427),
    .CO(_15918_[0]),
    .S(_15919_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32026_ (.A(net19733),
    .B(net427),
    .CO(_15920_[0]),
    .S(_15921_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32027_ (.A(net19739),
    .B(net19197),
    .CO(_15923_[0]),
    .S(_15924_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32028_ (.A(net19739),
    .B(net19198),
    .CO(_15925_[0]),
    .S(_15926_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32029_ (.A(net19739),
    .B(net427),
    .CO(_15927_[0]),
    .S(_15928_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32030_ (.A(_15930_[0]),
    .B(_15929_[0]),
    .CO(_15931_[0]),
    .S(_15932_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32031_ (.A(_15929_[0]),
    .B(_15930_[0]),
    .CO(_15933_[0]),
    .S(_15934_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32032_ (.A(_15935_[0]),
    .B(net19719),
    .CO(_15936_[0]),
    .S(_15937_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32033_ (.A(net19719),
    .B(_15935_[0]),
    .CO(_15938_[0]),
    .S(_15939_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32034_ (.A(net19721),
    .B(net18648),
    .CO(_15941_[0]),
    .S(_15942_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32035_ (.A(_15940_[0]),
    .B(net18649),
    .CO(_15943_[0]),
    .S(_15944_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32036_ (.A(_15935_[0]),
    .B(_15940_[0]),
    .CO(_15945_[0]),
    .S(_15946_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32037_ (.A(_15935_[0]),
    .B(_15940_[0]),
    .CO(_15947_[0]),
    .S(_15948_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32038_ (.A(net19189),
    .B(net18648),
    .CO(_15950_[0]),
    .S(_15951_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32039_ (.A(net19189),
    .B(net389),
    .CO(_15952_[0]),
    .S(_15953_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32040_ (.A(net19189),
    .B(net389),
    .CO(_15954_[0]),
    .S(_15955_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32041_ (.A(net19195),
    .B(net18648),
    .CO(_15957_[0]),
    .S(_15958_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32042_ (.A(net19192),
    .B(net18648),
    .CO(_15959_[0]),
    .S(_15960_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32043_ (.A(net19192),
    .B(net389),
    .CO(_15961_[0]),
    .S(_15962_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32044_ (.A(net19192),
    .B(net389),
    .CO(_15963_[0]),
    .S(_15964_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32045_ (.A(_15965_[0]),
    .B(_15966_[0]),
    .CO(_15967_[0]),
    .S(_15968_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32046_ (.A(net19171),
    .B(net19174),
    .CO(_15969_[0]),
    .S(_15970_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32047_ (.A(net19171),
    .B(net441),
    .CO(_15972_[0]),
    .S(_15973_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32048_ (.A(_15971_[0]),
    .B(net19171),
    .CO(_15974_[0]),
    .S(_15975_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32049_ (.A(net19177),
    .B(net19175),
    .CO(_15977_[0]),
    .S(_15978_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32050_ (.A(_15976_[0]),
    .B(net19174),
    .CO(_15979_[0]),
    .S(_15980_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32051_ (.A(net687),
    .B(net19180),
    .CO(_15981_[0]),
    .S(_15982_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32052_ (.A(_15976_[0]),
    .B(_15971_[0]),
    .CO(_15983_[0]),
    .S(_15984_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32053_ (.A(net19696),
    .B(net19175),
    .CO(_15986_[0]),
    .S(_15987_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32054_ (.A(net19696),
    .B(net19181),
    .CO(_15988_[0]),
    .S(_15989_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32055_ (.A(net19696),
    .B(net19181),
    .CO(_15990_[0]),
    .S(_15991_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32056_ (.A(net19699),
    .B(net19176),
    .CO(_15993_[0]),
    .S(_15994_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32057_ (.A(net19699),
    .B(net19175),
    .CO(_15995_[0]),
    .S(_15996_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32058_ (.A(net19699),
    .B(net19181),
    .CO(_15997_[0]),
    .S(_15998_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32059_ (.A(net19701),
    .B(net19181),
    .CO(_15999_[0]),
    .S(_16000_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32060_ (.A(_16001_[0]),
    .B(_16002_[0]),
    .CO(_16003_[0]),
    .S(_16004_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32061_ (.A(net19147),
    .B(net18565),
    .CO(_16005_[0]),
    .S(_16006_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32062_ (.A(net19147),
    .B(net527),
    .CO(_16008_[0]),
    .S(_16009_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32063_ (.A(net19145),
    .B(_16007_[0]),
    .CO(_16010_[0]),
    .S(_16011_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32064_ (.A(net19670),
    .B(net18565),
    .CO(_16013_[0]),
    .S(_16014_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32065_ (.A(net19669),
    .B(net18565),
    .CO(_16015_[0]),
    .S(_16016_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32066_ (.A(net19671),
    .B(net528),
    .CO(_16017_[0]),
    .S(_16018_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32067_ (.A(net19669),
    .B(net527),
    .CO(_16019_[0]),
    .S(_16020_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32068_ (.A(_03083_),
    .B(net18565),
    .CO(_16022_[0]),
    .S(_16023_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32069_ (.A(net19658),
    .B(net18567),
    .CO(_16024_[0]),
    .S(_16025_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32070_ (.A(net19660),
    .B(net18567),
    .CO(_16026_[0]),
    .S(_16027_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32071_ (.A(net19668),
    .B(net18564),
    .CO(_16029_[0]),
    .S(_16030_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32072_ (.A(net19663),
    .B(net18565),
    .CO(_16031_[0]),
    .S(_16032_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32073_ (.A(net19667),
    .B(net18567),
    .CO(_16033_[0]),
    .S(_16034_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32074_ (.A(net19667),
    .B(net18567),
    .CO(_16035_[0]),
    .S(_16036_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32075_ (.A(_16038_[0]),
    .B(_16037_[0]),
    .CO(_16039_[0]),
    .S(_16040_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32076_ (.A(_16037_[0]),
    .B(_16038_[0]),
    .CO(_16041_[0]),
    .S(_16042_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32077_ (.A(net19122),
    .B(net19138),
    .CO(_16044_[0]),
    .S(_16045_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32078_ (.A(_16043_[0]),
    .B(_16037_[0]),
    .CO(_16046_[0]),
    .S(_16047_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32079_ (.A(net19133),
    .B(net404),
    .CO(_16049_[0]),
    .S(_16050_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32080_ (.A(net405),
    .B(_16048_[0]),
    .CO(_16051_[0]),
    .S(_16052_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32081_ (.A(net19133),
    .B(net19138),
    .CO(_16053_[0]),
    .S(_16054_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32082_ (.A(_16048_[0]),
    .B(net478),
    .CO(_16055_[0]),
    .S(_16056_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32083_ (.A(net19650),
    .B(net19125),
    .CO(_16058_[0]),
    .S(_16059_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32084_ (.A(net19650),
    .B(net19139),
    .CO(_16060_[0]),
    .S(_16061_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32085_ (.A(net19653),
    .B(net19139),
    .CO(_16062_[0]),
    .S(_16063_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32086_ (.A(net19127),
    .B(net19126),
    .CO(_16065_[0]),
    .S(_16066_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32087_ (.A(_03833_),
    .B(net19125),
    .CO(_16067_[0]),
    .S(_16068_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32088_ (.A(net19131),
    .B(net19139),
    .CO(_16069_[0]),
    .S(_16070_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32089_ (.A(net19128),
    .B(net19136),
    .CO(_16071_[0]),
    .S(_16072_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32090_ (.A(_04571_),
    .B(_16074_[0]),
    .CO(_16075_[0]),
    .S(_16076_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32091_ (.A(net19609),
    .B(net509),
    .CO(_16077_[0]),
    .S(_16078_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32092_ (.A(_04571_),
    .B(_16079_[0]),
    .CO(_16080_[0]),
    .S(_16081_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32093_ (.A(net512),
    .B(net19601),
    .CO(_16083_[0]),
    .S(_16084_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32094_ (.A(net512),
    .B(net19601),
    .CO(_16085_[0]),
    .S(_16086_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32095_ (.A(net19617),
    .B(net19619),
    .CO(_16087_[0]),
    .S(_16088_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32096_ (.A(_16082_[0]),
    .B(_16079_[0]),
    .CO(_16089_[0]),
    .S(_16090_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32097_ (.A(net19606),
    .B(net19602),
    .CO(_16092_[0]),
    .S(_16093_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32098_ (.A(net19606),
    .B(net19619),
    .CO(_16094_[0]),
    .S(_16095_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32099_ (.A(net19606),
    .B(net19619),
    .CO(_16096_[0]),
    .S(_16097_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32100_ (.A(net19615),
    .B(net19602),
    .CO(_16099_[0]),
    .S(_16100_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32101_ (.A(net19614),
    .B(net19602),
    .CO(_16101_[0]),
    .S(_16102_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32102_ (.A(net19611),
    .B(net19618),
    .CO(_16103_[0]),
    .S(_16104_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32103_ (.A(_16106_[0]),
    .B(_16105_[0]),
    .CO(_16107_[0]),
    .S(_16108_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32104_ (.A(net19564),
    .B(net19017),
    .CO(_16109_[0]),
    .S(_16110_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32105_ (.A(_16111_[0]),
    .B(_16105_[0]),
    .CO(_16112_[0]),
    .S(_16113_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32106_ (.A(_16114_[0]),
    .B(net19018),
    .CO(_16115_[0]),
    .S(_16116_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32107_ (.A(_16114_[0]),
    .B(net19017),
    .CO(_16117_[0]),
    .S(_16118_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32108_ (.A(net19570),
    .B(net19060),
    .CO(_16119_[0]),
    .S(_16120_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32109_ (.A(_16114_[0]),
    .B(net19059),
    .CO(_16121_[0]),
    .S(_16122_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32110_ (.A(net19568),
    .B(net19019),
    .CO(_16124_[0]),
    .S(_16125_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32111_ (.A(net19569),
    .B(net19060),
    .CO(_16126_[0]),
    .S(_16127_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32112_ (.A(net19569),
    .B(net19060),
    .CO(_16128_[0]),
    .S(_16129_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32113_ (.A(net19058),
    .B(net19019),
    .CO(_16131_[0]),
    .S(_16132_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32114_ (.A(_05303_),
    .B(net19019),
    .CO(_16133_[0]),
    .S(_16134_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32115_ (.A(net19057),
    .B(net19060),
    .CO(_16135_[0]),
    .S(_16136_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32116_ (.A(_16137_[0]),
    .B(_16138_[0]),
    .CO(_16139_[0]),
    .S(_16140_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32117_ (.A(_16137_[0]),
    .B(net19008),
    .CO(_16141_[0]),
    .S(_16142_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32118_ (.A(_16137_[0]),
    .B(_05987_),
    .CO(_16144_[0]),
    .S(_16145_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32119_ (.A(_16146_[0]),
    .B(net19009),
    .CO(_16147_[0]),
    .S(_16148_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32120_ (.A(_16146_[0]),
    .B(net19009),
    .CO(_16149_[0]),
    .S(_16150_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32121_ (.A(net19542),
    .B(net19012),
    .CO(_16151_[0]),
    .S(_16152_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32122_ (.A(_16146_[0]),
    .B(_05987_),
    .CO(_16153_[0]),
    .S(_16154_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32123_ (.A(net19530),
    .B(net19010),
    .CO(_16156_[0]),
    .S(_16157_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32124_ (.A(net19530),
    .B(net19014),
    .CO(_16158_[0]),
    .S(_16159_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32125_ (.A(net19530),
    .B(net19014),
    .CO(_16160_[0]),
    .S(_16161_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32126_ (.A(net19541),
    .B(net19010),
    .CO(_16163_[0]),
    .S(_16164_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32127_ (.A(net19541),
    .B(net19010),
    .CO(_16165_[0]),
    .S(_16166_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32128_ (.A(net19541),
    .B(net19014),
    .CO(_16167_[0]),
    .S(_16168_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32129_ (.A(_16170_[0]),
    .B(_16169_[0]),
    .CO(_16171_[0]),
    .S(_16172_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32130_ (.A(net19456),
    .B(net517),
    .CO(_16173_[0]),
    .S(_16174_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32131_ (.A(net19455),
    .B(_06726_),
    .CO(_16176_[0]),
    .S(_16177_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32132_ (.A(net397),
    .B(net518),
    .CO(_16179_[0]),
    .S(_16180_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32133_ (.A(_16178_[0]),
    .B(net18958),
    .CO(_16181_[0]),
    .S(_16182_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32134_ (.A(net19465),
    .B(net18999),
    .CO(_16183_[0]),
    .S(_16184_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _32135_ (.A(_16178_[0]),
    .B(_06726_),
    .CO(_16185_[0]),
    .S(_16186_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32136_ (.A(net19458),
    .B(net519),
    .CO(_16188_[0]),
    .S(_16189_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32137_ (.A(net19462),
    .B(net19000),
    .CO(_16190_[0]),
    .S(_16191_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32138_ (.A(net19462),
    .B(net19000),
    .CO(_16192_[0]),
    .S(_16193_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32139_ (.A(_06763_),
    .B(net519),
    .CO(_16195_[0]),
    .S(_16196_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32140_ (.A(_06763_),
    .B(net519),
    .CO(_16197_[0]),
    .S(_16198_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32141_ (.A(net18997),
    .B(net19000),
    .CO(_16199_[0]),
    .S(_16200_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32142_ (.A(\u0.r0.rcnt_next[0] ),
    .B(_16201_[0]),
    .CO(_16202_[0]),
    .S(\u0.r0.rcnt_next[1] ));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32143_ (.A(\u0.r0.rcnt_next[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_16203_[0]),
    .S(_16204_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32144_ (.A(\u0.r0.rcnt[0] ),
    .B(_16201_[0]),
    .CO(_16205_[0]),
    .S(_16206_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32145_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_16207_[0]),
    .S(_16208_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _32146_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_16209_[0]),
    .S(_16210_[0]));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dcnt[0]$_SDFFE_PN0P_  (.D(_00405_),
    .CLK(clknet_leaf_67_clk),
    .Q(\dcnt[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dcnt[1]$_SDFFE_PN0P_  (.D(_00406_),
    .CLK(clknet_leaf_67_clk),
    .Q(\dcnt[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dcnt[2]$_SDFFE_PP0P_  (.D(_00407_),
    .CLK(clknet_leaf_64_clk),
    .Q(\dcnt[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dcnt[3]$_SDFFE_PN0P_  (.D(_00408_),
    .CLK(clknet_leaf_64_clk),
    .Q(\dcnt[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \done$_DFF_P_  (.D(_00160_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(net259));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \ld_r$_DFF_P_  (.D(net21539),
    .CLK(clknet_leaf_349_clk),
    .Q(ld_r));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa00_sr[0]$_DFF_P_  (.D(_00032_),
    .CLK(clknet_leaf_257_clk),
    .Q(\sa00_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[1]$_DFF_P_  (.D(_00033_),
    .CLK(clknet_5_25__leaf_clk),
    .Q(\sa00_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[2]$_DFF_P_  (.D(_00034_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\sa00_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[3]$_DFF_P_  (.D(_00035_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\sa00_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[4]$_DFF_P_  (.D(_00036_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(\sa00_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[5]$_DFF_P_  (.D(_00037_),
    .CLK(clknet_5_25__leaf_clk),
    .Q(\sa00_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[6]$_DFF_P_  (.D(_00038_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\sa00_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa00_sr[7]$_DFF_P_  (.D(_00039_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\sa00_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa01_sr[0]$_DFF_P_  (.D(_00040_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(\sa01_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa01_sr[1]$_DFF_P_  (.D(_00041_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(\sa01_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa01_sr[2]$_DFF_P_  (.D(_00042_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\sa01_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa01_sr[3]$_DFF_P_  (.D(_00043_),
    .CLK(clknet_leaf_106_clk),
    .Q(\sa01_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa01_sr[4]$_DFF_P_  (.D(_00044_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(\sa01_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa01_sr[5]$_DFF_P_  (.D(_00045_),
    .CLK(clknet_leaf_106_clk),
    .Q(\sa01_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa01_sr[6]$_DFF_P_  (.D(_00046_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\sa01_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa01_sr[7]$_DFF_P_  (.D(_00047_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\sa01_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa02_sr[0]$_DFF_P_  (.D(_00048_),
    .CLK(clknet_leaf_221_clk),
    .Q(\sa02_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[1]$_DFF_P_  (.D(_00049_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\sa02_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[2]$_DFF_P_  (.D(_00050_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\sa02_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[3]$_DFF_P_  (.D(_00051_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\sa02_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[4]$_DFF_P_  (.D(_00052_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\sa02_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[5]$_DFF_P_  (.D(_00053_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\sa02_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[6]$_DFF_P_  (.D(_00054_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\sa02_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa02_sr[7]$_DFF_P_  (.D(_00055_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\sa02_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa03_sr[0]$_DFF_P_  (.D(_00056_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(\sa03_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa03_sr[1]$_DFF_P_  (.D(_00057_),
    .CLK(clknet_leaf_315_clk),
    .Q(\sa03_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[2]$_DFF_P_  (.D(_00058_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(\sa03_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[3]$_DFF_P_  (.D(_00059_),
    .CLK(clknet_leaf_290_clk),
    .Q(\sa03_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[4]$_DFF_P_  (.D(_00060_),
    .CLK(clknet_leaf_290_clk),
    .Q(\sa03_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[5]$_DFF_P_  (.D(_00061_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(\sa03_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa03_sr[6]$_DFF_P_  (.D(_00062_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(\sa03_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa03_sr[7]$_DFF_P_  (.D(_00063_),
    .CLK(clknet_leaf_290_clk),
    .Q(\sa03_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[0]$_DFF_P_  (.D(_00072_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\sa10_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[1]$_DFF_P_  (.D(_00073_),
    .CLK(clknet_leaf_58_clk),
    .Q(\sa10_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa10_sr[2]$_DFF_P_  (.D(_00074_),
    .CLK(clknet_leaf_86_clk),
    .Q(\sa10_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa10_sr[3]$_DFF_P_  (.D(_00075_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(\sa10_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa10_sr[4]$_DFF_P_  (.D(_00076_),
    .CLK(clknet_leaf_91_clk),
    .Q(\sa10_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa10_sr[5]$_DFF_P_  (.D(_00077_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\sa10_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa10_sr[6]$_DFF_P_  (.D(_00078_),
    .CLK(clknet_leaf_75_clk),
    .Q(\sa10_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa10_sr[7]$_DFF_P_  (.D(_00079_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(\sa10_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[0]$_DFF_P_  (.D(_00080_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\sa11_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa11_sr[1]$_DFF_P_  (.D(_00081_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\sa11_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa11_sr[2]$_DFF_P_  (.D(_00082_),
    .CLK(clknet_leaf_123_clk),
    .Q(\sa11_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa11_sr[3]$_DFF_P_  (.D(_00083_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\sa11_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa11_sr[4]$_DFF_P_  (.D(_00084_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\sa11_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa11_sr[5]$_DFF_P_  (.D(_00085_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\sa11_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa11_sr[6]$_DFF_P_  (.D(_00086_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\sa11_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa11_sr[7]$_DFF_P_  (.D(_00087_),
    .CLK(clknet_leaf_123_clk),
    .Q(\sa11_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa12_sr[0]$_DFF_P_  (.D(_00088_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\sa12_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[1]$_DFF_P_  (.D(_00089_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(\sa12_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[2]$_DFF_P_  (.D(_00090_),
    .CLK(clknet_leaf_277_clk),
    .Q(\sa12_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa12_sr[3]$_DFF_P_  (.D(_00091_),
    .CLK(clknet_leaf_289_clk),
    .Q(\sa12_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[4]$_DFF_P_  (.D(_00092_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\sa12_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[5]$_DFF_P_  (.D(_00093_),
    .CLK(clknet_leaf_289_clk),
    .Q(\sa12_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa12_sr[6]$_DFF_P_  (.D(_00094_),
    .CLK(clknet_leaf_277_clk),
    .Q(\sa12_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa12_sr[7]$_DFF_P_  (.D(_00095_),
    .CLK(clknet_leaf_231_clk),
    .Q(\sa12_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa13_sr[0]$_DFF_P_  (.D(_00064_),
    .CLK(clknet_leaf_301_clk),
    .Q(\sa10_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa13_sr[1]$_DFF_P_  (.D(_00065_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\sa10_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa13_sr[2]$_DFF_P_  (.D(_00066_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(\sa10_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa13_sr[3]$_DFF_P_  (.D(_00067_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\sa10_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa13_sr[4]$_DFF_P_  (.D(_00068_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(\sa10_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa13_sr[5]$_DFF_P_  (.D(_00069_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\sa10_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa13_sr[6]$_DFF_P_  (.D(_00070_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\sa10_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa13_sr[7]$_DFF_P_  (.D(_00071_),
    .CLK(clknet_leaf_301_clk),
    .Q(\sa10_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa20_sr[0]$_DFF_P_  (.D(_00112_),
    .CLK(clknet_5_30__leaf_clk),
    .Q(\sa20_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa20_sr[1]$_DFF_P_  (.D(_00113_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa20_sr[2]$_DFF_P_  (.D(_00114_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa20_sr[3]$_DFF_P_  (.D(_00115_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa20_sr[4]$_DFF_P_  (.D(_00116_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa20_sr[5]$_DFF_P_  (.D(_00117_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\sa20_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa20_sr[6]$_DFF_P_  (.D(_00118_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa20_sr[7]$_DFF_P_  (.D(_00119_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\sa20_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[0]$_DFF_P_  (.D(_00120_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\sa21_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[1]$_DFF_P_  (.D(_00121_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\sa21_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[2]$_DFF_P_  (.D(_00122_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\sa21_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa21_sr[3]$_DFF_P_  (.D(_00123_),
    .CLK(clknet_leaf_96_clk),
    .Q(\sa21_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa21_sr[4]$_DFF_P_  (.D(_00124_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\sa21_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa21_sr[5]$_DFF_P_  (.D(_00125_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\sa21_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa21_sr[6]$_DFF_P_  (.D(_00126_),
    .CLK(clknet_leaf_96_clk),
    .Q(\sa21_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa21_sr[7]$_DFF_P_  (.D(_00127_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\sa21_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa22_sr[0]$_DFF_P_  (.D(_00096_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa22_sr[1]$_DFF_P_  (.D(_00097_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa22_sr[2]$_DFF_P_  (.D(_00098_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa22_sr[3]$_DFF_P_  (.D(_00099_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa22_sr[4]$_DFF_P_  (.D(_00100_),
    .CLK(clknet_leaf_191_clk),
    .Q(\sa20_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa22_sr[5]$_DFF_P_  (.D(_00101_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(\sa20_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa22_sr[6]$_DFF_P_  (.D(_00102_),
    .CLK(clknet_leaf_191_clk),
    .Q(\sa20_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa22_sr[7]$_DFF_P_  (.D(_00103_),
    .CLK(clknet_leaf_246_clk),
    .Q(\sa20_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[0]$_DFF_P_  (.D(_00104_),
    .CLK(clknet_leaf_399_clk),
    .Q(\sa21_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa23_sr[1]$_DFF_P_  (.D(_00105_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(\sa21_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa23_sr[2]$_DFF_P_  (.D(_00106_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\sa21_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa23_sr[3]$_DFF_P_  (.D(_00107_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\sa21_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa23_sr[4]$_DFF_P_  (.D(_00108_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\sa21_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa23_sr[5]$_DFF_P_  (.D(_00109_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\sa21_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa23_sr[6]$_DFF_P_  (.D(_00110_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\sa21_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa23_sr[7]$_DFF_P_  (.D(_00111_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\sa21_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa30_sr[0]$_DFF_P_  (.D(_00152_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\sa30_sr[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa30_sr[1]$_DFF_P_  (.D(_00153_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\sa30_sr[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa30_sr[2]$_DFF_P_  (.D(_00154_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(\sa30_sr[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa30_sr[3]$_DFF_P_  (.D(_00155_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(\sa30_sr[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa30_sr[4]$_DFF_P_  (.D(_00156_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(\sa30_sr[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa30_sr[5]$_DFF_P_  (.D(_00157_),
    .CLK(clknet_leaf_273_clk),
    .Q(\sa30_sr[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa30_sr[6]$_DFF_P_  (.D(_00158_),
    .CLK(clknet_leaf_270_clk),
    .Q(\sa30_sr[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa30_sr[7]$_DFF_P_  (.D(_00159_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\sa30_sr[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa31_sr[0]$_DFF_P_  (.D(_00128_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(\sa30_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa31_sr[1]$_DFF_P_  (.D(_00129_),
    .CLK(clknet_leaf_130_clk),
    .Q(\sa30_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa31_sr[2]$_DFF_P_  (.D(_00130_),
    .CLK(clknet_leaf_126_clk),
    .Q(\sa30_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa31_sr[3]$_DFF_P_  (.D(_00131_),
    .CLK(clknet_leaf_127_clk),
    .Q(\sa30_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa31_sr[4]$_DFF_P_  (.D(_00132_),
    .CLK(clknet_leaf_130_clk),
    .Q(\sa30_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa31_sr[5]$_DFF_P_  (.D(_00133_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(\sa30_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa31_sr[6]$_DFF_P_  (.D(_00134_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(\sa30_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa31_sr[7]$_DFF_P_  (.D(_00135_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(\sa30_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[0]$_DFF_P_  (.D(_00136_),
    .CLK(clknet_leaf_207_clk),
    .Q(\sa31_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[1]$_DFF_P_  (.D(_00137_),
    .CLK(clknet_leaf_207_clk),
    .Q(\sa31_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa32_sr[2]$_DFF_P_  (.D(_00138_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\sa31_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa32_sr[3]$_DFF_P_  (.D(_00139_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\sa31_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa32_sr[4]$_DFF_P_  (.D(_00140_),
    .CLK(clknet_leaf_246_clk),
    .Q(\sa31_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa32_sr[5]$_DFF_P_  (.D(_00141_),
    .CLK(clknet_leaf_249_clk),
    .Q(\sa31_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa32_sr[6]$_DFF_P_  (.D(_00142_),
    .CLK(clknet_5_25__leaf_clk),
    .Q(\sa31_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa32_sr[7]$_DFF_P_  (.D(_00143_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\sa31_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[0]$_DFF_P_  (.D(_00144_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(\sa32_sub[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[1]$_DFF_P_  (.D(_00145_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(\sa32_sub[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa33_sr[2]$_DFF_P_  (.D(_00146_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\sa32_sub[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[3]$_DFF_P_  (.D(_00147_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\sa32_sub[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[4]$_DFF_P_  (.D(_00148_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\sa32_sub[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[5]$_DFF_P_  (.D(_00149_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\sa32_sub[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \sa33_sr[6]$_DFF_P_  (.D(_00150_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\sa32_sub[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \sa33_sr[7]$_DFF_P_  (.D(_00151_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(\sa32_sub[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[0]$_DFFE_PP_  (.D(_00409_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\text_in_r[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[100]$_DFFE_PP_  (.D(_00410_),
    .CLK(clknet_leaf_144_clk),
    .Q(\text_in_r[100] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[101]$_DFFE_PP_  (.D(_00411_),
    .CLK(clknet_leaf_362_clk),
    .Q(\text_in_r[101] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[102]$_DFFE_PP_  (.D(_00412_),
    .CLK(clknet_leaf_362_clk),
    .Q(\text_in_r[102] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[103]$_DFFE_PP_  (.D(_00413_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\text_in_r[103] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[104]$_DFFE_PP_  (.D(_00414_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\text_in_r[104] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[105]$_DFFE_PP_  (.D(_00415_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\text_in_r[105] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[106]$_DFFE_PP_  (.D(_00416_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\text_in_r[106] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[107]$_DFFE_PP_  (.D(_00417_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\text_in_r[107] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[108]$_DFFE_PP_  (.D(_00418_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\text_in_r[108] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[109]$_DFFE_PP_  (.D(_00419_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\text_in_r[109] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[10]$_DFFE_PP_  (.D(_00420_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[110]$_DFFE_PP_  (.D(_00421_),
    .CLK(clknet_leaf_358_clk),
    .Q(\text_in_r[110] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[111]$_DFFE_PP_  (.D(_00422_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\text_in_r[111] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[112]$_DFFE_PP_  (.D(_00423_),
    .CLK(clknet_leaf_39_clk),
    .Q(\text_in_r[112] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[113]$_DFFE_PP_  (.D(_00424_),
    .CLK(clknet_leaf_377_clk),
    .Q(\text_in_r[113] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[114]$_DFFE_PP_  (.D(_00425_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\text_in_r[114] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[115]$_DFFE_PP_  (.D(_00426_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\text_in_r[115] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[116]$_DFFE_PP_  (.D(_00427_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\text_in_r[116] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[117]$_DFFE_PP_  (.D(_00428_),
    .CLK(clknet_leaf_349_clk),
    .Q(\text_in_r[117] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[118]$_DFFE_PP_  (.D(_00429_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\text_in_r[118] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[119]$_DFFE_PP_  (.D(_00430_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\text_in_r[119] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[11]$_DFFE_PP_  (.D(_00431_),
    .CLK(clknet_leaf_370_clk),
    .Q(\text_in_r[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[120]$_DFFE_PP_  (.D(_00432_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\text_in_r[120] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[121]$_DFFE_PP_  (.D(_00433_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\text_in_r[121] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[122]$_DFFE_PP_  (.D(_00434_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\text_in_r[122] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[123]$_DFFE_PP_  (.D(_00435_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\text_in_r[123] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[124]$_DFFE_PP_  (.D(_00436_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\text_in_r[124] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[125]$_DFFE_PP_  (.D(_00437_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\text_in_r[125] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[126]$_DFFE_PP_  (.D(_00438_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\text_in_r[126] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[127]$_DFFE_PP_  (.D(_00439_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\text_in_r[127] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[12]$_DFFE_PP_  (.D(_00440_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\text_in_r[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[13]$_DFFE_PP_  (.D(_00441_),
    .CLK(clknet_leaf_5_clk),
    .Q(\text_in_r[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[14]$_DFFE_PP_  (.D(_00442_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\text_in_r[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[15]$_DFFE_PP_  (.D(_00443_),
    .CLK(clknet_leaf_382_clk),
    .Q(\text_in_r[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[16]$_DFFE_PP_  (.D(_00444_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\text_in_r[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[17]$_DFFE_PP_  (.D(_00445_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\text_in_r[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[18]$_DFFE_PP_  (.D(_00446_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\text_in_r[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[19]$_DFFE_PP_  (.D(_00447_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\text_in_r[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[1]$_DFFE_PP_  (.D(_00448_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(\text_in_r[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[20]$_DFFE_PP_  (.D(_00449_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(\text_in_r[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[21]$_DFFE_PP_  (.D(_00450_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\text_in_r[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[22]$_DFFE_PP_  (.D(_00451_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\text_in_r[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[23]$_DFFE_PP_  (.D(_00452_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\text_in_r[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[24]$_DFFE_PP_  (.D(_00453_),
    .CLK(clknet_leaf_318_clk),
    .Q(\text_in_r[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[25]$_DFFE_PP_  (.D(_00454_),
    .CLK(clknet_leaf_303_clk),
    .Q(\text_in_r[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[26]$_DFFE_PP_  (.D(_00455_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\text_in_r[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[27]$_DFFE_PP_  (.D(_00456_),
    .CLK(clknet_leaf_303_clk),
    .Q(\text_in_r[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[28]$_DFFE_PP_  (.D(_00457_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\text_in_r[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[29]$_DFFE_PP_  (.D(_00458_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\text_in_r[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[2]$_DFFE_PP_  (.D(_00459_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\text_in_r[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[30]$_DFFE_PP_  (.D(_00460_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\text_in_r[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[31]$_DFFE_PP_  (.D(_00461_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(\text_in_r[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[32]$_DFFE_PP_  (.D(_00462_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(\text_in_r[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[33]$_DFFE_PP_  (.D(_00463_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(\text_in_r[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[34]$_DFFE_PP_  (.D(_00464_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(\text_in_r[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[35]$_DFFE_PP_  (.D(_00465_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(\text_in_r[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[36]$_DFFE_PP_  (.D(_00466_),
    .CLK(clknet_leaf_283_clk),
    .Q(\text_in_r[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[37]$_DFFE_PP_  (.D(_00467_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(\text_in_r[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[38]$_DFFE_PP_  (.D(_00468_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(\text_in_r[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[39]$_DFFE_PP_  (.D(_00469_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(\text_in_r[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[3]$_DFFE_PP_  (.D(_00470_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(\text_in_r[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[40]$_DFFE_PP_  (.D(_00471_),
    .CLK(clknet_leaf_207_clk),
    .Q(\text_in_r[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[41]$_DFFE_PP_  (.D(_00472_),
    .CLK(clknet_5_30__leaf_clk),
    .Q(\text_in_r[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[42]$_DFFE_PP_  (.D(_00473_),
    .CLK(clknet_leaf_206_clk),
    .Q(\text_in_r[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[43]$_DFFE_PP_  (.D(_00474_),
    .CLK(clknet_5_30__leaf_clk),
    .Q(\text_in_r[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[44]$_DFFE_PP_  (.D(_00475_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\text_in_r[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[45]$_DFFE_PP_  (.D(_00476_),
    .CLK(clknet_leaf_250_clk),
    .Q(\text_in_r[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[46]$_DFFE_PP_  (.D(_00477_),
    .CLK(clknet_leaf_205_clk),
    .Q(\text_in_r[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[47]$_DFFE_PP_  (.D(_00478_),
    .CLK(clknet_5_25__leaf_clk),
    .Q(\text_in_r[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[48]$_DFFE_PP_  (.D(_00479_),
    .CLK(clknet_5_25__leaf_clk),
    .Q(\text_in_r[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[49]$_DFFE_PP_  (.D(_00480_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\text_in_r[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[4]$_DFFE_PP_  (.D(_00481_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\text_in_r[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[50]$_DFFE_PP_  (.D(_00482_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\text_in_r[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[51]$_DFFE_PP_  (.D(_00483_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\text_in_r[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[52]$_DFFE_PP_  (.D(_00484_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\text_in_r[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[53]$_DFFE_PP_  (.D(_00485_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\text_in_r[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[54]$_DFFE_PP_  (.D(_00486_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(\text_in_r[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[55]$_DFFE_PP_  (.D(_00487_),
    .CLK(clknet_leaf_138_clk),
    .Q(\text_in_r[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[56]$_DFFE_PP_  (.D(_00488_),
    .CLK(clknet_leaf_223_clk),
    .Q(\text_in_r[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[57]$_DFFE_PP_  (.D(_00489_),
    .CLK(clknet_leaf_221_clk),
    .Q(\text_in_r[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[58]$_DFFE_PP_  (.D(_00490_),
    .CLK(clknet_5_30__leaf_clk),
    .Q(\text_in_r[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[59]$_DFFE_PP_  (.D(_00491_),
    .CLK(clknet_leaf_209_clk),
    .Q(\text_in_r[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[5]$_DFFE_PP_  (.D(_00492_),
    .CLK(clknet_leaf_352_clk),
    .Q(\text_in_r[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[60]$_DFFE_PP_  (.D(_00493_),
    .CLK(clknet_leaf_223_clk),
    .Q(\text_in_r[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[61]$_DFFE_PP_  (.D(_00494_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(\text_in_r[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[62]$_DFFE_PP_  (.D(_00495_),
    .CLK(clknet_leaf_257_clk),
    .Q(\text_in_r[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[63]$_DFFE_PP_  (.D(_00496_),
    .CLK(clknet_5_25__leaf_clk),
    .Q(\text_in_r[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[64]$_DFFE_PP_  (.D(_00497_),
    .CLK(clknet_leaf_125_clk),
    .Q(\text_in_r[64] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[65]$_DFFE_PP_  (.D(_00498_),
    .CLK(clknet_leaf_126_clk),
    .Q(\text_in_r[65] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[66]$_DFFE_PP_  (.D(_00499_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\text_in_r[66] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[67]$_DFFE_PP_  (.D(_00500_),
    .CLK(clknet_leaf_142_clk),
    .Q(\text_in_r[67] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[68]$_DFFE_PP_  (.D(_00501_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\text_in_r[68] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[69]$_DFFE_PP_  (.D(_00502_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\text_in_r[69] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[6]$_DFFE_PP_  (.D(_00503_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\text_in_r[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[70]$_DFFE_PP_  (.D(_00504_),
    .CLK(clknet_5_11__leaf_clk),
    .Q(\text_in_r[70] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[71]$_DFFE_PP_  (.D(_00505_),
    .CLK(clknet_leaf_154_clk),
    .Q(\text_in_r[71] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[72]$_DFFE_PP_  (.D(_00506_),
    .CLK(clknet_leaf_1_clk),
    .Q(\text_in_r[72] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[73]$_DFFE_PP_  (.D(_00507_),
    .CLK(clknet_leaf_423_clk),
    .Q(\text_in_r[73] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[74]$_DFFE_PP_  (.D(_00508_),
    .CLK(clknet_leaf_91_clk),
    .Q(\text_in_r[74] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[75]$_DFFE_PP_  (.D(_00509_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\text_in_r[75] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[76]$_DFFE_PP_  (.D(_00510_),
    .CLK(clknet_leaf_417_clk),
    .Q(\text_in_r[76] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[77]$_DFFE_PP_  (.D(_00511_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\text_in_r[77] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[78]$_DFFE_PP_  (.D(_00512_),
    .CLK(clknet_leaf_81_clk),
    .Q(\text_in_r[78] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[79]$_DFFE_PP_  (.D(_00513_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(\text_in_r[79] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[7]$_DFFE_PP_  (.D(_00514_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\text_in_r[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[80]$_DFFE_PP_  (.D(_00515_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(\text_in_r[80] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[81]$_DFFE_PP_  (.D(_00516_),
    .CLK(clknet_leaf_102_clk),
    .Q(\text_in_r[81] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[82]$_DFFE_PP_  (.D(_00517_),
    .CLK(clknet_leaf_102_clk),
    .Q(\text_in_r[82] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[83]$_DFFE_PP_  (.D(_00518_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(\text_in_r[83] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[84]$_DFFE_PP_  (.D(_00519_),
    .CLK(clknet_leaf_71_clk),
    .Q(\text_in_r[84] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[85]$_DFFE_PP_  (.D(_00520_),
    .CLK(clknet_leaf_81_clk),
    .Q(\text_in_r[85] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[86]$_DFFE_PP_  (.D(_00521_),
    .CLK(clknet_leaf_86_clk),
    .Q(\text_in_r[86] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[87]$_DFFE_PP_  (.D(_00522_),
    .CLK(clknet_leaf_82_clk),
    .Q(\text_in_r[87] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[88]$_DFFE_PP_  (.D(_00523_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\text_in_r[88] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[89]$_DFFE_PP_  (.D(_00524_),
    .CLK(clknet_leaf_111_clk),
    .Q(\text_in_r[89] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[8]$_DFFE_PP_  (.D(_00525_),
    .CLK(clknet_leaf_369_clk),
    .Q(\text_in_r[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[90]$_DFFE_PP_  (.D(_00526_),
    .CLK(clknet_leaf_111_clk),
    .Q(\text_in_r[90] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[91]$_DFFE_PP_  (.D(_00527_),
    .CLK(clknet_leaf_141_clk),
    .Q(\text_in_r[91] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[92]$_DFFE_PP_  (.D(_00528_),
    .CLK(clknet_5_11__leaf_clk),
    .Q(\text_in_r[92] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[93]$_DFFE_PP_  (.D(_00529_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\text_in_r[93] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[94]$_DFFE_PP_  (.D(_00530_),
    .CLK(clknet_leaf_138_clk),
    .Q(\text_in_r[94] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[95]$_DFFE_PP_  (.D(_00531_),
    .CLK(clknet_leaf_138_clk),
    .Q(\text_in_r[95] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[96]$_DFFE_PP_  (.D(_00532_),
    .CLK(clknet_leaf_139_clk),
    .Q(\text_in_r[96] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[97]$_DFFE_PP_  (.D(_00533_),
    .CLK(clknet_leaf_143_clk),
    .Q(\text_in_r[97] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[98]$_DFFE_PP_  (.D(_00534_),
    .CLK(clknet_5_11__leaf_clk),
    .Q(\text_in_r[98] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[99]$_DFFE_PP_  (.D(_00535_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\text_in_r[99] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_in_r[9]$_DFFE_PP_  (.D(_00536_),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\text_in_r[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[0]$_DFF_P_  (.D(_00265_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(net260));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[100]$_DFF_P_  (.D(_00165_),
    .CLK(clknet_leaf_167_clk),
    .Q(net261));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[101]$_DFF_P_  (.D(_00166_),
    .CLK(clknet_leaf_358_clk),
    .Q(net262));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[102]$_DFF_P_  (.D(_00167_),
    .CLK(clknet_leaf_355_clk),
    .Q(net263));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[103]$_DFF_P_  (.D(_00168_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(net264));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[104]$_DFF_P_  (.D(_00169_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(net265));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[105]$_DFF_P_  (.D(_00170_),
    .CLK(clknet_leaf_178_clk),
    .Q(net266));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[106]$_DFF_P_  (.D(_00171_),
    .CLK(clknet_leaf_185_clk),
    .Q(net267));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[107]$_DFF_P_  (.D(_00172_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(net268));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[108]$_DFF_P_  (.D(_00173_),
    .CLK(clknet_leaf_273_clk),
    .Q(net269));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[109]$_DFF_P_  (.D(_00174_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(net270));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[10]$_DFF_P_  (.D(_00195_),
    .CLK(clknet_leaf_7_clk),
    .Q(net271));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[110]$_DFF_P_  (.D(_00175_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(net272));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[111]$_DFF_P_  (.D(_00176_),
    .CLK(clknet_leaf_168_clk),
    .Q(net273));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[112]$_DFF_P_  (.D(_00177_),
    .CLK(clknet_leaf_166_clk),
    .Q(net274));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[113]$_DFF_P_  (.D(_00178_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(net275));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[114]$_DFF_P_  (.D(_00179_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(net276));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[115]$_DFF_P_  (.D(_00180_),
    .CLK(clknet_leaf_166_clk),
    .Q(net277));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[116]$_DFF_P_  (.D(_00181_),
    .CLK(clknet_leaf_355_clk),
    .Q(net278));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[117]$_DFF_P_  (.D(_00182_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(net279));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[118]$_DFF_P_  (.D(_00183_),
    .CLK(clknet_leaf_25_clk),
    .Q(net280));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[119]$_DFF_P_  (.D(_00184_),
    .CLK(clknet_leaf_168_clk),
    .Q(net281));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[11]$_DFF_P_  (.D(_00196_),
    .CLK(clknet_leaf_376_clk),
    .Q(net282));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[120]$_DFF_P_  (.D(_00185_),
    .CLK(clknet_leaf_169_clk),
    .Q(net283));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[121]$_DFF_P_  (.D(_00186_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(net284));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[122]$_DFF_P_  (.D(_00187_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(net285));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[123]$_DFF_P_  (.D(_00188_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(net286));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[124]$_DFF_P_  (.D(_00189_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(net287));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[125]$_DFF_P_  (.D(_00190_),
    .CLK(clknet_leaf_270_clk),
    .Q(net288));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[126]$_DFF_P_  (.D(_00191_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(net289));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[127]$_DFF_P_  (.D(_00192_),
    .CLK(clknet_leaf_169_clk),
    .Q(net290));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[12]$_DFF_P_  (.D(_00197_),
    .CLK(clknet_5_0__leaf_clk),
    .Q(net291));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[13]$_DFF_P_  (.D(_00198_),
    .CLK(clknet_leaf_7_clk),
    .Q(net292));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[14]$_DFF_P_  (.D(_00199_),
    .CLK(clknet_leaf_29_clk),
    .Q(net293));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[15]$_DFF_P_  (.D(_00200_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(net294));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[16]$_DFF_P_  (.D(_00201_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(net295));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[17]$_DFF_P_  (.D(_00202_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(net296));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[18]$_DFF_P_  (.D(_00203_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(net297));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[19]$_DFF_P_  (.D(_00204_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(net298));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[1]$_DFF_P_  (.D(_00266_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(net299));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[20]$_DFF_P_  (.D(_00205_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(net300));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[21]$_DFF_P_  (.D(_00206_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(net301));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[22]$_DFF_P_  (.D(_00207_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(net302));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[23]$_DFF_P_  (.D(_00208_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(net303));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[24]$_DFF_P_  (.D(_00209_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(net304));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[25]$_DFF_P_  (.D(_00210_),
    .CLK(clknet_leaf_315_clk),
    .Q(net305));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[26]$_DFF_P_  (.D(_00211_),
    .CLK(clknet_leaf_318_clk),
    .Q(net306));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[27]$_DFF_P_  (.D(_00212_),
    .CLK(clknet_5_21__leaf_clk),
    .Q(net307));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[28]$_DFF_P_  (.D(_00213_),
    .CLK(clknet_5_20__leaf_clk),
    .Q(net308));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[29]$_DFF_P_  (.D(_00214_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(net309));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[2]$_DFF_P_  (.D(_00267_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(net310));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[30]$_DFF_P_  (.D(_00215_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(net311));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[31]$_DFF_P_  (.D(_00216_),
    .CLK(clknet_leaf_313_clk),
    .Q(net312));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[32]$_DFF_P_  (.D(_00217_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(net313));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[33]$_DFF_P_  (.D(_00218_),
    .CLK(clknet_5_30__leaf_clk),
    .Q(net314));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[34]$_DFF_P_  (.D(_00219_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(net315));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[35]$_DFF_P_  (.D(_00220_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(net316));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[36]$_DFF_P_  (.D(_00221_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(net317));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[37]$_DFF_P_  (.D(_00222_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(net318));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[38]$_DFF_P_  (.D(_00223_),
    .CLK(clknet_5_28__leaf_clk),
    .Q(net319));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[39]$_DFF_P_  (.D(_00224_),
    .CLK(clknet_leaf_283_clk),
    .Q(net320));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[3]$_DFF_P_  (.D(_00268_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(net321));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[40]$_DFF_P_  (.D(_00225_),
    .CLK(clknet_5_27__leaf_clk),
    .Q(net322));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[41]$_DFF_P_  (.D(_00226_),
    .CLK(clknet_leaf_206_clk),
    .Q(net323));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[42]$_DFF_P_  (.D(_00227_),
    .CLK(clknet_leaf_205_clk),
    .Q(net324));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[43]$_DFF_P_  (.D(_00228_),
    .CLK(clknet_5_30__leaf_clk),
    .Q(net325));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[44]$_DFF_P_  (.D(_00229_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(net326));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[45]$_DFF_P_  (.D(_00230_),
    .CLK(clknet_5_25__leaf_clk),
    .Q(net327));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[46]$_DFF_P_  (.D(_00231_),
    .CLK(clknet_leaf_241_clk),
    .Q(net328));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[47]$_DFF_P_  (.D(_00232_),
    .CLK(clknet_leaf_241_clk),
    .Q(net329));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[48]$_DFF_P_  (.D(_00233_),
    .CLK(clknet_leaf_249_clk),
    .Q(net330));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[49]$_DFF_P_  (.D(_00234_),
    .CLK(clknet_leaf_254_clk),
    .Q(net331));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[4]$_DFF_P_  (.D(_00269_),
    .CLK(clknet_5_17__leaf_clk),
    .Q(net332));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[50]$_DFF_P_  (.D(_00235_),
    .CLK(clknet_leaf_185_clk),
    .Q(net333));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[51]$_DFF_P_  (.D(_00236_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(net334));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[52]$_DFF_P_  (.D(_00237_),
    .CLK(clknet_leaf_252_clk),
    .Q(net335));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[53]$_DFF_P_  (.D(_00238_),
    .CLK(clknet_leaf_254_clk),
    .Q(net336));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[54]$_DFF_P_  (.D(_00239_),
    .CLK(clknet_leaf_152_clk),
    .Q(net337));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[55]$_DFF_P_  (.D(_00240_),
    .CLK(clknet_leaf_252_clk),
    .Q(net338));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[56]$_DFF_P_  (.D(_00241_),
    .CLK(clknet_leaf_239_clk),
    .Q(net339));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[57]$_DFF_P_  (.D(_00242_),
    .CLK(clknet_leaf_239_clk),
    .Q(net340));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[58]$_DFF_P_  (.D(_00243_),
    .CLK(clknet_leaf_209_clk),
    .Q(net341));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[59]$_DFF_P_  (.D(_00244_),
    .CLK(clknet_5_30__leaf_clk),
    .Q(net342));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[5]$_DFF_P_  (.D(_00270_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(net343));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[60]$_DFF_P_  (.D(_00245_),
    .CLK(clknet_leaf_231_clk),
    .Q(net344));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[61]$_DFF_P_  (.D(_00246_),
    .CLK(clknet_5_29__leaf_clk),
    .Q(net345));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[62]$_DFF_P_  (.D(_00247_),
    .CLK(clknet_leaf_257_clk),
    .Q(net346));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[63]$_DFF_P_  (.D(_00248_),
    .CLK(clknet_leaf_250_clk),
    .Q(net347));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[64]$_DFF_P_  (.D(_00249_),
    .CLK(clknet_leaf_125_clk),
    .Q(net348));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[65]$_DFF_P_  (.D(_00250_),
    .CLK(clknet_5_11__leaf_clk),
    .Q(net349));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[66]$_DFF_P_  (.D(_00251_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(net350));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[67]$_DFF_P_  (.D(_00252_),
    .CLK(clknet_5_11__leaf_clk),
    .Q(net351));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[68]$_DFF_P_  (.D(_00253_),
    .CLK(clknet_leaf_57_clk),
    .Q(net352));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[69]$_DFF_P_  (.D(_00254_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(net353));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[6]$_DFF_P_  (.D(_00271_),
    .CLK(clknet_leaf_352_clk),
    .Q(net354));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[70]$_DFF_P_  (.D(_00255_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(net355));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[71]$_DFF_P_  (.D(_00256_),
    .CLK(clknet_leaf_138_clk),
    .Q(net356));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[72]$_DFF_P_  (.D(_00257_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(net357));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[73]$_DFF_P_  (.D(_00258_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(net358));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[74]$_DFF_P_  (.D(_00259_),
    .CLK(clknet_leaf_77_clk),
    .Q(net359));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[75]$_DFF_P_  (.D(_00260_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(net360));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[76]$_DFF_P_  (.D(_00261_),
    .CLK(clknet_leaf_417_clk),
    .Q(net361));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[77]$_DFF_P_  (.D(_00262_),
    .CLK(clknet_leaf_424_clk),
    .Q(net362));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[78]$_DFF_P_  (.D(_00263_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(net363));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[79]$_DFF_P_  (.D(_00264_),
    .CLK(clknet_leaf_71_clk),
    .Q(net364));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[7]$_DFF_P_  (.D(_00272_),
    .CLK(clknet_5_16__leaf_clk),
    .Q(net365));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[80]$_DFF_P_  (.D(_00273_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(net366));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[81]$_DFF_P_  (.D(_00274_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(net367));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[82]$_DFF_P_  (.D(_00275_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(net368));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[83]$_DFF_P_  (.D(_00276_),
    .CLK(clknet_leaf_82_clk),
    .Q(net369));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[84]$_DFF_P_  (.D(_00277_),
    .CLK(clknet_leaf_61_clk),
    .Q(net370));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[85]$_DFF_P_  (.D(_00278_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(net371));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[86]$_DFF_P_  (.D(_00279_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(net372));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[87]$_DFF_P_  (.D(_00280_),
    .CLK(clknet_leaf_61_clk),
    .Q(net373));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[88]$_DFF_P_  (.D(_00281_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(net374));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[89]$_DFF_P_  (.D(_00282_),
    .CLK(clknet_leaf_127_clk),
    .Q(net375));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[8]$_DFF_P_  (.D(_00193_),
    .CLK(clknet_leaf_377_clk),
    .Q(net376));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[90]$_DFF_P_  (.D(_00283_),
    .CLK(clknet_5_10__leaf_clk),
    .Q(net377));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[91]$_DFF_P_  (.D(_00284_),
    .CLK(clknet_leaf_141_clk),
    .Q(net378));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[92]$_DFF_P_  (.D(_00285_),
    .CLK(clknet_5_11__leaf_clk),
    .Q(net379));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[93]$_DFF_P_  (.D(_00286_),
    .CLK(clknet_leaf_57_clk),
    .Q(net380));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[94]$_DFF_P_  (.D(_00287_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(net381));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[95]$_DFF_P_  (.D(_00288_),
    .CLK(clknet_leaf_58_clk),
    .Q(net382));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[96]$_DFF_P_  (.D(_00161_),
    .CLK(clknet_leaf_150_clk),
    .Q(net383));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[97]$_DFF_P_  (.D(_00162_),
    .CLK(clknet_leaf_178_clk),
    .Q(net384));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[98]$_DFF_P_  (.D(_00163_),
    .CLK(clknet_leaf_150_clk),
    .Q(net385));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[99]$_DFF_P_  (.D(_00164_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(net386));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \text_out[9]$_DFF_P_  (.D(_00194_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(net387));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[24]$_SDFF_PP1_  (.D(_00537_),
    .CLK(clknet_leaf_42_clk),
    .Q(\u0.r0.out[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[25]$_SDFF_PP0_  (.D(_00538_),
    .CLK(clknet_leaf_45_clk),
    .Q(\u0.r0.out[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[26]$_SDFF_PP0_  (.D(_00539_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.r0.out[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[27]$_SDFF_PP0_  (.D(_00540_),
    .CLK(clknet_leaf_53_clk),
    .Q(\u0.r0.out[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[28]$_SDFF_PP0_  (.D(_00541_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.r0.out[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[29]$_SDFF_PP0_  (.D(_00542_),
    .CLK(clknet_leaf_35_clk),
    .Q(\u0.r0.out[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[30]$_SDFF_PP0_  (.D(_00543_),
    .CLK(clknet_leaf_35_clk),
    .Q(\u0.r0.out[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.out[31]$_SDFF_PP0_  (.D(_00544_),
    .CLK(clknet_leaf_45_clk),
    .Q(\u0.r0.out[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.rcnt[0]$_SDFF_PP0_  (.D(_00545_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.r0.rcnt[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.rcnt[1]$_SDFF_PP0_  (.D(_00546_),
    .CLK(clknet_leaf_39_clk),
    .Q(\u0.r0.rcnt[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.rcnt[2]$_SDFF_PP0_  (.D(_00547_),
    .CLK(clknet_leaf_42_clk),
    .Q(\u0.r0.rcnt[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.r0.rcnt[3]$_SDFF_PP0_  (.D(_00548_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.r0.rcnt[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[0]$_DFF_P_  (.D(_00000_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.subword[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[1]$_DFF_P_  (.D(_00001_),
    .CLK(clknet_leaf_376_clk),
    .Q(\u0.subword[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[2]$_DFF_P_  (.D(_00002_),
    .CLK(clknet_leaf_394_clk),
    .Q(\u0.subword[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[3]$_DFF_P_  (.D(_00003_),
    .CLK(clknet_leaf_376_clk),
    .Q(\u0.subword[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[4]$_DFF_P_  (.D(_00004_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.subword[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[5]$_DFF_P_  (.D(_00005_),
    .CLK(clknet_leaf_390_clk),
    .Q(\u0.subword[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[6]$_DFF_P_  (.D(_00006_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\u0.subword[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u0.d[7]$_DFF_P_  (.D(_00007_),
    .CLK(clknet_leaf_36_clk),
    .Q(\u0.subword[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[0]$_DFF_P_  (.D(_00008_),
    .CLK(clknet_leaf_417_clk),
    .Q(\u0.subword[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[1]$_DFF_P_  (.D(_00009_),
    .CLK(clknet_leaf_415_clk),
    .Q(\u0.subword[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[2]$_DFF_P_  (.D(_00010_),
    .CLK(clknet_leaf_410_clk),
    .Q(\u0.subword[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[3]$_DFF_P_  (.D(_00011_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\u0.subword[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[4]$_DFF_P_  (.D(_00012_),
    .CLK(clknet_leaf_411_clk),
    .Q(\u0.subword[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[5]$_DFF_P_  (.D(_00013_),
    .CLK(clknet_leaf_412_clk),
    .Q(\u0.subword[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[6]$_DFF_P_  (.D(_00014_),
    .CLK(clknet_leaf_411_clk),
    .Q(\u0.subword[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u1.d[7]$_DFF_P_  (.D(_00015_),
    .CLK(clknet_leaf_410_clk),
    .Q(\u0.subword[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[0]$_DFF_P_  (.D(_00016_),
    .CLK(clknet_leaf_431_clk),
    .Q(\u0.subword[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[1]$_DFF_P_  (.D(_00017_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.subword[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[2]$_DFF_P_  (.D(_00018_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.subword[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[3]$_DFF_P_  (.D(_00019_),
    .CLK(clknet_leaf_431_clk),
    .Q(\u0.subword[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[4]$_DFF_P_  (.D(_00020_),
    .CLK(clknet_leaf_1_clk),
    .Q(\u0.subword[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[5]$_DFF_P_  (.D(_00021_),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\u0.subword[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[6]$_DFF_P_  (.D(_00022_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\u0.subword[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u2.d[7]$_DFF_P_  (.D(_00023_),
    .CLK(clknet_leaf_29_clk),
    .Q(\u0.subword[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[0]$_DFF_P_  (.D(_00024_),
    .CLK(clknet_leaf_378_clk),
    .Q(\u0.subword[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[1]$_DFF_P_  (.D(_00025_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\u0.subword[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[2]$_DFF_P_  (.D(_00026_),
    .CLK(clknet_leaf_370_clk),
    .Q(\u0.subword[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[3]$_DFF_P_  (.D(_00027_),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\u0.subword[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[4]$_DFF_P_  (.D(_00028_),
    .CLK(clknet_leaf_389_clk),
    .Q(\u0.subword[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[5]$_DFF_P_  (.D(_00029_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\u0.subword[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[6]$_DFF_P_  (.D(_00030_),
    .CLK(clknet_leaf_382_clk),
    .Q(\u0.subword[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.u3.d[7]$_DFF_P_  (.D(_00031_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\u0.subword[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][0]$_DFF_P_  (.D(_00289_),
    .CLK(clknet_leaf_152_clk),
    .Q(\u0.w[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][10]$_DFF_P_  (.D(_00290_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.w[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][11]$_DFF_P_  (.D(_00291_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.w[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][12]$_DFF_P_  (.D(_00292_),
    .CLK(clknet_leaf_413_clk),
    .Q(\u0.w[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][13]$_DFF_P_  (.D(_00293_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][14]$_DFF_P_  (.D(_00294_),
    .CLK(clknet_leaf_22_clk),
    .Q(\u0.w[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][15]$_DFF_P_  (.D(_00295_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\u0.w[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][16]$_DFF_P_  (.D(_00296_),
    .CLK(clknet_leaf_75_clk),
    .Q(\u0.w[0][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][17]$_DFF_P_  (.D(_00297_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.w[0][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][18]$_DFF_P_  (.D(_00298_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.w[0][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][19]$_DFF_P_  (.D(_00299_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.w[0][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][1]$_DFF_P_  (.D(_00300_),
    .CLK(clknet_leaf_160_clk),
    .Q(\u0.w[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][20]$_DFF_P_  (.D(_00301_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\u0.w[0][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][21]$_DFF_P_  (.D(_00302_),
    .CLK(clknet_leaf_28_clk),
    .Q(\u0.w[0][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][22]$_DFF_P_  (.D(_00303_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.w[0][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][23]$_DFF_P_  (.D(_00304_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\u0.w[0][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][24]$_DFF_P_  (.D(_00305_),
    .CLK(clknet_leaf_43_clk),
    .Q(\u0.w[0][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][25]$_DFF_P_  (.D(_00306_),
    .CLK(clknet_leaf_54_clk),
    .Q(\u0.w[0][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][26]$_DFF_P_  (.D(_00307_),
    .CLK(clknet_leaf_160_clk),
    .Q(\u0.w[0][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][27]$_DFF_P_  (.D(_00308_),
    .CLK(clknet_leaf_159_clk),
    .Q(\u0.w[0][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][28]$_DFF_P_  (.D(_00309_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\u0.w[0][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][29]$_DFF_P_  (.D(_00310_),
    .CLK(clknet_leaf_37_clk),
    .Q(\u0.w[0][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][2]$_DFF_P_  (.D(_00311_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\u0.w[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][30]$_DFF_P_  (.D(_00312_),
    .CLK(clknet_leaf_36_clk),
    .Q(\u0.w[0][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][31]$_DFF_P_  (.D(_00313_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.w[0][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][3]$_DFF_P_  (.D(_00314_),
    .CLK(clknet_leaf_154_clk),
    .Q(\u0.w[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][4]$_DFF_P_  (.D(_00315_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\u0.w[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][5]$_DFF_P_  (.D(_00316_),
    .CLK(clknet_leaf_363_clk),
    .Q(\u0.w[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][6]$_DFF_P_  (.D(_00317_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\u0.w[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][7]$_DFF_P_  (.D(_00318_),
    .CLK(clknet_leaf_354_clk),
    .Q(\u0.w[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][8]$_DFF_P_  (.D(_00319_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.w[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[0][9]$_DFF_P_  (.D(_00320_),
    .CLK(clknet_leaf_425_clk),
    .Q(\u0.w[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][0]$_DFF_P_  (.D(_00321_),
    .CLK(clknet_leaf_143_clk),
    .Q(\u0.w[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][10]$_DFF_P_  (.D(_00322_),
    .CLK(clknet_leaf_15_clk),
    .Q(\u0.w[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][11]$_DFF_P_  (.D(_00323_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.w[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][12]$_DFF_P_  (.D(_00324_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\u0.w[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][13]$_DFF_P_  (.D(_00325_),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\u0.w[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][14]$_DFF_P_  (.D(_00326_),
    .CLK(clknet_leaf_25_clk),
    .Q(\u0.w[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][15]$_DFF_P_  (.D(_00327_),
    .CLK(clknet_leaf_49_clk),
    .Q(\u0.w[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][16]$_DFF_P_  (.D(_00328_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.w[1][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][17]$_DFF_P_  (.D(_00329_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.w[1][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][18]$_DFF_P_  (.D(_00330_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.w[1][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][19]$_DFF_P_  (.D(_00331_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\u0.w[1][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][1]$_DFF_P_  (.D(_00332_),
    .CLK(clknet_leaf_142_clk),
    .Q(\u0.w[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][20]$_DFF_P_  (.D(_00333_),
    .CLK(clknet_leaf_19_clk),
    .Q(\u0.w[1][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][21]$_DFF_P_  (.D(_00334_),
    .CLK(clknet_leaf_21_clk),
    .Q(\u0.w[1][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][22]$_DFF_P_  (.D(_00335_),
    .CLK(clknet_leaf_11_clk),
    .Q(\u0.w[1][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][23]$_DFF_P_  (.D(_00336_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\u0.w[1][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][24]$_DFF_P_  (.D(_00337_),
    .CLK(clknet_leaf_77_clk),
    .Q(\u0.w[1][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][25]$_DFF_P_  (.D(_00338_),
    .CLK(clknet_leaf_49_clk),
    .Q(\u0.w[1][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][26]$_DFF_P_  (.D(_00339_),
    .CLK(clknet_5_9__leaf_clk),
    .Q(\u0.w[1][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][27]$_DFF_P_  (.D(_00340_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\u0.w[1][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][28]$_DFF_P_  (.D(_00341_),
    .CLK(clknet_leaf_22_clk),
    .Q(\u0.w[1][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][29]$_DFF_P_  (.D(_00342_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\u0.w[1][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][2]$_DFF_P_  (.D(_00343_),
    .CLK(clknet_leaf_144_clk),
    .Q(\u0.w[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][30]$_DFF_P_  (.D(_00344_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.w[1][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][31]$_DFF_P_  (.D(_00345_),
    .CLK(clknet_leaf_54_clk),
    .Q(\u0.w[1][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][3]$_DFF_P_  (.D(_00346_),
    .CLK(clknet_leaf_139_clk),
    .Q(\u0.w[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][4]$_DFF_P_  (.D(_00347_),
    .CLK(clknet_5_12__leaf_clk),
    .Q(\u0.w[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][5]$_DFF_P_  (.D(_00348_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\u0.w[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][6]$_DFF_P_  (.D(_00349_),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\u0.w[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][7]$_DFF_P_  (.D(_00350_),
    .CLK(clknet_leaf_354_clk),
    .Q(\u0.w[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][8]$_DFF_P_  (.D(_00351_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.w[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[1][9]$_DFF_P_  (.D(_00352_),
    .CLK(clknet_leaf_425_clk),
    .Q(\u0.w[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][0]$_DFF_P_  (.D(_00353_),
    .CLK(clknet_leaf_161_clk),
    .Q(\u0.w[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][10]$_DFF_P_  (.D(_00354_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.w[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][11]$_DFF_P_  (.D(_00355_),
    .CLK(clknet_leaf_424_clk),
    .Q(\u0.w[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][12]$_DFF_P_  (.D(_00356_),
    .CLK(clknet_leaf_413_clk),
    .Q(\u0.w[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][13]$_DFF_P_  (.D(_00357_),
    .CLK(clknet_leaf_0_clk),
    .Q(\u0.w[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][14]$_DFF_P_  (.D(_00358_),
    .CLK(clknet_leaf_32_clk),
    .Q(\u0.w[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][15]$_DFF_P_  (.D(_00359_),
    .CLK(clknet_leaf_49_clk),
    .Q(\u0.w[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][16]$_DFF_P_  (.D(_00360_),
    .CLK(clknet_leaf_75_clk),
    .Q(\u0.w[2][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][17]$_DFF_P_  (.D(_00361_),
    .CLK(clknet_leaf_15_clk),
    .Q(\u0.w[2][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][18]$_DFF_P_  (.D(_00362_),
    .CLK(clknet_leaf_19_clk),
    .Q(\u0.w[2][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][19]$_DFF_P_  (.D(_00363_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\u0.w[2][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][1]$_DFF_P_  (.D(_00364_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.w[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][20]$_DFF_P_  (.D(_00365_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\u0.w[2][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][21]$_DFF_P_  (.D(_00366_),
    .CLK(clknet_leaf_30_clk),
    .Q(\u0.w[2][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][22]$_DFF_P_  (.D(_00367_),
    .CLK(clknet_leaf_28_clk),
    .Q(\u0.w[2][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][23]$_DFF_P_  (.D(_00368_),
    .CLK(clknet_leaf_21_clk),
    .Q(\u0.w[2][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][24]$_DFF_P_  (.D(_00369_),
    .CLK(clknet_leaf_167_clk),
    .Q(\u0.w[2][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][25]$_DFF_P_  (.D(_00370_),
    .CLK(clknet_leaf_53_clk),
    .Q(\u0.w[2][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][26]$_DFF_P_  (.D(_00371_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.w[2][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][27]$_DFF_P_  (.D(_00372_),
    .CLK(clknet_leaf_159_clk),
    .Q(\u0.w[2][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][28]$_DFF_P_  (.D(_00373_),
    .CLK(clknet_leaf_32_clk),
    .Q(\u0.w[2][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][29]$_DFF_P_  (.D(_00374_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\u0.w[2][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][2]$_DFF_P_  (.D(_00375_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.w[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][30]$_DFF_P_  (.D(_00376_),
    .CLK(clknet_leaf_37_clk),
    .Q(\u0.w[2][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][31]$_DFF_P_  (.D(_00377_),
    .CLK(clknet_leaf_43_clk),
    .Q(\u0.w[2][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][3]$_DFF_P_  (.D(_00378_),
    .CLK(clknet_leaf_161_clk),
    .Q(\u0.w[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][4]$_DFF_P_  (.D(_00379_),
    .CLK(clknet_5_13__leaf_clk),
    .Q(\u0.w[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][5]$_DFF_P_  (.D(_00380_),
    .CLK(clknet_leaf_363_clk),
    .Q(\u0.w[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][6]$_DFF_P_  (.D(_00381_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\u0.w[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][7]$_DFF_P_  (.D(_00382_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\u0.w[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][8]$_DFF_P_  (.D(_00383_),
    .CLK(clknet_5_3__leaf_clk),
    .Q(\u0.w[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[2][9]$_DFF_P_  (.D(_00384_),
    .CLK(clknet_leaf_423_clk),
    .Q(\u0.w[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][0]$_DFF_P_  (.D(net20811),
    .CLK(clknet_leaf_376_clk),
    .Q(\u0.tmp_w[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][10]$_DFF_P_  (.D(_07622_),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\u0.tmp_w[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][11]$_DFF_P_  (.D(net20578),
    .CLK(clknet_leaf_415_clk),
    .Q(\u0.tmp_w[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][12]$_DFF_P_  (.D(_07639_),
    .CLK(clknet_leaf_412_clk),
    .Q(\u0.tmp_w[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][13]$_DFF_P_  (.D(net20712),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\u0.tmp_w[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][14]$_DFF_P_  (.D(net20708),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\u0.tmp_w[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][15]$_DFF_P_  (.D(net20847),
    .CLK(clknet_leaf_30_clk),
    .Q(\u0.tmp_w[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][16]$_DFF_P_  (.D(net20832),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\u0.tmp_w[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][17]$_DFF_P_  (.D(net20835),
    .CLK(clknet_leaf_399_clk),
    .Q(\u0.tmp_w[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][18]$_DFF_P_  (.D(net20779),
    .CLK(clknet_leaf_394_clk),
    .Q(\u0.tmp_w[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][19]$_DFF_P_  (.D(_07330_),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\u0.tmp_w[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][1]$_DFF_P_  (.D(net20818),
    .CLK(clknet_leaf_378_clk),
    .Q(\u0.tmp_w[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][20]$_DFF_P_  (.D(net20781),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\u0.tmp_w[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][21]$_DFF_P_  (.D(net20788),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\u0.tmp_w[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][22]$_DFF_P_  (.D(_07666_),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\u0.tmp_w[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][23]$_DFF_P_  (.D(net20845),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\u0.tmp_w[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][24]$_DFF_P_  (.D(net20471),
    .CLK(clknet_5_20__leaf_clk),
    .Q(\u0.tmp_w[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][25]$_DFF_P_  (.D(net20474),
    .CLK(clknet_5_16__leaf_clk),
    .Q(\u0.tmp_w[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][26]$_DFF_P_  (.D(net20810),
    .CLK(clknet_leaf_385_clk),
    .Q(\u0.tmp_w[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][27]$_DFF_P_  (.D(_07706_),
    .CLK(clknet_leaf_389_clk),
    .Q(\u0.tmp_w[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][28]$_DFF_P_  (.D(net20577),
    .CLK(clknet_5_22__leaf_clk),
    .Q(\u0.tmp_w[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][29]$_DFF_P_  (.D(_07727_),
    .CLK(clknet_leaf_390_clk),
    .Q(\u0.tmp_w[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][2]$_DFF_P_  (.D(net20767),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\u0.tmp_w[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][30]$_DFF_P_  (.D(net20838),
    .CLK(clknet_leaf_385_clk),
    .Q(\u0.tmp_w[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][31]$_DFF_P_  (.D(_00399_),
    .CLK(clknet_leaf_313_clk),
    .Q(\u0.tmp_w[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][3]$_DFF_P_  (.D(net20593),
    .CLK(clknet_leaf_372_clk),
    .Q(\u0.tmp_w[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][4]$_DFF_P_  (.D(net20860),
    .CLK(clknet_5_5__leaf_clk),
    .Q(\u0.tmp_w[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][5]$_DFF_P_  (.D(net20756),
    .CLK(clknet_leaf_372_clk),
    .Q(\u0.tmp_w[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][6]$_DFF_P_  (.D(net20858),
    .CLK(clknet_leaf_369_clk),
    .Q(\u0.tmp_w[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][7]$_DFF_P_  (.D(net20857),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\u0.tmp_w[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][8]$_DFF_P_  (.D(net20821),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\u0.tmp_w[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \u0.w[3][9]$_DFF_P_  (.D(net20831),
    .CLK(clknet_5_0__leaf_clk),
    .Q(\u0.tmp_w[9] ));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Right_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Right_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Right_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Right_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Right_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Right_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Right_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Right_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Right_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Right_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Right_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Right_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Right_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Right_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Right_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Right_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Right_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Right_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Right_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Right_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Right_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Right_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Right_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Right_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Right_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Right_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Right_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Right_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Right_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Right_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Right_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Right_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Right_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Right_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Right_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Right_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Right_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Right_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Right_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Right_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Right_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Right_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Right_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Right_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Right_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Right_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Right_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Right_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Right_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Right_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_371 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_372 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_373 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_374 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_375 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_376 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_377 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_378 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_379 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_380 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_381 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_382 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_383 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_384 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_385 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_386 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_387 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_388 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_389 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_390 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_391 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_392 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_393 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_394 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_395 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_396 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_397 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_398 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_399 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_400 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_401 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_402 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_403 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_404 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_405 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_406 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_407 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_408 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_409 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_410 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_411 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_412 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_413 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_414 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_415 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_416 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_417 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_418 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_419 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_420 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_421 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_422 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_423 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_424 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_425 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_426 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_427 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_428 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_429 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_430 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_431 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_432 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_433 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_434 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_435 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_436 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_437 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_438 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_439 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_440 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Left_441 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Left_442 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Left_443 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Left_444 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Left_445 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Left_446 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Left_447 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Left_448 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Left_449 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Left_450 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Left_451 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Left_452 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Left_453 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Left_454 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Left_455 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Left_456 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Left_457 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Left_458 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Left_459 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Left_460 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Left_461 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Left_462 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Left_463 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Left_464 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Left_465 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Left_466 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Left_467 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Left_468 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Left_469 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Left_470 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Left_471 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Left_472 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Left_473 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Left_474 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Left_475 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Left_476 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Left_477 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Left_478 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Left_479 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Left_480 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Left_481 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Left_482 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Left_483 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Left_484 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Left_485 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Left_486 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Left_487 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Left_488 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Left_489 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Left_490 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Left_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17799 (.I(_01093_),
    .Z(net17799));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17802 (.I(_01064_),
    .Z(net17802));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17774 (.I(_01780_),
    .Z(net17774));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17765 (.I(_01837_),
    .Z(net17765));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17772 (.I(_01790_),
    .Z(net17772));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17767 (.I(_01820_),
    .Z(net17767));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17773 (.I(_01780_),
    .Z(net17773));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17778 (.I(_01722_),
    .Z(net17778));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17770 (.I(_01797_),
    .Z(net17770));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17771 (.I(_01790_),
    .Z(net17771));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17784 (.I(_01698_),
    .Z(net17784));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17776 (.I(_01763_),
    .Z(net17776));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17858 (.I(_14536_),
    .Z(net17858));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17780 (.I(_01719_),
    .Z(net17780));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17850 (.I(_14587_),
    .Z(net17850));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18014 (.I(_06955_),
    .Z(net18014));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17814 (.I(_00940_),
    .Z(net17814));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17781 (.I(_01716_),
    .Z(net17781));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17789 (.I(_01269_),
    .Z(net17789));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17782 (.I(_01699_),
    .Z(net17782));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18240 (.I(_14435_),
    .Z(net18240));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place18178 (.I(_00995_),
    .Z(net18178));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17783 (.I(_01698_),
    .Z(net17783));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17786 (.I(_01673_),
    .Z(net17786));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17788 (.I(_01347_),
    .Z(net17788));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17810 (.I(_00990_),
    .Z(net17810));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17791 (.I(_01252_),
    .Z(net17791));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17816 (.I(_00940_),
    .Z(net17816));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17817 (.I(_00940_),
    .Z(net17817));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17805 (.I(_01028_),
    .Z(net17805));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17809 (.I(_01020_),
    .Z(net17809));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17796 (.I(_01146_),
    .Z(net17796));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17797 (.I(_01133_),
    .Z(net17797));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17798 (.I(_01112_),
    .Z(net17798));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17801 (.I(_01064_),
    .Z(net17801));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17815 (.I(net17814),
    .Z(net17815));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17807 (.I(_01025_),
    .Z(net17807));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17804 (.I(_01040_),
    .Z(net17804));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18194 (.I(net18189),
    .Z(net18194));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17812 (.I(_00979_),
    .Z(net17812));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17806 (.I(_01025_),
    .Z(net17806));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17811 (.I(_00990_),
    .Z(net17811));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17813 (.I(_00950_),
    .Z(net17813));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18012 (.I(_06958_),
    .Z(net18012));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18298 (.I(_12982_),
    .Z(net18298));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17988 (.I(_15936_[0]),
    .Z(net17988));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18001 (.I(_15709_[0]),
    .Z(net18001));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17828 (.I(_15383_),
    .Z(net17828));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18438 (.I(_06929_),
    .Z(net18438));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18310 (.I(_12919_),
    .Z(net18310));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18309 (.I(_12919_),
    .Z(net18309));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17989 (.I(_15933_[0]),
    .Z(net17989));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18292 (.I(net18291),
    .Z(net18292));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18297 (.I(net18296),
    .Z(net18297));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19156 (.I(net19155),
    .Z(net19156));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17991 (.I(_15932_[0]),
    .Z(net17991));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17854 (.I(net17852),
    .Z(net17854));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17995 (.I(_15717_[0]),
    .Z(net17995));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17981 (.I(_15959_[0]),
    .Z(net17981));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17831 (.I(_15322_),
    .Z(net17831));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17836 (.I(_15295_),
    .Z(net17836));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17837 (.I(_15295_),
    .Z(net17837));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17843 (.I(_14737_),
    .Z(net17843));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17999 (.I(net17998),
    .Z(net17999));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17863 (.I(_14490_),
    .Z(net17863));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17941 (.I(_11444_),
    .Z(net17941));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17861 (.I(_14502_),
    .Z(net17861));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17842 (.I(_15034_),
    .Z(net17842));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18010 (.I(_06994_),
    .Z(net18010));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17853 (.I(net17852),
    .Z(net17853));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18003 (.I(_15708_[0]),
    .Z(net18003));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17973 (.I(_16019_[0]),
    .Z(net17973));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17908 (.I(net17907),
    .Z(net17908));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17845 (.I(_14667_),
    .Z(net17845));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17847 (.I(_14616_),
    .Z(net17847));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17855 (.I(_14549_),
    .Z(net17855));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17851 (.I(_14579_),
    .Z(net17851));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17859 (.I(_14533_),
    .Z(net17859));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17852 (.I(_14551_),
    .Z(net17852));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17856 (.I(_14544_),
    .Z(net17856));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17921 (.I(_12142_),
    .Z(net17921));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17867 (.I(_14438_),
    .Z(net17867));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17997 (.I(_15712_[0]),
    .Z(net17997));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17860 (.I(_14525_),
    .Z(net17860));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17870 (.I(_13993_),
    .Z(net17870));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17862 (.I(_14490_),
    .Z(net17862));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17885 (.I(net526),
    .Z(net17885));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17868 (.I(_14387_),
    .Z(net17868));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17866 (.I(_14438_),
    .Z(net17866));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17864 (.I(_14463_),
    .Z(net17864));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17873 (.I(_13852_),
    .Z(net17873));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17871 (.I(_13947_),
    .Z(net17871));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17869 (.I(_14201_),
    .Z(net17869));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17879 (.I(_13782_),
    .Z(net17879));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17874 (.I(net603),
    .Z(net17874));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18160 (.I(_01725_),
    .Z(net18160));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17965 (.I(_10597_),
    .Z(net17965));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17883 (.I(_13750_),
    .Z(net17883));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17875 (.I(_13827_),
    .Z(net17875));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17872 (.I(_13861_),
    .Z(net17872));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17877 (.I(net635),
    .Z(net17877));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17876 (.I(_13811_),
    .Z(net17876));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17880 (.I(_13761_),
    .Z(net17880));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17881 (.I(_13755_),
    .Z(net17881));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17884 (.I(_13706_),
    .Z(net17884));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17909 (.I(net17908),
    .Z(net17909));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17958 (.I(_10622_),
    .Z(net17958));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17928 (.I(_11633_),
    .Z(net17928));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17905 (.I(_12997_),
    .Z(net17905));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17949 (.I(_10718_),
    .Z(net17949));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17903 (.I(net17902),
    .Z(net17903));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17925 (.I(net642),
    .Z(net17925));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17918 (.I(_12203_),
    .Z(net17918));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17907 (.I(_12989_),
    .Z(net17907));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17891 (.I(_13095_),
    .Z(net17891));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17967 (.I(net17966),
    .Z(net17967));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17895 (.I(_13075_),
    .Z(net17895));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17893 (.I(_13093_),
    .Z(net17893));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17913 (.I(_12365_),
    .Z(net17913));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17896 (.I(_13060_),
    .Z(net17896));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17898 (.I(_13052_),
    .Z(net17898));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17904 (.I(net17902),
    .Z(net17904));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17959 (.I(_10622_),
    .Z(net17959));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17923 (.I(_12133_),
    .Z(net17923));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17900 (.I(_13033_),
    .Z(net17900));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17910 (.I(_12951_),
    .Z(net17910));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17902 (.I(_13000_),
    .Z(net17902));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17906 (.I(net17905),
    .Z(net17906));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17911 (.I(_12682_),
    .Z(net17911));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17914 (.I(_12316_),
    .Z(net17914));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17912 (.I(_12365_),
    .Z(net17912));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place17924 (.I(_12133_),
    .Z(net17924));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17917 (.I(_12205_),
    .Z(net17917));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17915 (.I(_12308_),
    .Z(net17915));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17962 (.I(_10613_),
    .Z(net17962));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17916 (.I(_12225_),
    .Z(net17916));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17930 (.I(_11588_),
    .Z(net17930));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17945 (.I(_11246_),
    .Z(net17945));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17919 (.I(_12145_),
    .Z(net17919));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17936 (.I(_11490_),
    .Z(net17936));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17922 (.I(net642),
    .Z(net17922));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17926 (.I(_12125_),
    .Z(net17926));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17929 (.I(_11633_),
    .Z(net17929));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17960 (.I(_10618_),
    .Z(net17960));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17979 (.I(_16004_[0]),
    .Z(net17979));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17998 (.I(_15712_[0]),
    .Z(net17998));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17940 (.I(_11444_),
    .Z(net17940));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17931 (.I(_11580_),
    .Z(net17931));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17934 (.I(_11493_),
    .Z(net17934));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17932 (.I(_11543_),
    .Z(net17932));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17937 (.I(_11480_),
    .Z(net17937));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17952 (.I(_10706_),
    .Z(net17952));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17938 (.I(_11467_),
    .Z(net17938));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17933 (.I(_11538_),
    .Z(net17933));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17935 (.I(_11490_),
    .Z(net17935));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17939 (.I(_11454_),
    .Z(net17939));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17942 (.I(_11424_),
    .Z(net17942));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17950 (.I(_10718_),
    .Z(net17950));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17946 (.I(_11244_),
    .Z(net17946));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17947 (.I(_10942_),
    .Z(net17947));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17977 (.I(_16010_[0]),
    .Z(net17977));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17944 (.I(_11292_),
    .Z(net17944));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17971 (.I(_16029_[0]),
    .Z(net17971));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17948 (.I(_10905_),
    .Z(net17948));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17953 (.I(_10692_),
    .Z(net17953));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17951 (.I(_10706_),
    .Z(net17951));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17956 (.I(_10647_),
    .Z(net17956));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17954 (.I(_10672_),
    .Z(net17954));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17955 (.I(_10649_),
    .Z(net17955));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17970 (.I(_10495_),
    .Z(net17970));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17957 (.I(_10626_),
    .Z(net17957));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17961 (.I(_10613_),
    .Z(net17961));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17963 (.I(_10607_),
    .Z(net17963));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17969 (.I(_10495_),
    .Z(net17969));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17964 (.I(_10602_),
    .Z(net17964));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17966 (.I(_10561_),
    .Z(net17966));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17968 (.I(_10495_),
    .Z(net17968));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17990 (.I(_15933_[0]),
    .Z(net17990));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18016 (.I(_06943_),
    .Z(net18016));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17972 (.I(_16026_[0]),
    .Z(net17972));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18009 (.I(_07009_),
    .Z(net18009));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18176 (.I(_01045_),
    .Z(net18176));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17976 (.I(_16010_[0]),
    .Z(net17976));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17974 (.I(_16015_[0]),
    .Z(net17974));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17975 (.I(_16013_[0]),
    .Z(net17975));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17978 (.I(_16008_[0]),
    .Z(net17978));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17982 (.I(_15954_[0]),
    .Z(net17982));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17987 (.I(net17986),
    .Z(net17987));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17980 (.I(_16003_[0]),
    .Z(net17980));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17986 (.I(_15938_[0]),
    .Z(net17986));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17985 (.I(_15941_[0]),
    .Z(net17985));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17983 (.I(_15947_[0]),
    .Z(net17983));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18002 (.I(_15708_[0]),
    .Z(net18002));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17984 (.I(_15943_[0]),
    .Z(net17984));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18189 (.I(_00939_),
    .Z(net18189));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17992 (.I(_15931_[0]),
    .Z(net17992));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17993 (.I(_15728_[0]),
    .Z(net17993));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18007 (.I(_07132_),
    .Z(net18007));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18000 (.I(_15709_[0]),
    .Z(net18000));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17994 (.I(_15721_[0]),
    .Z(net17994));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17996 (.I(_15715_[0]),
    .Z(net17996));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18004 (.I(_15707_[0]),
    .Z(net18004));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18181 (.I(_00973_),
    .Z(net18181));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18005 (.I(_07207_),
    .Z(net18005));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18188 (.I(net18186),
    .Z(net18188));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18006 (.I(_07132_),
    .Z(net18006));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18008 (.I(_07123_),
    .Z(net18008));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18165 (.I(_01193_),
    .Z(net18165));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18162 (.I(_01510_),
    .Z(net18162));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18013 (.I(_06958_),
    .Z(net18013));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18148 (.I(_02406_),
    .Z(net18148));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18066 (.I(_04781_),
    .Z(net18066));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18187 (.I(net18186),
    .Z(net18187));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18011 (.I(_06983_),
    .Z(net18011));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18186 (.I(_00939_),
    .Z(net18186));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18015 (.I(_06944_),
    .Z(net18015));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18041 (.I(_05509_),
    .Z(net18041));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18067 (.I(_04781_),
    .Z(net18067));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18024 (.I(_06351_),
    .Z(net18024));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18023 (.I(_06489_),
    .Z(net18023));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18034 (.I(_06122_),
    .Z(net18034));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18029 (.I(_06209_),
    .Z(net18029));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18020 (.I(_06823_),
    .Z(net18020));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18096 (.I(_04047_),
    .Z(net18096));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18039 (.I(_05528_),
    .Z(net18039));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18025 (.I(_06303_),
    .Z(net18025));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18026 (.I(_06234_),
    .Z(net18026));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18027 (.I(_06216_),
    .Z(net18027));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18033 (.I(_06167_),
    .Z(net18033));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18028 (.I(_06209_),
    .Z(net18028));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18051 (.I(_05393_),
    .Z(net18051));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18032 (.I(_06180_),
    .Z(net18032));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18101 (.I(net18100),
    .Z(net18101));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18038 (.I(_05550_),
    .Z(net18038));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18037 (.I(_05653_),
    .Z(net18037));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18036 (.I(_05812_),
    .Z(net18036));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18042 (.I(_05503_),
    .Z(net18042));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18040 (.I(_05509_),
    .Z(net18040));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18046 (.I(_05431_),
    .Z(net18046));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18132 (.I(net18131),
    .Z(net18132));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18072 (.I(_04754_),
    .Z(net18072));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18047 (.I(_05429_),
    .Z(net18047));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18103 (.I(_04009_),
    .Z(net18103));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18053 (.I(_05338_),
    .Z(net18053));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18056 (.I(_04925_),
    .Z(net18056));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18049 (.I(_05406_),
    .Z(net18049));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18052 (.I(_05373_),
    .Z(net18052));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18050 (.I(_05393_),
    .Z(net18050));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18060 (.I(_04852_),
    .Z(net18060));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18076 (.I(net18075),
    .Z(net18076));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18058 (.I(_04858_),
    .Z(net18058));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18115 (.I(_03938_),
    .Z(net18115));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18063 (.I(_04785_),
    .Z(net18063));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18061 (.I(_04826_),
    .Z(net18061));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18064 (.I(_04781_),
    .Z(net18064));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18071 (.I(_04767_),
    .Z(net18071));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18097 (.I(net18096),
    .Z(net18097));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18074 (.I(_04728_),
    .Z(net18074));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18102 (.I(_04015_),
    .Z(net18102));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18082 (.I(_04626_),
    .Z(net18082));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18078 (.I(_04663_),
    .Z(net18078));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18124 (.I(_03235_),
    .Z(net18124));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18173 (.I(_01073_),
    .Z(net18173));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18084 (.I(_04431_),
    .Z(net18084));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18091 (.I(_04093_),
    .Z(net18091));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place18111 (.I(_03973_),
    .Z(net18111));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18089 (.I(_04115_),
    .Z(net18089));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18087 (.I(_04233_),
    .Z(net18087));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18085 (.I(_04233_),
    .Z(net18085));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18088 (.I(_04117_),
    .Z(net18088));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18090 (.I(_04109_),
    .Z(net18090));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18092 (.I(_04083_),
    .Z(net18092));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18107 (.I(net18106),
    .Z(net18107));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18095 (.I(_04047_),
    .Z(net18095));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18098 (.I(_04042_),
    .Z(net18098));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18099 (.I(_04021_),
    .Z(net18099));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18100 (.I(_04015_),
    .Z(net18100));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18104 (.I(_04004_),
    .Z(net18104));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18105 (.I(_03982_),
    .Z(net18105));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18108 (.I(_03980_),
    .Z(net18108));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18130 (.I(_02717_),
    .Z(net18130));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18109 (.I(net18108),
    .Z(net18109));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18122 (.I(_03254_),
    .Z(net18122));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18113 (.I(net18112),
    .Z(net18113));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place18112 (.I(_03965_),
    .Z(net18112));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18119 (.I(_03286_),
    .Z(net18119));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18114 (.I(_03938_),
    .Z(net18114));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18121 (.I(_03286_),
    .Z(net18121));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18120 (.I(_03286_),
    .Z(net18120));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18125 (.I(_03235_),
    .Z(net18125));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18117 (.I(_03400_),
    .Z(net18117));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18116 (.I(_03405_),
    .Z(net18116));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18127 (.I(_03162_),
    .Z(net18127));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18147 (.I(_02429_),
    .Z(net18147));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18128 (.I(_02742_),
    .Z(net18128));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18159 (.I(_01725_),
    .Z(net18159));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18155 (.I(_01833_),
    .Z(net18155));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18158 (.I(_01725_),
    .Z(net18158));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18152 (.I(_01906_),
    .Z(net18152));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18143 (.I(_02466_),
    .Z(net18143));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18131 (.I(_02643_),
    .Z(net18131));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18133 (.I(_02548_),
    .Z(net18133));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18149 (.I(_02406_),
    .Z(net18149));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18138 (.I(_02508_),
    .Z(net18138));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18134 (.I(_02538_),
    .Z(net18134));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18135 (.I(_02534_),
    .Z(net18135));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18137 (.I(net18136),
    .Z(net18137));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18145 (.I(_02431_),
    .Z(net18145));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18136 (.I(_02522_),
    .Z(net18136));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18141 (.I(_02487_),
    .Z(net18141));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18139 (.I(_02508_),
    .Z(net18139));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18140 (.I(_02490_),
    .Z(net18140));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18142 (.I(_02471_),
    .Z(net18142));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18144 (.I(_02445_),
    .Z(net18144));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18146 (.I(_02431_),
    .Z(net18146));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18169 (.I(_01132_),
    .Z(net18169));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18154 (.I(_01833_),
    .Z(net18154));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18156 (.I(_01770_),
    .Z(net18156));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18150 (.I(_02397_),
    .Z(net18150));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18151 (.I(_02344_),
    .Z(net18151));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18166 (.I(_01186_),
    .Z(net18166));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18153 (.I(_01885_),
    .Z(net18153));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18157 (.I(_01769_),
    .Z(net18157));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18232 (.I(_14489_),
    .Z(net18232));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18161 (.I(_01715_),
    .Z(net18161));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18305 (.I(_12974_),
    .Z(net18305));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18222 (.I(_14565_),
    .Z(net18222));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18185 (.I(_00939_),
    .Z(net18185));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18163 (.I(_01342_),
    .Z(net18163));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18206 (.I(net18205),
    .Z(net18206));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18180 (.I(_00973_),
    .Z(net18180));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18177 (.I(_00995_),
    .Z(net18177));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18167 (.I(_01153_),
    .Z(net18167));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18170 (.I(_01103_),
    .Z(net18170));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18168 (.I(_01136_),
    .Z(net18168));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18183 (.I(_00971_),
    .Z(net18183));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18174 (.I(_01069_),
    .Z(net18174));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18175 (.I(_01055_),
    .Z(net18175));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18182 (.I(_00971_),
    .Z(net18182));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18179 (.I(_00989_),
    .Z(net18179));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18239 (.I(_14435_),
    .Z(net18239));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18184 (.I(_00939_),
    .Z(net18184));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18238 (.I(net18236),
    .Z(net18238));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18221 (.I(_14600_),
    .Z(net18221));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18204 (.I(net406),
    .Z(net18204));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18201 (.I(net400),
    .Z(net18201));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18251 (.I(_14212_),
    .Z(net18251));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18291 (.I(_13034_),
    .Z(net18291));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18234 (.I(_14470_),
    .Z(net18234));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18304 (.I(net18303),
    .Z(net18304));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18200 (.I(_15866_[0]),
    .Z(net18200));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18199 (.I(_15328_),
    .Z(net18199));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18279 (.I(_13113_),
    .Z(net18279));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18282 (.I(_13112_),
    .Z(net18282));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18294 (.I(net18293),
    .Z(net18294));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18289 (.I(_13056_),
    .Z(net18289));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18208 (.I(_14998_),
    .Z(net18208));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18207 (.I(net18205),
    .Z(net18207));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18215 (.I(_14656_),
    .Z(net18215));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18223 (.I(net18222),
    .Z(net18223));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18209 (.I(_14922_),
    .Z(net18209));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18211 (.I(_14744_),
    .Z(net18211));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19155 (.I(_03151_),
    .Z(net19155));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18303 (.I(_12974_),
    .Z(net18303));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18250 (.I(_14386_),
    .Z(net18250));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18228 (.I(_14534_),
    .Z(net18228));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18216 (.I(_14649_),
    .Z(net18216));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18210 (.I(_14859_),
    .Z(net18210));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18236 (.I(_14435_),
    .Z(net18236));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18212 (.I(_14707_),
    .Z(net18212));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18213 (.I(_14695_),
    .Z(net18213));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18217 (.I(_14643_),
    .Z(net18217));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18214 (.I(_14658_),
    .Z(net18214));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18224 (.I(_14563_),
    .Z(net18224));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18218 (.I(_14624_),
    .Z(net18218));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18225 (.I(_14562_),
    .Z(net18225));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18219 (.I(_14610_),
    .Z(net18219));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18220 (.I(_14600_),
    .Z(net18220));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18226 (.I(_14543_),
    .Z(net18226));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18227 (.I(_14535_),
    .Z(net18227));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18235 (.I(_14462_),
    .Z(net18235));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18233 (.I(_14472_),
    .Z(net18233));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18231 (.I(_14520_),
    .Z(net18231));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18229 (.I(_14531_),
    .Z(net18229));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19110 (.I(net19097),
    .Z(net19110));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19109 (.I(net19097),
    .Z(net19109));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18365 (.I(_16149_[0]),
    .Z(net18365));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18283 (.I(_13100_),
    .Z(net18283));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18368 (.I(_16140_[0]),
    .Z(net18368));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18272 (.I(_13674_),
    .Z(net18272));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18355 (.I(_16185_[0]),
    .Z(net18355));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18352 (.I(_10447_),
    .Z(net18352));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18540 (.I(net18532),
    .Z(net18540));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18333 (.I(_11361_),
    .Z(net18333));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18329 (.I(_11400_),
    .Z(net18329));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place18318 (.I(net485),
    .Z(net18318));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18321 (.I(_11622_),
    .Z(net18321));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18320 (.I(net486),
    .Z(net18320));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18267 (.I(_13801_),
    .Z(net18267));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18275 (.I(_13365_),
    .Z(net18275));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18265 (.I(_13825_),
    .Z(net18265));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18270 (.I(_13776_),
    .Z(net18270));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18255 (.I(_13903_),
    .Z(net18255));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18363 (.I(_16160_[0]),
    .Z(net18363));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18276 (.I(_13211_),
    .Z(net18276));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18257 (.I(_13870_),
    .Z(net18257));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18261 (.I(net18260),
    .Z(net18261));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18268 (.I(_13801_),
    .Z(net18268));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18260 (.I(_13836_),
    .Z(net18260));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18274 (.I(_13392_),
    .Z(net18274));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18264 (.I(_13826_),
    .Z(net18264));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18266 (.I(_13803_),
    .Z(net18266));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18269 (.I(_13781_),
    .Z(net18269));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18300 (.I(_12974_),
    .Z(net18300));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18301 (.I(_12974_),
    .Z(net18301));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18271 (.I(_13716_),
    .Z(net18271));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18280 (.I(_13113_),
    .Z(net18280));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18273 (.I(_13672_),
    .Z(net18273));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18277 (.I(_13191_),
    .Z(net18277));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18299 (.I(net18298),
    .Z(net18299));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18287 (.I(_13077_),
    .Z(net18287));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18281 (.I(_13112_),
    .Z(net18281));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18284 (.I(_13092_),
    .Z(net18284));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18285 (.I(_13085_),
    .Z(net18285));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18288 (.I(_13056_),
    .Z(net18288));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18286 (.I(_13081_),
    .Z(net18286));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18290 (.I(_13050_),
    .Z(net18290));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18293 (.I(_13032_),
    .Z(net18293));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place18316 (.I(net18315),
    .Z(net18316));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18295 (.I(_13020_),
    .Z(net18295));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18296 (.I(_12996_),
    .Z(net18296));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18302 (.I(_12974_),
    .Z(net18302));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18449 (.I(_06310_),
    .Z(net18449));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18455 (.I(_06199_),
    .Z(net18455));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18454 (.I(_06218_),
    .Z(net18454));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18444 (.I(_06878_),
    .Z(net18444));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18312 (.I(_12915_),
    .Z(net18312));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18585 (.I(net18584),
    .Z(net18585));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18534 (.I(net18532),
    .Z(net18534));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18526 (.I(net18525),
    .Z(net18526));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18335 (.I(_11361_),
    .Z(net18335));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18596 (.I(net692),
    .Z(net18596));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18358 (.I(_16176_[0]),
    .Z(net18358));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18317 (.I(_12124_),
    .Z(net18317));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18343 (.I(_10646_),
    .Z(net18343));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18344 (.I(_10625_),
    .Z(net18344));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18346 (.I(_10596_),
    .Z(net18346));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18410 (.I(_15805_[0]),
    .Z(net18410));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18330 (.I(_11400_),
    .Z(net18330));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 place18319 (.I(net18318),
    .Z(net18319));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18323 (.I(_11537_),
    .Z(net18323));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18322 (.I(_11559_),
    .Z(net18322));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18324 (.I(_11453_),
    .Z(net18324));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18327 (.I(_11411_),
    .Z(net18327));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18326 (.I(_11416_),
    .Z(net18326));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18328 (.I(_11400_),
    .Z(net18328));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18334 (.I(_11361_),
    .Z(net18334));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18325 (.I(_11430_),
    .Z(net18325));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18349 (.I(_10536_),
    .Z(net18349));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18424 (.I(net18423),
    .Z(net18424));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18338 (.I(_11359_),
    .Z(net18338));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18350 (.I(_10536_),
    .Z(net18350));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18331 (.I(_11393_),
    .Z(net18331));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18431 (.I(_06993_),
    .Z(net18431));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18332 (.I(_11366_),
    .Z(net18332));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18337 (.I(_11359_),
    .Z(net18337));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18339 (.I(_11357_),
    .Z(net18339));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18336 (.I(_11359_),
    .Z(net18336));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18340 (.I(_11323_),
    .Z(net18340));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18345 (.I(_10621_),
    .Z(net18345));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18341 (.I(_11103_),
    .Z(net18341));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18342 (.I(_10761_),
    .Z(net18342));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18404 (.I(net18403),
    .Z(net18404));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18505 (.I(_04671_),
    .Z(net18505));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18595 (.I(net18586),
    .Z(net18595));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18348 (.I(_10565_),
    .Z(net18348));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18347 (.I(_10575_),
    .Z(net18347));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18786 (.I(_14414_),
    .Z(net18786));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18351 (.I(_10498_),
    .Z(net18351));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18353 (.I(_16197_[0]),
    .Z(net18353));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18594 (.I(net18586),
    .Z(net18594));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18544 (.I(net18543),
    .Z(net18544));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18380 (.I(_16049_[0]),
    .Z(net18380));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18376 (.I(_16108_[0]),
    .Z(net18376));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18357 (.I(_16176_[0]),
    .Z(net18357));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18369 (.I(_16139_[0]),
    .Z(net18369));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18354 (.I(_16192_[0]),
    .Z(net18354));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18356 (.I(_16181_[0]),
    .Z(net18356));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18359 (.I(_16173_[0]),
    .Z(net18359));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18374 (.I(_16109_[0]),
    .Z(net18374));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18361 (.I(_16171_[0]),
    .Z(net18361));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18360 (.I(_16172_[0]),
    .Z(net18360));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18362 (.I(_16165_[0]),
    .Z(net18362));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18389 (.I(_15969_[0]),
    .Z(net18389));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18364 (.I(_16151_[0]),
    .Z(net18364));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18366 (.I(_16144_[0]),
    .Z(net18366));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18367 (.I(_16141_[0]),
    .Z(net18367));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18548 (.I(net18532),
    .Z(net18548));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18373 (.I(net18372),
    .Z(net18373));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18370 (.I(_16133_[0]),
    .Z(net18370));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18371 (.I(_16121_[0]),
    .Z(net18371));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18372 (.I(_16112_[0]),
    .Z(net18372));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18375 (.I(net18374),
    .Z(net18375));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18377 (.I(_16107_[0]),
    .Z(net18377));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18383 (.I(_16040_[0]),
    .Z(net18383));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18379 (.I(_16051_[0]),
    .Z(net18379));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18465 (.I(_06051_),
    .Z(net18465));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18546 (.I(net18543),
    .Z(net18546));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18501 (.I(_04706_),
    .Z(net18501));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18381 (.I(_16046_[0]),
    .Z(net18381));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18547 (.I(net18543),
    .Z(net18547));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18382 (.I(_16041_[0]),
    .Z(net18382));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18384 (.I(_16039_[0]),
    .Z(net18384));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18472 (.I(_05440_),
    .Z(net18472));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18385 (.I(_15995_[0]),
    .Z(net18385));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18545 (.I(net18543),
    .Z(net18545));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18386 (.I(_15990_[0]),
    .Z(net18386));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18387 (.I(_15974_[0]),
    .Z(net18387));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18436 (.I(net520),
    .Z(net18436));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18433 (.I(_06975_),
    .Z(net18433));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18538 (.I(net18532),
    .Z(net18538));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18393 (.I(_15909_[0]),
    .Z(net18393));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18390 (.I(_15968_[0]),
    .Z(net18390));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18396 (.I(_15900_[0]),
    .Z(net18396));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place18397 (.I(_15900_[0]),
    .Z(net18397));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18399 (.I(_15849_[0]),
    .Z(net18399));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18394 (.I(_15904_[0]),
    .Z(net18394));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18395 (.I(_15901_[0]),
    .Z(net18395));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18403 (.I(_15836_[0]),
    .Z(net18403));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18400 (.I(_15845_[0]),
    .Z(net18400));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18430 (.I(_06993_),
    .Z(net18430));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18401 (.I(_15840_[0]),
    .Z(net18401));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18408 (.I(_15808_[0]),
    .Z(net18408));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18402 (.I(_15837_[0]),
    .Z(net18402));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18405 (.I(_15835_[0]),
    .Z(net18405));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18409 (.I(net18408),
    .Z(net18409));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18406 (.I(_15817_[0]),
    .Z(net18406));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18407 (.I(_15808_[0]),
    .Z(net18407));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18411 (.I(_15804_[0]),
    .Z(net18411));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18427 (.I(_07035_),
    .Z(net18427));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18413 (.I(_15785_[0]),
    .Z(net18413));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18417 (.I(_15772_[0]),
    .Z(net18417));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18412 (.I(_15792_[0]),
    .Z(net18412));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18414 (.I(_15781_[0]),
    .Z(net18414));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18415 (.I(_15776_[0]),
    .Z(net18415));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18421 (.I(_15687_[0]),
    .Z(net18421));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18416 (.I(_15773_[0]),
    .Z(net18416));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18418 (.I(_15771_[0]),
    .Z(net18418));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18422 (.I(_15685_[0]),
    .Z(net18422));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18419 (.I(_15696_[0]),
    .Z(net18419));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18420 (.I(_15689_[0]),
    .Z(net18420));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18539 (.I(net18538),
    .Z(net18539));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18543 (.I(net18532),
    .Z(net18543));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18541 (.I(net18532),
    .Z(net18541));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18439 (.I(_06929_),
    .Z(net18439));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18432 (.I(_06980_),
    .Z(net18432));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18426 (.I(_07048_),
    .Z(net18426));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18428 (.I(_07034_),
    .Z(net18428));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18429 (.I(_07000_),
    .Z(net18429));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18437 (.I(_06931_),
    .Z(net18437));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18434 (.I(_06965_),
    .Z(net18434));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18435 (.I(_06931_),
    .Z(net18435));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18447 (.I(_06641_),
    .Z(net18447));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18446 (.I(net476),
    .Z(net18446));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18442 (.I(_06898_),
    .Z(net18442));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18445 (.I(_06786_),
    .Z(net18445));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18441 (.I(_06898_),
    .Z(net18441));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18452 (.I(_06249_),
    .Z(net18452));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18537 (.I(net18532),
    .Z(net18537));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18443 (.I(_06878_),
    .Z(net18443));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18450 (.I(net18449),
    .Z(net18450));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18448 (.I(_06310_),
    .Z(net18448));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18479 (.I(_05392_),
    .Z(net18479));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18469 (.I(_05466_),
    .Z(net18469));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18510 (.I(_04593_),
    .Z(net18510));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18451 (.I(_06262_),
    .Z(net18451));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18453 (.I(_06218_),
    .Z(net18453));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place18502 (.I(_04700_),
    .Z(net18502));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18467 (.I(_05529_),
    .Z(net18467));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18458 (.I(_06158_),
    .Z(net18458));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18457 (.I(_06161_),
    .Z(net18457));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18503 (.I(_04700_),
    .Z(net18503));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18464 (.I(_06051_),
    .Z(net18464));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18462 (.I(_06120_),
    .Z(net18462));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18459 (.I(_06154_),
    .Z(net18459));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18468 (.I(_05529_),
    .Z(net18468));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18460 (.I(_06126_),
    .Z(net18460));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18461 (.I(_06120_),
    .Z(net18461));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18463 (.I(_06061_),
    .Z(net18463));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18593 (.I(net18586),
    .Z(net18593));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18466 (.I(_05646_),
    .Z(net18466));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18482 (.I(_05391_),
    .Z(net18482));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18727 (.I(_15150_),
    .Z(net18727));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18722 (.I(net18708),
    .Z(net18722));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18488 (.I(_04896_),
    .Z(net18488));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18476 (.I(_05394_),
    .Z(net18476));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18500 (.I(_04709_),
    .Z(net18500));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18592 (.I(net692),
    .Z(net18592));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18474 (.I(_05403_),
    .Z(net18474));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18486 (.I(net18485),
    .Z(net18486));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18475 (.I(_05394_),
    .Z(net18475));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18478 (.I(_05392_),
    .Z(net18478));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18481 (.I(_05391_),
    .Z(net18481));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18483 (.I(_05363_),
    .Z(net18483));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18484 (.I(_05345_),
    .Z(net18484));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18487 (.I(_04909_),
    .Z(net18487));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18490 (.I(_04857_),
    .Z(net18490));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18485 (.I(_05307_),
    .Z(net18485));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18597 (.I(net18596),
    .Z(net18597));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18491 (.I(_04833_),
    .Z(net18491));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18493 (.I(_04753_),
    .Z(net18493));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18558 (.I(_03345_),
    .Z(net18558));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18492 (.I(_04796_),
    .Z(net18492));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18489 (.I(_04865_),
    .Z(net18489));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18499 (.I(_04714_),
    .Z(net18499));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18496 (.I(net18495),
    .Z(net18496));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18495 (.I(_04724_),
    .Z(net18495));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18494 (.I(_04742_),
    .Z(net18494));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18498 (.I(_04716_),
    .Z(net18498));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18509 (.I(_04597_),
    .Z(net18509));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18497 (.I(_04717_),
    .Z(net18497));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18504 (.I(_04696_),
    .Z(net18504));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18506 (.I(_04666_),
    .Z(net18506));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18591 (.I(net18586),
    .Z(net18591));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18523 (.I(net18522),
    .Z(net18523));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18507 (.I(_04656_),
    .Z(net18507));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18508 (.I(_04631_),
    .Z(net18508));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18512 (.I(_04139_),
    .Z(net18512));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18517 (.I(_03985_),
    .Z(net18517));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18511 (.I(_04150_),
    .Z(net18511));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18590 (.I(net691),
    .Z(net18590));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18514 (.I(_04049_),
    .Z(net18514));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18566 (.I(net18565),
    .Z(net18566));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18524 (.I(net18522),
    .Z(net18524));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18562 (.I(_03227_),
    .Z(net18562));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18522 (.I(_03967_),
    .Z(net18522));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18527 (.I(net18525),
    .Z(net18527));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18531 (.I(net18530),
    .Z(net18531));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18528 (.I(_03926_),
    .Z(net18528));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18601 (.I(net691),
    .Z(net18601));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18530 (.I(_03896_),
    .Z(net18530));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18529 (.I(_03896_),
    .Z(net18529));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18609 (.I(net18605),
    .Z(net18609));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18567 (.I(net527),
    .Z(net18567));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18560 (.I(_03243_),
    .Z(net18560));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18602 (.I(net691),
    .Z(net18602));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18600 (.I(net692),
    .Z(net18600));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18559 (.I(_03243_),
    .Z(net18559));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18608 (.I(net18605),
    .Z(net18608));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18607 (.I(net18606),
    .Z(net18607));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18646 (.I(_01623_),
    .Z(net18646));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18721 (.I(net18720),
    .Z(net18721));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18720 (.I(net18708),
    .Z(net18720));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18719 (.I(net18708),
    .Z(net18719));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18631 (.I(net18623),
    .Z(net18631));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18630 (.I(net18623),
    .Z(net18630));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18629 (.I(net18623),
    .Z(net18629));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18628 (.I(net18623),
    .Z(net18628));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18570 (.I(_02566_),
    .Z(net18570));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18589 (.I(net692),
    .Z(net18589));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18561 (.I(_03227_),
    .Z(net18561));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18565 (.I(_16002_[0]),
    .Z(net18565));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18574 (.I(_02480_),
    .Z(net18574));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18636 (.I(_01646_),
    .Z(net18636));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18627 (.I(net18623),
    .Z(net18627));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18637 (.I(net18636),
    .Z(net18637));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18603 (.I(_02388_),
    .Z(net18603));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18577 (.I(_02462_),
    .Z(net18577));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18584 (.I(_02396_),
    .Z(net18584));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18564 (.I(_16002_[0]),
    .Z(net18564));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18563 (.I(_03197_),
    .Z(net18563));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18616 (.I(_01774_),
    .Z(net18616));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18580 (.I(_02401_),
    .Z(net18580));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18626 (.I(net18623),
    .Z(net18626));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18606 (.I(net18605),
    .Z(net18606));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18604 (.I(_02388_),
    .Z(net18604));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18582 (.I(_02401_),
    .Z(net18582));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18568 (.I(_02624_),
    .Z(net18568));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18569 (.I(_02566_),
    .Z(net18569));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18576 (.I(_02462_),
    .Z(net18576));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18573 (.I(_02480_),
    .Z(net18573));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18571 (.I(_02506_),
    .Z(net18571));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18575 (.I(_02463_),
    .Z(net18575));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18572 (.I(_02480_),
    .Z(net18572));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18581 (.I(_02401_),
    .Z(net18581));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18578 (.I(_02443_),
    .Z(net18578));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18579 (.I(_02401_),
    .Z(net18579));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18587 (.I(net18586),
    .Z(net18587));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18634 (.I(_01670_),
    .Z(net18634));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18583 (.I(_02396_),
    .Z(net18583));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 place18586 (.I(_02391_),
    .Z(net18586));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18788 (.I(net18786),
    .Z(net18788));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18625 (.I(net18623),
    .Z(net18625));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18624 (.I(net18623),
    .Z(net18624));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18726 (.I(_15150_),
    .Z(net18726));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18632 (.I(net18623),
    .Z(net18632));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18621 (.I(_01691_),
    .Z(net18621));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18698 (.I(net18684),
    .Z(net18698));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18697 (.I(net18684),
    .Z(net18697));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18680 (.I(net18676),
    .Z(net18680));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18679 (.I(net18676),
    .Z(net18679));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18678 (.I(net18676),
    .Z(net18678));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18645 (.I(net18636),
    .Z(net18645));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18644 (.I(net18636),
    .Z(net18644));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18718 (.I(net18708),
    .Z(net18718));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18643 (.I(net18636),
    .Z(net18643));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18620 (.I(_01691_),
    .Z(net18620));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18677 (.I(net18676),
    .Z(net18677));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20435 (.I(net20433),
    .Z(net20435));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18244 (.I(net18240),
    .Z(net18244));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place18623 (.I(_01670_),
    .Z(net18623));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18962 (.I(net18961),
    .Z(net18962));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18902 (.I(net18901),
    .Z(net18902));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18901 (.I(_12053_),
    .Z(net18901));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18694 (.I(net18684),
    .Z(net18694));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18693 (.I(net18691),
    .Z(net18693));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18676 (.I(_00946_),
    .Z(net18676));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18692 (.I(net18691),
    .Z(net18692));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18691 (.I(net18684),
    .Z(net18691));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18690 (.I(net18684),
    .Z(net18690));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18689 (.I(net18688),
    .Z(net18689));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18675 (.I(net18670),
    .Z(net18675));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18701 (.I(net18684),
    .Z(net18701));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place18688 (.I(net18684),
    .Z(net18688));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18717 (.I(net18708),
    .Z(net18717));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18687 (.I(net18684),
    .Z(net18687));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18686 (.I(net18684),
    .Z(net18686));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18974 (.I(net18973),
    .Z(net18974));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18652 (.I(net389),
    .Z(net18652));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer78 (.I(_01730_),
    .Z(net465));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18716 (.I(net18708),
    .Z(net18716));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18973 (.I(net18971),
    .Z(net18973));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18656 (.I(_01110_),
    .Z(net18656));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18715 (.I(net18708),
    .Z(net18715));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18972 (.I(net18971),
    .Z(net18972));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18746 (.I(_14493_),
    .Z(net18746));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18742 (.I(_14530_),
    .Z(net18742));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18714 (.I(net18708),
    .Z(net18714));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18243 (.I(net18242),
    .Z(net18243));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18751 (.I(net18750),
    .Z(net18751));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18785 (.I(_14414_),
    .Z(net18785));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18663 (.I(net18662),
    .Z(net18663));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18655 (.I(_01110_),
    .Z(net18655));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18668 (.I(_01024_),
    .Z(net18668));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18671 (.I(net18670),
    .Z(net18671));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19029 (.I(net19022),
    .Z(net19029));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19027 (.I(net19022),
    .Z(net19027));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18753 (.I(net18750),
    .Z(net18753));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18762 (.I(net18761),
    .Z(net18762));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18725 (.I(net18724),
    .Z(net18725));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18763 (.I(net18750),
    .Z(net18763));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18672 (.I(net18670),
    .Z(net18672));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18737 (.I(net18734),
    .Z(net18737));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18723 (.I(net18708),
    .Z(net18723));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19120 (.I(_03946_),
    .Z(net19120));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18993 (.I(net18992),
    .Z(net18993));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18683 (.I(net18682),
    .Z(net18683));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18665 (.I(_01057_),
    .Z(net18665));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18736 (.I(net18734),
    .Z(net18736));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18734 (.I(_15150_),
    .Z(net18734));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18657 (.I(_01106_),
    .Z(net18657));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18654 (.I(_01120_),
    .Z(net18654));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18733 (.I(net18731),
    .Z(net18733));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18730 (.I(net18729),
    .Z(net18730));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18658 (.I(_01104_),
    .Z(net18658));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18662 (.I(_01072_),
    .Z(net18662));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18670 (.I(_00946_),
    .Z(net18670));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18667 (.I(_01024_),
    .Z(net18667));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18659 (.I(_01099_),
    .Z(net18659));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18660 (.I(_01080_),
    .Z(net18660));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18669 (.I(_00988_),
    .Z(net18669));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18661 (.I(_01072_),
    .Z(net18661));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18664 (.I(_01057_),
    .Z(net18664));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18666 (.I(_01024_),
    .Z(net18666));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18713 (.I(net18708),
    .Z(net18713));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18682 (.I(_00943_),
    .Z(net18682));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18732 (.I(net18731),
    .Z(net18732));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18696 (.I(net18694),
    .Z(net18696));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18731 (.I(_15150_),
    .Z(net18731));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18705 (.I(_15245_),
    .Z(net18705));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18712 (.I(net18708),
    .Z(net18712));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18704 (.I(_15245_),
    .Z(net18704));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18710 (.I(net18709),
    .Z(net18710));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18761 (.I(net18750),
    .Z(net18761));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18754 (.I(net18750),
    .Z(net18754));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18706 (.I(_15219_),
    .Z(net18706));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18744 (.I(_14519_),
    .Z(net18744));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18724 (.I(_15150_),
    .Z(net18724));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18760 (.I(net18750),
    .Z(net18760));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18758 (.I(net18750),
    .Z(net18758));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18757 (.I(net18754),
    .Z(net18757));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18756 (.I(net18754),
    .Z(net18756));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18755 (.I(net18754),
    .Z(net18755));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18759 (.I(net18750),
    .Z(net18759));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18740 (.I(_14638_),
    .Z(net18740));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18784 (.I(net18783),
    .Z(net18784));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18749 (.I(_14446_),
    .Z(net18749));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18783 (.I(_14414_),
    .Z(net18783));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18782 (.I(net18781),
    .Z(net18782));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18764 (.I(_14434_),
    .Z(net18764));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18739 (.I(_14638_),
    .Z(net18739));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18709 (.I(net18708),
    .Z(net18709));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18707 (.I(_15201_),
    .Z(net18707));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18770 (.I(net18764),
    .Z(net18770));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18769 (.I(net18768),
    .Z(net18769));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18768 (.I(net18764),
    .Z(net18768));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18752 (.I(net18750),
    .Z(net18752));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18992 (.I(_06782_),
    .Z(net18992));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18988 (.I(_06782_),
    .Z(net18988));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18738 (.I(_14648_),
    .Z(net18738));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18708 (.I(_15196_),
    .Z(net18708));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18735 (.I(net18734),
    .Z(net18735));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18767 (.I(net18764),
    .Z(net18767));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18766 (.I(net18764),
    .Z(net18766));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18987 (.I(net18985),
    .Z(net18987));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18741 (.I(_14582_),
    .Z(net18741));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18825 (.I(net18813),
    .Z(net18825));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18796 (.I(_13793_),
    .Z(net18796));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18780 (.I(net18771),
    .Z(net18780));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18781 (.I(_14414_),
    .Z(net18781));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18779 (.I(net18771),
    .Z(net18779));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18778 (.I(net18771),
    .Z(net18778));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18777 (.I(net18771),
    .Z(net18777));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18776 (.I(net18771),
    .Z(net18776));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18775 (.I(net18771),
    .Z(net18775));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18774 (.I(net18771),
    .Z(net18774));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18773 (.I(net18771),
    .Z(net18773));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18792 (.I(_13922_),
    .Z(net18792));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18748 (.I(_14446_),
    .Z(net18748));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18772 (.I(net18771),
    .Z(net18772));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18824 (.I(net18813),
    .Z(net18824));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18810 (.I(net18806),
    .Z(net18810));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18765 (.I(net18764),
    .Z(net18765));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18801 (.I(_13753_),
    .Z(net18801));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18797 (.I(_13793_),
    .Z(net18797));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18823 (.I(net18813),
    .Z(net18823));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18986 (.I(net18985),
    .Z(net18986));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18822 (.I(net18813),
    .Z(net18822));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18985 (.I(_06782_),
    .Z(net18985));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18771 (.I(_14414_),
    .Z(net18771));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18743 (.I(_14519_),
    .Z(net18743));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18745 (.I(_14493_),
    .Z(net18745));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18747 (.I(_14493_),
    .Z(net18747));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18750 (.I(_14441_),
    .Z(net18750));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18991 (.I(_06782_),
    .Z(net18991));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18787 (.I(net18786),
    .Z(net18787));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18990 (.I(net18988),
    .Z(net18990));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18791 (.I(_13922_),
    .Z(net18791));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18989 (.I(net18988),
    .Z(net18989));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18952 (.I(_16080_[0]),
    .Z(net18952));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18950 (.I(_16096_[0]),
    .Z(net18950));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18911 (.I(_11363_),
    .Z(net18911));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18819 (.I(net18818),
    .Z(net18819));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18949 (.I(_09544_),
    .Z(net18949));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18964 (.I(net18961),
    .Z(net18964));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19051 (.I(net19038),
    .Z(net19051));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18818 (.I(net18813),
    .Z(net18818));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18904 (.I(_11528_),
    .Z(net18904));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19090 (.I(net19082),
    .Z(net19090));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18813 (.I(_13701_),
    .Z(net18813));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18817 (.I(net18813),
    .Z(net18817));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18816 (.I(net18813),
    .Z(net18816));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18794 (.I(_13796_),
    .Z(net18794));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18815 (.I(net18813),
    .Z(net18815));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18814 (.I(net18813),
    .Z(net18814));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18800 (.I(_13753_),
    .Z(net18800));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18798 (.I(_13775_),
    .Z(net18798));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18793 (.I(_13843_),
    .Z(net18793));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19054 (.I(net19038),
    .Z(net19054));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18866 (.I(net18854),
    .Z(net18866));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18865 (.I(net18854),
    .Z(net18865));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18864 (.I(net18854),
    .Z(net18864));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18820 (.I(net18813),
    .Z(net18820));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18802 (.I(_13721_),
    .Z(net18802));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18795 (.I(_13793_),
    .Z(net18795));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18809 (.I(net18806),
    .Z(net18809));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18799 (.I(_13753_),
    .Z(net18799));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19053 (.I(net19052),
    .Z(net19053));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18977 (.I(net18971),
    .Z(net18977));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18867 (.I(_12918_),
    .Z(net18867));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18976 (.I(net18971),
    .Z(net18976));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18804 (.I(_13721_),
    .Z(net18804));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18975 (.I(net18971),
    .Z(net18975));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18803 (.I(_13721_),
    .Z(net18803));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18899 (.I(net18894),
    .Z(net18899));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18898 (.I(net18894),
    .Z(net18898));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18971 (.I(_06827_),
    .Z(net18971));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18897 (.I(net18894),
    .Z(net18897));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18863 (.I(net18854),
    .Z(net18863));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18896 (.I(net18894),
    .Z(net18896));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18808 (.I(net18806),
    .Z(net18808));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18807 (.I(net18806),
    .Z(net18807));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18806 (.I(_13709_),
    .Z(net18806));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18805 (.I(_13719_),
    .Z(net18805));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18862 (.I(net18854),
    .Z(net18862));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18861 (.I(net18854),
    .Z(net18861));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19092 (.I(net19082),
    .Z(net19092));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18848 (.I(_12994_),
    .Z(net18848));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18860 (.I(net18854),
    .Z(net18860));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18834 (.I(_13139_),
    .Z(net18834));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18833 (.I(_13174_),
    .Z(net18833));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18894 (.I(_12121_),
    .Z(net18894));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18893 (.I(net18887),
    .Z(net18893));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18892 (.I(net18887),
    .Z(net18892));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18891 (.I(net18887),
    .Z(net18891));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18878 (.I(net18875),
    .Z(net18878));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18890 (.I(net18887),
    .Z(net18890));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18884 (.I(_12201_),
    .Z(net18884));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18871 (.I(_12863_),
    .Z(net18871));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18870 (.I(_12863_),
    .Z(net18870));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18881 (.I(net18875),
    .Z(net18881));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18853 (.I(_12946_),
    .Z(net18853));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18838 (.I(_13091_),
    .Z(net18838));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18845 (.I(_13024_),
    .Z(net18845));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18882 (.I(_12208_),
    .Z(net18882));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18248 (.I(_14435_),
    .Z(net18248));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18970 (.I(_06827_),
    .Z(net18970));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18969 (.I(net18967),
    .Z(net18969));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18839 (.I(_13058_),
    .Z(net18839));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18836 (.I(_13129_),
    .Z(net18836));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18918 (.I(net18916),
    .Z(net18918));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18917 (.I(net18916),
    .Z(net18917));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18851 (.I(_12976_),
    .Z(net18851));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18847 (.I(_12994_),
    .Z(net18847));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18880 (.I(net18875),
    .Z(net18880));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18837 (.I(_13091_),
    .Z(net18837));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18888 (.I(net18887),
    .Z(net18888));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18883 (.I(_12201_),
    .Z(net18883));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18841 (.I(_13030_),
    .Z(net18841));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18842 (.I(_13025_),
    .Z(net18842));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18843 (.I(_13025_),
    .Z(net18843));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18840 (.I(_13030_),
    .Z(net18840));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18879 (.I(net18875),
    .Z(net18879));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18844 (.I(_13024_),
    .Z(net18844));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18846 (.I(_13022_),
    .Z(net18846));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18875 (.I(_12212_),
    .Z(net18875));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18877 (.I(net18875),
    .Z(net18877));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18849 (.I(_12981_),
    .Z(net18849));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18869 (.I(_12918_),
    .Z(net18869));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18850 (.I(_12976_),
    .Z(net18850));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18852 (.I(_12946_),
    .Z(net18852));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18868 (.I(_12918_),
    .Z(net18868));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18854 (.I(_12943_),
    .Z(net18854));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19091 (.I(net19082),
    .Z(net19091));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18900 (.I(_12053_),
    .Z(net18900));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18872 (.I(_12478_),
    .Z(net18872));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18953 (.I(_16077_[0]),
    .Z(net18953));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19184 (.I(_01777_),
    .Z(net19184));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19107 (.I(net19097),
    .Z(net19107));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18945 (.I(_09840_),
    .Z(net18945));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18932 (.I(_10699_),
    .Z(net18932));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18906 (.I(_11429_),
    .Z(net18906));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18944 (.I(_09851_),
    .Z(net18944));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18247 (.I(_14435_),
    .Z(net18247));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18246 (.I(_14435_),
    .Z(net18246));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18978 (.I(_06820_),
    .Z(net18978));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19037 (.I(net19035),
    .Z(net19037));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18876 (.I(net18875),
    .Z(net18876));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18873 (.I(_12391_),
    .Z(net18873));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18889 (.I(net18887),
    .Z(net18889));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18886 (.I(_12174_),
    .Z(net18886));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19036 (.I(net19035),
    .Z(net19036));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18885 (.I(_12174_),
    .Z(net18885));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18874 (.I(_12224_),
    .Z(net18874));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18895 (.I(net18894),
    .Z(net18895));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18903 (.I(net18902),
    .Z(net18903));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19035 (.I(net19022),
    .Z(net19035));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18943 (.I(_09934_),
    .Z(net18943));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19034 (.I(net19022),
    .Z(net19034));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19033 (.I(net19022),
    .Z(net19033));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18934 (.I(_10688_),
    .Z(net18934));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18916 (.I(net18915),
    .Z(net18916));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19032 (.I(net19022),
    .Z(net19032));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place18887 (.I(_12121_),
    .Z(net18887));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18930 (.I(_10703_),
    .Z(net18930));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18910 (.I(_11363_),
    .Z(net18910));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18905 (.I(_11429_),
    .Z(net18905));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19031 (.I(net19030),
    .Z(net19031));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18968 (.I(net18967),
    .Z(net18968));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18967 (.I(_06827_),
    .Z(net18967));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19030 (.I(net19022),
    .Z(net19030));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18914 (.I(_11356_),
    .Z(net18914));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19088 (.I(net19082),
    .Z(net19088));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18913 (.I(_11356_),
    .Z(net18913));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18907 (.I(_11408_),
    .Z(net18907));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19089 (.I(net19082),
    .Z(net19089));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18998 (.I(_06726_),
    .Z(net18998));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18919 (.I(_11186_),
    .Z(net18919));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19001 (.I(net19000),
    .Z(net19001));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18965 (.I(net18961),
    .Z(net18965));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19026 (.I(net19022),
    .Z(net19026));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19173 (.I(_15965_[0]),
    .Z(net19173));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18908 (.I(_11392_),
    .Z(net18908));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18909 (.I(_11363_),
    .Z(net18909));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place18915 (.I(_15706_[0]),
    .Z(net18915));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18912 (.I(_11356_),
    .Z(net18912));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18984 (.I(net18978),
    .Z(net18984));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18920 (.I(net18919),
    .Z(net18920));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18983 (.I(net18978),
    .Z(net18983));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18928 (.I(_10729_),
    .Z(net18928));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18923 (.I(_11088_),
    .Z(net18923));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18966 (.I(_06827_),
    .Z(net18966));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18927 (.I(_10746_),
    .Z(net18927));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18924 (.I(_10867_),
    .Z(net18924));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18982 (.I(net18978),
    .Z(net18982));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18925 (.I(_10771_),
    .Z(net18925));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18935 (.I(_10677_),
    .Z(net18935));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18931 (.I(_10699_),
    .Z(net18931));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18929 (.I(_10703_),
    .Z(net18929));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18926 (.I(_10746_),
    .Z(net18926));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18979 (.I(net18978),
    .Z(net18979));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18933 (.I(_10688_),
    .Z(net18933));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18995 (.I(_06763_),
    .Z(net18995));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19172 (.I(net19171),
    .Z(net19172));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19025 (.I(net19022),
    .Z(net19025));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19024 (.I(net19022),
    .Z(net19024));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18947 (.I(_09840_),
    .Z(net18947));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19528 (.I(net19515),
    .Z(net19528));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18940 (.I(_10595_),
    .Z(net18940));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18936 (.I(_10666_),
    .Z(net18936));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19087 (.I(net19082),
    .Z(net19087));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18960 (.I(_06851_),
    .Z(net18960));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18937 (.I(_10645_),
    .Z(net18937));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18938 (.I(_10615_),
    .Z(net18938));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19086 (.I(net19082),
    .Z(net19086));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18939 (.I(_10595_),
    .Z(net18939));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18941 (.I(_10497_),
    .Z(net18941));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18942 (.I(_10446_),
    .Z(net18942));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19019 (.I(net19018),
    .Z(net19019));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18946 (.I(_09840_),
    .Z(net18946));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18981 (.I(net18978),
    .Z(net18981));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18957 (.I(_06928_),
    .Z(net18957));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19052 (.I(net19038),
    .Z(net19052));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18948 (.I(_09744_),
    .Z(net18948));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18980 (.I(net18978),
    .Z(net18980));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18951 (.I(_16089_[0]),
    .Z(net18951));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18963 (.I(net18961),
    .Z(net18963));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer140 (.I(_16007_[0]),
    .Z(net527));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place18954 (.I(_16076_[0]),
    .Z(net18954));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18955 (.I(_16075_[0]),
    .Z(net18955));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18956 (.I(_06971_),
    .Z(net18956));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place18958 (.I(_16170_[0]),
    .Z(net18958));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18961 (.I(_06827_),
    .Z(net18961));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18994 (.I(_06782_),
    .Z(net18994));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19014 (.I(net19012),
    .Z(net19014));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18245 (.I(_14435_),
    .Z(net18245));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18997 (.I(_06763_),
    .Z(net18997));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18996 (.I(_06763_),
    .Z(net18996));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19028 (.I(net19022),
    .Z(net19028));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19119 (.I(_03946_),
    .Z(net19119));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17587 (.I(_11293_),
    .Z(net17587));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19050 (.I(net19038),
    .Z(net19050));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19038 (.I(_05322_),
    .Z(net19038));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19039 (.I(net19038),
    .Z(net19039));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19049 (.I(net19038),
    .Z(net19049));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19048 (.I(net19038),
    .Z(net19048));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19047 (.I(net19038),
    .Z(net19047));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19000 (.I(net18998),
    .Z(net19000));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18999 (.I(net18998),
    .Z(net18999));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17543 (.I(_13136_),
    .Z(net17543));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19085 (.I(net19082),
    .Z(net19085));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19084 (.I(net19083),
    .Z(net19084));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19083 (.I(net19082),
    .Z(net19083));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19003 (.I(_06162_),
    .Z(net19003));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19002 (.I(_06299_),
    .Z(net19002));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19004 (.I(_06162_),
    .Z(net19004));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19106 (.I(net19097),
    .Z(net19106));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19009 (.I(_16138_[0]),
    .Z(net19009));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19010 (.I(net19009),
    .Z(net19010));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19007 (.I(_06075_),
    .Z(net19007));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19055 (.I(_05303_),
    .Z(net19055));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19006 (.I(_06157_),
    .Z(net19006));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19011 (.I(_06032_),
    .Z(net19011));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19095 (.I(_04599_),
    .Z(net19095));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19105 (.I(net19097),
    .Z(net19105));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19104 (.I(net19103),
    .Z(net19104));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19060 (.I(net19059),
    .Z(net19060));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19059 (.I(_16111_[0]),
    .Z(net19059));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19016 (.I(_05450_),
    .Z(net19016));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19012 (.I(_05987_),
    .Z(net19012));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19041 (.I(net19038),
    .Z(net19041));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20432 (.I(_14517_),
    .Z(net20432));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19015 (.I(_05450_),
    .Z(net19015));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19044 (.I(net19038),
    .Z(net19044));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19022 (.I(_05342_),
    .Z(net19022));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19023 (.I(net19022),
    .Z(net19023));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19021 (.I(net19020),
    .Z(net19021));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19005 (.I(_06157_),
    .Z(net19005));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19077 (.I(_04655_),
    .Z(net19077));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19008 (.I(_16138_[0]),
    .Z(net19008));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19020 (.I(_05361_),
    .Z(net19020));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19013 (.I(net19012),
    .Z(net19013));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19040 (.I(net19038),
    .Z(net19040));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19018 (.I(_16106_[0]),
    .Z(net19018));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19017 (.I(_16106_[0]),
    .Z(net19017));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19046 (.I(net19038),
    .Z(net19046));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19058 (.I(_05303_),
    .Z(net19058));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19043 (.I(net19041),
    .Z(net19043));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19042 (.I(net19041),
    .Z(net19042));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19045 (.I(net19038),
    .Z(net19045));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19057 (.I(_05303_),
    .Z(net19057));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19056 (.I(_05303_),
    .Z(net19056));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19171 (.I(_15965_[0]),
    .Z(net19171));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19118 (.I(_03946_),
    .Z(net19118));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19117 (.I(_03946_),
    .Z(net19117));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19116 (.I(_03946_),
    .Z(net19116));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19115 (.I(_03946_),
    .Z(net19115));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19103 (.I(net19097),
    .Z(net19103));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19075 (.I(_04655_),
    .Z(net19075));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19081 (.I(_04630_),
    .Z(net19081));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19061 (.I(_05060_),
    .Z(net19061));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19074 (.I(_04704_),
    .Z(net19074));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19114 (.I(_03946_),
    .Z(net19114));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19266 (.I(net19263),
    .Z(net19266));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19160 (.I(_03122_),
    .Z(net19160));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19163 (.I(net19160),
    .Z(net19163));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19162 (.I(net19160),
    .Z(net19162));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19097 (.I(_04592_),
    .Z(net19097));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19154 (.I(_03151_),
    .Z(net19154));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19122 (.I(_16037_[0]),
    .Z(net19122));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19102 (.I(net19101),
    .Z(net19102));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19072 (.I(_04705_),
    .Z(net19072));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19101 (.I(net19097),
    .Z(net19101));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19100 (.I(net19097),
    .Z(net19100));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19123 (.I(net19122),
    .Z(net19123));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19153 (.I(_03151_),
    .Z(net19153));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19152 (.I(net19149),
    .Z(net19152));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19132 (.I(_03833_),
    .Z(net19132));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19099 (.I(net19098),
    .Z(net19099));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19065 (.I(_04752_),
    .Z(net19065));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19069 (.I(net19068),
    .Z(net19069));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19067 (.I(_04723_),
    .Z(net19067));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19062 (.I(_04769_),
    .Z(net19062));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19064 (.I(_04752_),
    .Z(net19064));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19066 (.I(_04723_),
    .Z(net19066));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19068 (.I(_04708_),
    .Z(net19068));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19071 (.I(_04705_),
    .Z(net19071));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19070 (.I(_04707_),
    .Z(net19070));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19073 (.I(_04704_),
    .Z(net19073));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19131 (.I(_03833_),
    .Z(net19131));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19082 (.I(_04605_),
    .Z(net19082));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19079 (.I(_04632_),
    .Z(net19079));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19078 (.I(_04632_),
    .Z(net19078));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19080 (.I(_04630_),
    .Z(net19080));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19108 (.I(net19097),
    .Z(net19108));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19112 (.I(_03946_),
    .Z(net19112));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19315 (.I(net19303),
    .Z(net19315));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19124 (.I(_16037_[0]),
    .Z(net19124));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19126 (.I(net403),
    .Z(net19126));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19514 (.I(_06056_),
    .Z(net19514));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19130 (.I(_03833_),
    .Z(net19130));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19121 (.I(_03946_),
    .Z(net19121));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19127 (.I(_03833_),
    .Z(net19127));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19128 (.I(_03833_),
    .Z(net19128));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19316 (.I(net19303),
    .Z(net19316));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19314 (.I(net647),
    .Z(net19314));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19529 (.I(net19515),
    .Z(net19529));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19125 (.I(net404),
    .Z(net19125));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19167 (.I(net19160),
    .Z(net19167));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19161 (.I(net19160),
    .Z(net19161));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19166 (.I(net19160),
    .Z(net19166));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19262 (.I(_15807_[0]),
    .Z(net19262));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19313 (.I(net19303),
    .Z(net19313));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19148 (.I(net19147),
    .Z(net19148));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19165 (.I(net19160),
    .Z(net19165));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19164 (.I(net19160),
    .Z(net19164));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19261 (.I(net19259),
    .Z(net19261));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19149 (.I(_03151_),
    .Z(net19149));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19257 (.I(net19256),
    .Z(net19257));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19144 (.I(_03193_),
    .Z(net19144));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19139 (.I(net19138),
    .Z(net19139));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19256 (.I(_13669_),
    .Z(net19256));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19183 (.I(_01777_),
    .Z(net19183));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19135 (.I(net19133),
    .Z(net19135));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19600 (.I(net19588),
    .Z(net19600));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19129 (.I(_03833_),
    .Z(net19129));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19176 (.I(net19175),
    .Z(net19176));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19136 (.I(_16043_[0]),
    .Z(net19136));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19179 (.I(_15976_[0]),
    .Z(net19179));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19240 (.I(net19233),
    .Z(net19240));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19239 (.I(net19233),
    .Z(net19239));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19134 (.I(net19133),
    .Z(net19134));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19133 (.I(_16048_[0]),
    .Z(net19133));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19137 (.I(_16043_[0]),
    .Z(net19137));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19138 (.I(_16043_[0]),
    .Z(net19138));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19151 (.I(net19149),
    .Z(net19151));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19140 (.I(_03340_),
    .Z(net19140));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19141 (.I(net19140),
    .Z(net19141));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19170 (.I(net19168),
    .Z(net19170));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19145 (.I(_16001_[0]),
    .Z(net19145));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19142 (.I(_03284_),
    .Z(net19142));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19147 (.I(_16001_[0]),
    .Z(net19147));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19168 (.I(_03122_),
    .Z(net19168));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19146 (.I(_16001_[0]),
    .Z(net19146));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19143 (.I(_03193_),
    .Z(net19143));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19169 (.I(net19168),
    .Z(net19169));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19150 (.I(net19149),
    .Z(net19150));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19238 (.I(net19233),
    .Z(net19238));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19237 (.I(net19233),
    .Z(net19237));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19174 (.I(_15966_[0]),
    .Z(net19174));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19175 (.I(_15966_[0]),
    .Z(net19175));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place19178 (.I(net19177),
    .Z(net19178));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19312 (.I(net647),
    .Z(net19312));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19271 (.I(_12947_),
    .Z(net19271));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19270 (.I(_12947_),
    .Z(net19270));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19512 (.I(_06056_),
    .Z(net19512));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19223 (.I(_14488_),
    .Z(net19223));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place19212 (.I(_15076_),
    .Z(net19212));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19209 (.I(net651),
    .Z(net19209));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19194 (.I(net19192),
    .Z(net19194));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19192 (.I(_01614_),
    .Z(net19192));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19195 (.I(net19192),
    .Z(net19195));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19191 (.I(net19189),
    .Z(net19191));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19273 (.I(_15770_[0]),
    .Z(net19273));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19304 (.I(net647),
    .Z(net19304));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19180 (.I(_15971_[0]),
    .Z(net19180));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19181 (.I(net442),
    .Z(net19181));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19303 (.I(_12128_),
    .Z(net19303));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19274 (.I(net19273),
    .Z(net19274));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19300 (.I(net19297),
    .Z(net19300));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19275 (.I(net19273),
    .Z(net19275));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19283 (.I(_12861_),
    .Z(net19283));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19249 (.I(_13669_),
    .Z(net19249));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19198 (.I(net19197),
    .Z(net19198));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19190 (.I(net19189),
    .Z(net19190));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19182 (.I(_01777_),
    .Z(net19182));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19197 (.I(net19196),
    .Z(net19197));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19188 (.I(_01643_),
    .Z(net19188));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19196 (.I(_15898_[0]),
    .Z(net19196));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19199 (.I(net19197),
    .Z(net19199));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19189 (.I(_01619_),
    .Z(net19189));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19193 (.I(net19192),
    .Z(net19193));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19269 (.I(_12947_),
    .Z(net19269));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19268 (.I(net19267),
    .Z(net19268));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19311 (.I(net647),
    .Z(net19311));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19226 (.I(net19225),
    .Z(net19226));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19227 (.I(net19224),
    .Z(net19227));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19208 (.I(net19207),
    .Z(net19208));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19228 (.I(net19224),
    .Z(net19228));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19248 (.I(_13669_),
    .Z(net19248));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19251 (.I(_13669_),
    .Z(net19251));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19201 (.I(_00987_),
    .Z(net19201));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19255 (.I(_13669_),
    .Z(net19255));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19207 (.I(_15865_[0]),
    .Z(net19207));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19205 (.I(net19204),
    .Z(net19205));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19220 (.I(_14495_),
    .Z(net19220));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19200 (.I(_01019_),
    .Z(net19200));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19242 (.I(_15802_[0]),
    .Z(net19242));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19310 (.I(net647),
    .Z(net19310));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19258 (.I(_13669_),
    .Z(net19258));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19206 (.I(_15903_[0]),
    .Z(net19206));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19254 (.I(_13669_),
    .Z(net19254));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19202 (.I(net19201),
    .Z(net19202));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19232 (.I(_13800_),
    .Z(net19232));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19272 (.I(net19271),
    .Z(net19272));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19234 (.I(net19233),
    .Z(net19234));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19217 (.I(_14521_),
    .Z(net19217));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19203 (.I(_00948_),
    .Z(net19203));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19210 (.I(_15874_[0]),
    .Z(net19210));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19218 (.I(net19217),
    .Z(net19218));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19204 (.I(_15903_[0]),
    .Z(net19204));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19211 (.I(net19210),
    .Z(net19211));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19231 (.I(_13808_),
    .Z(net19231));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19235 (.I(net19233),
    .Z(net19235));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19214 (.I(net19213),
    .Z(net19214));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19213 (.I(_14581_),
    .Z(net19213));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19253 (.I(net19252),
    .Z(net19253));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19215 (.I(_14555_),
    .Z(net19215));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19216 (.I(_14521_),
    .Z(net19216));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19252 (.I(_13669_),
    .Z(net19252));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19247 (.I(_13714_),
    .Z(net19247));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19225 (.I(net19224),
    .Z(net19225));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19222 (.I(_14488_),
    .Z(net19222));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19219 (.I(_14495_),
    .Z(net19219));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19221 (.I(_14488_),
    .Z(net19221));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19224 (.I(_15834_[0]),
    .Z(net19224));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19230 (.I(net19229),
    .Z(net19230));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19229 (.I(_15839_[0]),
    .Z(net19229));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19241 (.I(_13779_),
    .Z(net19241));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19246 (.I(net19244),
    .Z(net19246));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19233 (.I(_13790_),
    .Z(net19233));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19243 (.I(net430),
    .Z(net19243));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19265 (.I(net19263),
    .Z(net19265));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19263 (.I(_12947_),
    .Z(net19263));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19264 (.I(net19263),
    .Z(net19264));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19260 (.I(net19259),
    .Z(net19260));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19278 (.I(net19277),
    .Z(net19278));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19411 (.I(net19400),
    .Z(net19411));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19331 (.I(_12052_),
    .Z(net19331));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place19322 (.I(net19317),
    .Z(net19322));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19321 (.I(net19317),
    .Z(net19321));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19309 (.I(net19303),
    .Z(net19309));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19245 (.I(net19244),
    .Z(net19245));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19244 (.I(_13714_),
    .Z(net19244));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19308 (.I(net19303),
    .Z(net19308));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19250 (.I(_13669_),
    .Z(net19250));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19307 (.I(net19303),
    .Z(net19307));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19320 (.I(net19317),
    .Z(net19320));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19277 (.I(net19273),
    .Z(net19277));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19276 (.I(net19275),
    .Z(net19276));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19285 (.I(_15769_[0]),
    .Z(net19285));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19281 (.I(_12861_),
    .Z(net19281));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19404 (.I(net19400),
    .Z(net19404));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19783 (.I(net19780),
    .Z(net19783));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19319 (.I(net19317),
    .Z(net19319));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19318 (.I(net19317),
    .Z(net19318));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19295 (.I(net19294),
    .Z(net19295));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19294 (.I(_15778_[0]),
    .Z(net19294));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19290 (.I(_12856_),
    .Z(net19290));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19293 (.I(_12856_),
    .Z(net19293));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19289 (.I(net19287),
    .Z(net19289));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19280 (.I(net19279),
    .Z(net19280));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19286 (.I(net19285),
    .Z(net19286));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19279 (.I(_12861_),
    .Z(net19279));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19292 (.I(_12856_),
    .Z(net19292));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19291 (.I(_12856_),
    .Z(net19291));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19284 (.I(_15769_[0]),
    .Z(net19284));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19343 (.I(net19341),
    .Z(net19343));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19361 (.I(net19352),
    .Z(net19361));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19287 (.I(_12856_),
    .Z(net19287));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19288 (.I(net19287),
    .Z(net19288));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19370 (.I(net19363),
    .Z(net19370));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19410 (.I(net19409),
    .Z(net19410));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19371 (.I(net19363),
    .Z(net19371));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19298 (.I(net19297),
    .Z(net19298));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19317 (.I(_12095_),
    .Z(net19317));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19328 (.I(net19317),
    .Z(net19328));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19385 (.I(net19374),
    .Z(net19385));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19384 (.I(net19383),
    .Z(net19384));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19338 (.I(_12047_),
    .Z(net19338));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19299 (.I(net19297),
    .Z(net19299));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19296 (.I(_15778_[0]),
    .Z(net19296));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19337 (.I(_12047_),
    .Z(net19337));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19334 (.I(net19333),
    .Z(net19334));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19372 (.I(net19363),
    .Z(net19372));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19409 (.I(net19400),
    .Z(net19409));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19326 (.I(net19317),
    .Z(net19326));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19325 (.I(net19317),
    .Z(net19325));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19297 (.I(_15775_[0]),
    .Z(net19297));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19302 (.I(net19301),
    .Z(net19302));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19301 (.I(net646),
    .Z(net19301));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19408 (.I(net19407),
    .Z(net19408));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place19324 (.I(net19322),
    .Z(net19324));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19323 (.I(net19322),
    .Z(net19323));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19327 (.I(net19317),
    .Z(net19327));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19330 (.I(_12052_),
    .Z(net19330));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19407 (.I(net19400),
    .Z(net19407));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19329 (.I(_12052_),
    .Z(net19329));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19360 (.I(net19359),
    .Z(net19360));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19359 (.I(net19352),
    .Z(net19359));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19358 (.I(net19352),
    .Z(net19358));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19339 (.I(_15746_[0]),
    .Z(net19339));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19351 (.I(net19341),
    .Z(net19351));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19357 (.I(net19352),
    .Z(net19357));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19356 (.I(net19352),
    .Z(net19356));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19355 (.I(net19352),
    .Z(net19355));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19354 (.I(net19352),
    .Z(net19354));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20679 (.I(net20669),
    .Z(net20679));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21513 (.I(net21490),
    .Z(net21513));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21512 (.I(net21490),
    .Z(net21512));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19341 (.I(_11333_),
    .Z(net19341));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21511 (.I(net21501),
    .Z(net21511));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19782 (.I(net19780),
    .Z(net19782));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19335 (.I(_12047_),
    .Z(net19335));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19336 (.I(_12047_),
    .Z(net19336));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19350 (.I(net19341),
    .Z(net19350));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19349 (.I(net19341),
    .Z(net19349));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19781 (.I(net19780),
    .Z(net19781));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19383 (.I(net19374),
    .Z(net19383));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19382 (.I(net19374),
    .Z(net19382));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19353 (.I(net19352),
    .Z(net19353));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19348 (.I(net19341),
    .Z(net19348));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19347 (.I(net19341),
    .Z(net19347));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19346 (.I(net19341),
    .Z(net19346));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19847 (.I(net19840),
    .Z(net19847));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19696 (.I(_02342_),
    .Z(net19696));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19381 (.I(net19374),
    .Z(net19381));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19846 (.I(net19840),
    .Z(net19846));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19821 (.I(net19820),
    .Z(net19821));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19362 (.I(net19352),
    .Z(net19362));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19380 (.I(net19374),
    .Z(net19380));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19368 (.I(net19363),
    .Z(net19368));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19367 (.I(net19363),
    .Z(net19367));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19366 (.I(net19363),
    .Z(net19366));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19352 (.I(_11317_),
    .Z(net19352));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19342 (.I(net19341),
    .Z(net19342));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19365 (.I(net19363),
    .Z(net19365));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19364 (.I(net19363),
    .Z(net19364));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19363 (.I(_11296_),
    .Z(net19363));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19379 (.I(net19374),
    .Z(net19379));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19378 (.I(net19374),
    .Z(net19378));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19377 (.I(net19374),
    .Z(net19377));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19406 (.I(net506),
    .Z(net19406));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19376 (.I(net19374),
    .Z(net19376));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19369 (.I(net19363),
    .Z(net19369));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19375 (.I(net19374),
    .Z(net19375));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19779 (.I(_14459_),
    .Z(net19779));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19405 (.I(net19400),
    .Z(net19405));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19394 (.I(_11237_),
    .Z(net19394));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19397 (.I(_11237_),
    .Z(net19397));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19396 (.I(_11237_),
    .Z(net19396));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19395 (.I(_11237_),
    .Z(net19395));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19392 (.I(net19386),
    .Z(net19392));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19391 (.I(net19386),
    .Z(net19391));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19390 (.I(net19386),
    .Z(net19390));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19389 (.I(net19386),
    .Z(net19389));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19388 (.I(net19386),
    .Z(net19388));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19426 (.I(_15673_[0]),
    .Z(net19426));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19486 (.I(net19483),
    .Z(net19486));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19485 (.I(net19483),
    .Z(net19485));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19393 (.I(_11237_),
    .Z(net19393));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19415 (.I(net19413),
    .Z(net19415));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19414 (.I(net19413),
    .Z(net19414));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19403 (.I(net505),
    .Z(net19403));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19413 (.I(_10492_),
    .Z(net19413));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19423 (.I(net19413),
    .Z(net19423));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19412 (.I(_10492_),
    .Z(net19412));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20451 (.I(_09847_),
    .Z(net20451));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19475 (.I(_06109_),
    .Z(net19475));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place19425 (.I(net494),
    .Z(net19425));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19474 (.I(_06109_),
    .Z(net19474));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19526 (.I(net19525),
    .Z(net19526));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19472 (.I(_06109_),
    .Z(net19472));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19464 (.I(net19463),
    .Z(net19464));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19525 (.I(net19515),
    .Z(net19525));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19454 (.I(net19446),
    .Z(net19454));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19402 (.I(net507),
    .Z(net19402));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19399 (.I(net19398),
    .Z(net19399));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19398 (.I(_15674_[0]),
    .Z(net19398));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19460 (.I(_06762_),
    .Z(net19460));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19429 (.I(_15679_[0]),
    .Z(net19429));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19453 (.I(net19450),
    .Z(net19453));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19400 (.I(_10503_),
    .Z(net19400));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19420 (.I(net19413),
    .Z(net19420));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19452 (.I(net19450),
    .Z(net19452));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19419 (.I(net19418),
    .Z(net19419));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19416 (.I(net19413),
    .Z(net19416));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19401 (.I(net19400),
    .Z(net19401));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19422 (.I(net19413),
    .Z(net19422));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19418 (.I(net19413),
    .Z(net19418));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19417 (.I(net19413),
    .Z(net19417));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19421 (.I(net19413),
    .Z(net19421));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19511 (.I(net19510),
    .Z(net19511));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19451 (.I(net19450),
    .Z(net19451));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19427 (.I(net495),
    .Z(net19427));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19524 (.I(net19515),
    .Z(net19524));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer111 (.I(_10622_),
    .Z(net498));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19473 (.I(_06109_),
    .Z(net19473));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19490 (.I(net19487),
    .Z(net19490));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19428 (.I(net496),
    .Z(net19428));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19523 (.I(net19515),
    .Z(net19523));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19695 (.I(net19686),
    .Z(net19695));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19489 (.I(net19487),
    .Z(net19489));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19471 (.I(_06109_),
    .Z(net19471));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19470 (.I(_06109_),
    .Z(net19470));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19694 (.I(net19686),
    .Z(net19694));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19559 (.I(_05335_),
    .Z(net19559));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19693 (.I(net19686),
    .Z(net19693));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19853 (.I(net19840),
    .Z(net19853));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19449 (.I(net19448),
    .Z(net19449));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19668 (.I(_03078_),
    .Z(net19668));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19459 (.I(_06762_),
    .Z(net19459));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19448 (.I(net19446),
    .Z(net19448));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19431 (.I(net502),
    .Z(net19431));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19430 (.I(net19429),
    .Z(net19430));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19654 (.I(net19650),
    .Z(net19654));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19447 (.I(net19446),
    .Z(net19447));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19432 (.I(_10261_),
    .Z(net19432));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19522 (.I(net19515),
    .Z(net19522));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19505 (.I(_06056_),
    .Z(net19505));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19488 (.I(net19487),
    .Z(net19488));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19510 (.I(_06056_),
    .Z(net19510));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19484 (.I(net19483),
    .Z(net19484));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19467 (.I(_06109_),
    .Z(net19467));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19483 (.I(_06090_),
    .Z(net19483));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19436 (.I(_09774_),
    .Z(net19436));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19434 (.I(_09883_),
    .Z(net19434));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19444 (.I(_08681_),
    .Z(net19444));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19433 (.I(_09888_),
    .Z(net19433));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19458 (.I(_06762_),
    .Z(net19458));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19446 (.I(_06800_),
    .Z(net19446));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19469 (.I(_06109_),
    .Z(net19469));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19468 (.I(_06109_),
    .Z(net19468));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19439 (.I(_09298_),
    .Z(net19439));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19442 (.I(_08763_),
    .Z(net19442));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19438 (.I(_09743_),
    .Z(net19438));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19437 (.I(_09753_),
    .Z(net19437));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19435 (.I(_09865_),
    .Z(net19435));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19457 (.I(net388),
    .Z(net19457));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19440 (.I(_09296_),
    .Z(net19440));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19441 (.I(_09289_),
    .Z(net19441));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19443 (.I(_08751_),
    .Z(net19443));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19445 (.I(_08155_),
    .Z(net19445));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19465 (.I(net391),
    .Z(net19465));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19463 (.I(_06762_),
    .Z(net19463));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19487 (.I(_06071_),
    .Z(net19487));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19508 (.I(net19505),
    .Z(net19508));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19504 (.I(_06056_),
    .Z(net19504));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19507 (.I(net19505),
    .Z(net19507));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19506 (.I(net19505),
    .Z(net19506));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19509 (.I(_06056_),
    .Z(net19509));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19482 (.I(net19476),
    .Z(net19482));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19481 (.I(net19476),
    .Z(net19481));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19480 (.I(net19476),
    .Z(net19480));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19466 (.I(_06109_),
    .Z(net19466));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19479 (.I(net19476),
    .Z(net19479));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19478 (.I(net19476),
    .Z(net19478));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19477 (.I(net19476),
    .Z(net19477));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19476 (.I(_06090_),
    .Z(net19476));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19521 (.I(net19515),
    .Z(net19521));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19503 (.I(_06056_),
    .Z(net19503));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19502 (.I(net19497),
    .Z(net19502));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19496 (.I(_06071_),
    .Z(net19496));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19495 (.I(net19493),
    .Z(net19495));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19494 (.I(net19493),
    .Z(net19494));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19493 (.I(_06071_),
    .Z(net19493));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19501 (.I(net19497),
    .Z(net19501));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19500 (.I(net19497),
    .Z(net19500));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19497 (.I(_06056_),
    .Z(net19497));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19499 (.I(net19497),
    .Z(net19499));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19498 (.I(net19497),
    .Z(net19498));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19520 (.I(net19515),
    .Z(net19520));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19519 (.I(net19515),
    .Z(net19519));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19653 (.I(net19650),
    .Z(net19653));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19518 (.I(net19515),
    .Z(net19518));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19517 (.I(net19515),
    .Z(net19517));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19516 (.I(net19515),
    .Z(net19516));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19515 (.I(_06050_),
    .Z(net19515));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19527 (.I(net19515),
    .Z(net19527));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20416 (.I(net20412),
    .Z(net20416));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20450 (.I(net20449),
    .Z(net20450));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20442 (.I(_12196_),
    .Z(net20442));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20441 (.I(_12314_),
    .Z(net20441));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19558 (.I(net19546),
    .Z(net19558));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19557 (.I(net19546),
    .Z(net19557));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19556 (.I(net19546),
    .Z(net19556));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19555 (.I(net19546),
    .Z(net19555));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19530 (.I(_06030_),
    .Z(net19530));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19984 (.I(net19975),
    .Z(net19984));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19554 (.I(net19546),
    .Z(net19554));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19533 (.I(net19532),
    .Z(net19533));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19532 (.I(_06030_),
    .Z(net19532));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19599 (.I(net19588),
    .Z(net19599));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19531 (.I(net19530),
    .Z(net19531));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20460 (.I(_09742_),
    .Z(net20460));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19553 (.I(net19546),
    .Z(net19553));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19550 (.I(net19546),
    .Z(net19550));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19552 (.I(net19546),
    .Z(net19552));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19551 (.I(net19546),
    .Z(net19551));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19541 (.I(_06024_),
    .Z(net19541));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19628 (.I(net19627),
    .Z(net19628));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19540 (.I(_06024_),
    .Z(net19540));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19537 (.I(_06024_),
    .Z(net19537));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19534 (.I(_16137_[0]),
    .Z(net19534));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19539 (.I(net19538),
    .Z(net19539));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19598 (.I(net19588),
    .Z(net19598));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19597 (.I(net19588),
    .Z(net19597));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19538 (.I(_06024_),
    .Z(net19538));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20695 (.I(net20685),
    .Z(net20695));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19580 (.I(net19571),
    .Z(net19580));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19581 (.I(net19571),
    .Z(net19581));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19579 (.I(net19571),
    .Z(net19579));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19578 (.I(net19571),
    .Z(net19578));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19577 (.I(net19571),
    .Z(net19577));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19569 (.I(_05302_),
    .Z(net19569));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19549 (.I(net19546),
    .Z(net19549));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19542 (.I(_16146_[0]),
    .Z(net19542));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19536 (.I(_06024_),
    .Z(net19536));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19535 (.I(_06024_),
    .Z(net19535));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19545 (.I(net19544),
    .Z(net19545));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19566 (.I(net19565),
    .Z(net19566));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20765 (.I(net20757),
    .Z(net20765));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20602 (.I(_07330_),
    .Z(net20602));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20764 (.I(net20757),
    .Z(net20764));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20614 (.I(_07330_),
    .Z(net20614));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20613 (.I(_07330_),
    .Z(net20613));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20612 (.I(net20611),
    .Z(net20612));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20611 (.I(_07330_),
    .Z(net20611));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20588 (.I(net20587),
    .Z(net20588));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20578 (.I(_07630_),
    .Z(net20578));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19548 (.I(net19546),
    .Z(net19548));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19544 (.I(net19543),
    .Z(net19544));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19543 (.I(_16146_[0]),
    .Z(net19543));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19560 (.I(net19559),
    .Z(net19560));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20490 (.I(_09198_),
    .Z(net20490));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19565 (.I(_16105_[0]),
    .Z(net19565));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19563 (.I(net19559),
    .Z(net19563));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19546 (.I(_05367_),
    .Z(net19546));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19547 (.I(net19546),
    .Z(net19547));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19562 (.I(net19559),
    .Z(net19562));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20439 (.I(_13616_),
    .Z(net20439));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21082 (.I(_10378_),
    .Z(net21082));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19927 (.I(_06414_),
    .Z(net19927));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19639 (.I(net19630),
    .Z(net19639));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19595 (.I(net19588),
    .Z(net19595));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19564 (.I(_16105_[0]),
    .Z(net19564));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19582 (.I(_04651_),
    .Z(net19582));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19587 (.I(_04651_),
    .Z(net19587));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19638 (.I(net19630),
    .Z(net19638));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19576 (.I(net19571),
    .Z(net19576));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19575 (.I(net19571),
    .Z(net19575));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19637 (.I(net19630),
    .Z(net19637));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19570 (.I(_16114_[0]),
    .Z(net19570));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19567 (.I(_05302_),
    .Z(net19567));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19568 (.I(_05302_),
    .Z(net19568));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20262 (.I(net20258),
    .Z(net20262));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19616 (.I(_04568_),
    .Z(net19616));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19607 (.I(net19606),
    .Z(net19607));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19594 (.I(net19593),
    .Z(net19594));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19593 (.I(net19588),
    .Z(net19593));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19592 (.I(net19588),
    .Z(net19592));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19586 (.I(_04651_),
    .Z(net19586));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19585 (.I(net19584),
    .Z(net19585));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19574 (.I(net19571),
    .Z(net19574));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19573 (.I(net19571),
    .Z(net19573));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19926 (.I(_06414_),
    .Z(net19926));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19571 (.I(_04674_),
    .Z(net19571));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20261 (.I(net20258),
    .Z(net20261));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20254 (.I(net20252),
    .Z(net20254));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19627 (.I(net19624),
    .Z(net19627));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19617 (.I(net512),
    .Z(net19617));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19982 (.I(net19975),
    .Z(net19982));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19981 (.I(net19975),
    .Z(net19981));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19584 (.I(_04651_),
    .Z(net19584));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19572 (.I(net19571),
    .Z(net19572));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19591 (.I(net19588),
    .Z(net19591));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19583 (.I(_04651_),
    .Z(net19583));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19596 (.I(net19588),
    .Z(net19596));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19980 (.I(net19975),
    .Z(net19980));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19590 (.I(net19588),
    .Z(net19590));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19589 (.I(net19588),
    .Z(net19589));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19979 (.I(net19978),
    .Z(net19979));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19640 (.I(_03878_),
    .Z(net19640));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19588 (.I(_04620_),
    .Z(net19588));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19606 (.I(_04574_),
    .Z(net19606));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19605 (.I(net19604),
    .Z(net19605));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19604 (.I(net19603),
    .Z(net19604));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19602 (.I(net509),
    .Z(net19602));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19601 (.I(_16074_[0]),
    .Z(net19601));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20418 (.I(_02422_),
    .Z(net20418));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19978 (.I(net19975),
    .Z(net19978));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19636 (.I(net19630),
    .Z(net19636));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19648 (.I(net19640),
    .Z(net19648));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19647 (.I(net19640),
    .Z(net19647));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19603 (.I(_04574_),
    .Z(net19603));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19646 (.I(net19640),
    .Z(net19646));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19645 (.I(net19640),
    .Z(net19645));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19767 (.I(net19766),
    .Z(net19767));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19613 (.I(_04568_),
    .Z(net19613));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19612 (.I(_04568_),
    .Z(net19612));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19634 (.I(net19630),
    .Z(net19634));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19615 (.I(_04568_),
    .Z(net19615));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19614 (.I(_04568_),
    .Z(net19614));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19609 (.I(_04571_),
    .Z(net19609));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19610 (.I(net510),
    .Z(net19610));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19608 (.I(_04571_),
    .Z(net19608));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19611 (.I(_04568_),
    .Z(net19611));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19936 (.I(_05457_),
    .Z(net19936));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19914 (.I(_06892_),
    .Z(net19914));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19895 (.I(_09295_),
    .Z(net19895));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19917 (.I(_06892_),
    .Z(net19917));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19951 (.I(net19950),
    .Z(net19951));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19859 (.I(net19857),
    .Z(net19859));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19619 (.I(net19618),
    .Z(net19619));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19644 (.I(net19640),
    .Z(net19644));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19621 (.I(_03993_),
    .Z(net19621));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19633 (.I(net19630),
    .Z(net19633));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19626 (.I(net19624),
    .Z(net19626));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19629 (.I(net19624),
    .Z(net19629));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19623 (.I(_03993_),
    .Z(net19623));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19652 (.I(net19650),
    .Z(net19652));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19823 (.I(_12051_),
    .Z(net19823));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19632 (.I(net19630),
    .Z(net19632));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19631 (.I(net19630),
    .Z(net19631));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19625 (.I(net19624),
    .Z(net19625));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19618 (.I(_16079_[0]),
    .Z(net19618));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19630 (.I(_03908_),
    .Z(net19630));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19620 (.I(_03993_),
    .Z(net19620));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19622 (.I(_03993_),
    .Z(net19622));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19983 (.I(net19975),
    .Z(net19983));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20942 (.I(_12842_),
    .Z(net20942));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19624 (.I(_03921_),
    .Z(net19624));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19857 (.I(_10556_),
    .Z(net19857));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20678 (.I(net20669),
    .Z(net20678));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19685 (.I(net19678),
    .Z(net19685));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19674 (.I(_02496_),
    .Z(net19674));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19662 (.I(_03083_),
    .Z(net19662));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19660 (.I(_03083_),
    .Z(net19660));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19659 (.I(_03083_),
    .Z(net19659));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19655 (.I(_03083_),
    .Z(net19655));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19658 (.I(_03083_),
    .Z(net19658));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19635 (.I(net19630),
    .Z(net19635));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19657 (.I(_03083_),
    .Z(net19657));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19656 (.I(_03083_),
    .Z(net19656));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19651 (.I(net19650),
    .Z(net19651));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19643 (.I(net19640),
    .Z(net19643));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19642 (.I(net19640),
    .Z(net19642));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19641 (.I(net19640),
    .Z(net19641));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19977 (.I(net19975),
    .Z(net19977));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19650 (.I(_03832_),
    .Z(net19650));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19692 (.I(net19686),
    .Z(net19692));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19649 (.I(_03832_),
    .Z(net19649));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19661 (.I(net19660),
    .Z(net19661));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19820 (.I(net19809),
    .Z(net19820));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19691 (.I(net19686),
    .Z(net19691));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19345 (.I(net19341),
    .Z(net19345));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19344 (.I(net19341),
    .Z(net19344));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19684 (.I(net19678),
    .Z(net19684));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19683 (.I(net19678),
    .Z(net19683));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19669 (.I(_16012_[0]),
    .Z(net19669));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19852 (.I(net19840),
    .Z(net19852));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19667 (.I(_03078_),
    .Z(net19667));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19666 (.I(net19665),
    .Z(net19666));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19675 (.I(_02496_),
    .Z(net19675));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19665 (.I(_03078_),
    .Z(net19665));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19664 (.I(net19663),
    .Z(net19664));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19663 (.I(_03078_),
    .Z(net19663));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19333 (.I(_15737_[0]),
    .Z(net19333));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19766 (.I(_15172_),
    .Z(net19766));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19851 (.I(net19840),
    .Z(net19851));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19677 (.I(_02496_),
    .Z(net19677));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19670 (.I(net19669),
    .Z(net19670));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19676 (.I(_02496_),
    .Z(net19676));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19671 (.I(net19669),
    .Z(net19671));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19778 (.I(_14459_),
    .Z(net19778));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19682 (.I(net19678),
    .Z(net19682));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19681 (.I(net19678),
    .Z(net19681));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19673 (.I(_02496_),
    .Z(net19673));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19680 (.I(net19678),
    .Z(net19680));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19672 (.I(_02496_),
    .Z(net19672));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19819 (.I(net19809),
    .Z(net19819));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19690 (.I(net19686),
    .Z(net19690));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19710 (.I(net19702),
    .Z(net19710));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19689 (.I(net19686),
    .Z(net19689));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19688 (.I(net19686),
    .Z(net19688));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19687 (.I(net19686),
    .Z(net19687));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19679 (.I(net19678),
    .Z(net19679));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19678 (.I(_02440_),
    .Z(net19678));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19764 (.I(net19759),
    .Z(net19764));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19763 (.I(net19759),
    .Z(net19763));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19756 (.I(net19747),
    .Z(net19756));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19755 (.I(net19747),
    .Z(net19755));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19709 (.I(net19708),
    .Z(net19709));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19698 (.I(net19696),
    .Z(net19698));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19686 (.I(_02384_),
    .Z(net19686));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19850 (.I(net19840),
    .Z(net19850));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19848 (.I(net19840),
    .Z(net19848));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19697 (.I(net19696),
    .Z(net19697));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19717 (.I(net19715),
    .Z(net19717));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19716 (.I(net19715),
    .Z(net19716));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19715 (.I(_01663_),
    .Z(net19715));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19706 (.I(net19702),
    .Z(net19706));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19705 (.I(net19702),
    .Z(net19705));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19701 (.I(net19699),
    .Z(net19701));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19700 (.I(net19699),
    .Z(net19700));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19699 (.I(_02337_),
    .Z(net19699));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19708 (.I(net19702),
    .Z(net19708));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19340 (.I(net19339),
    .Z(net19340));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19373 (.I(net19363),
    .Z(net19373));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19386 (.I(_11243_),
    .Z(net19386));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19762 (.I(net19759),
    .Z(net19762));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19761 (.I(net19759),
    .Z(net19761));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19760 (.I(net19759),
    .Z(net19760));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19704 (.I(net19702),
    .Z(net19704));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19703 (.I(net19702),
    .Z(net19703));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19751 (.I(net19747),
    .Z(net19751));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19707 (.I(net19702),
    .Z(net19707));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19702 (.I(_01695_),
    .Z(net19702));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19387 (.I(net19386),
    .Z(net19387));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19374 (.I(_11288_),
    .Z(net19374));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19718 (.I(_01645_),
    .Z(net19718));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19259 (.I(_15807_[0]),
    .Z(net19259));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19561 (.I(net19559),
    .Z(net19561));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19730 (.I(net19725),
    .Z(net19730));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19236 (.I(net19233),
    .Z(net19236));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19185 (.I(_01777_),
    .Z(net19185));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19721 (.I(_15940_[0]),
    .Z(net19721));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19729 (.I(net19725),
    .Z(net19729));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19785 (.I(_14384_),
    .Z(net19785));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19711 (.I(_01684_),
    .Z(net19711));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19738 (.I(net19736),
    .Z(net19738));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19714 (.I(net19712),
    .Z(net19714));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19712 (.I(_01663_),
    .Z(net19712));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21096 (.I(_10367_),
    .Z(net21096));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19713 (.I(net19712),
    .Z(net19713));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19726 (.I(net19725),
    .Z(net19726));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19737 (.I(net19736),
    .Z(net19737));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19753 (.I(net19747),
    .Z(net19753));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19728 (.I(net19725),
    .Z(net19728));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19723 (.I(net467),
    .Z(net19723));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19727 (.I(net19725),
    .Z(net19727));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19720 (.I(net19719),
    .Z(net19720));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19719 (.I(_15929_[0]),
    .Z(net19719));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19187 (.I(net19186),
    .Z(net19187));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19734 (.I(net19731),
    .Z(net19734));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19186 (.I(_01777_),
    .Z(net19186));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19113 (.I(_03946_),
    .Z(net19113));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18648 (.I(_15930_[0]),
    .Z(net18648));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19733 (.I(net19731),
    .Z(net19733));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19098 (.I(net19097),
    .Z(net19098));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18650 (.I(net18649),
    .Z(net18650));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18649 (.I(_15930_[0]),
    .Z(net18649));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19111 (.I(_04576_),
    .Z(net19111));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19096 (.I(_04596_),
    .Z(net19096));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18711 (.I(net18708),
    .Z(net18711));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18703 (.I(_15333_),
    .Z(net18703));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18702 (.I(_15333_),
    .Z(net18702));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18685 (.I(net18684),
    .Z(net18685));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place18684 (.I(_00902_),
    .Z(net18684));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19754 (.I(net19747),
    .Z(net19754));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19722 (.I(net19721),
    .Z(net19722));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19736 (.I(net19735),
    .Z(net19736));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19725 (.I(_01034_),
    .Z(net19725));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19752 (.I(net19747),
    .Z(net19752));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18681 (.I(_00943_),
    .Z(net18681));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place19724 (.I(_01576_),
    .Z(net19724));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18674 (.I(net18670),
    .Z(net18674));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19732 (.I(net19731),
    .Z(net19732));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18673 (.I(net18670),
    .Z(net18673));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18653 (.I(_15935_[0]),
    .Z(net18653));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18647 (.I(_01623_),
    .Z(net18647));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18642 (.I(net18636),
    .Z(net18642));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18641 (.I(net18636),
    .Z(net18641));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18640 (.I(net18636),
    .Z(net18640));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21510 (.I(net21501),
    .Z(net21510));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19759 (.I(_15172_),
    .Z(net19759));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19749 (.I(net19747),
    .Z(net19749));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18699 (.I(net18684),
    .Z(net18699));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19731 (.I(_00878_),
    .Z(net19731));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19744 (.I(net19742),
    .Z(net19744));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place19735 (.I(_15897_[0]),
    .Z(net19735));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19739 (.I(_00873_),
    .Z(net19739));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19740 (.I(net19739),
    .Z(net19740));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19746 (.I(net19742),
    .Z(net19746));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19741 (.I(_15906_[0]),
    .Z(net19741));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19743 (.I(net19742),
    .Z(net19743));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19817 (.I(net19809),
    .Z(net19817));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19742 (.I(_15261_),
    .Z(net19742));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19745 (.I(net19742),
    .Z(net19745));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19795 (.I(_15842_[0]),
    .Z(net19795));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19777 (.I(_14459_),
    .Z(net19777));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19748 (.I(net19747),
    .Z(net19748));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19747 (.I(_15251_),
    .Z(net19747));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19750 (.I(net19747),
    .Z(net19750));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19773 (.I(_15117_),
    .Z(net19773));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19758 (.I(net19757),
    .Z(net19758));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19757 (.I(_15172_),
    .Z(net19757));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19765 (.I(_15172_),
    .Z(net19765));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19772 (.I(_15117_),
    .Z(net19772));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21509 (.I(net21501),
    .Z(net21509));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19768 (.I(_15122_),
    .Z(net19768));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19784 (.I(_14384_),
    .Z(net19784));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19816 (.I(net19814),
    .Z(net19816));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19769 (.I(_15117_),
    .Z(net19769));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19771 (.I(_15117_),
    .Z(net19771));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21508 (.I(net21501),
    .Z(net21508));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19770 (.I(_15117_),
    .Z(net19770));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18639 (.I(net18636),
    .Z(net18639));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18638 (.I(net18636),
    .Z(net18638));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18619 (.I(_01768_),
    .Z(net18619));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20677 (.I(net20669),
    .Z(net20677));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20676 (.I(net20669),
    .Z(net20676));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20675 (.I(net20669),
    .Z(net20675));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19776 (.I(_14459_),
    .Z(net19776));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19818 (.I(net19809),
    .Z(net19818));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19775 (.I(_14459_),
    .Z(net19775));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19774 (.I(_15074_),
    .Z(net19774));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19856 (.I(net19854),
    .Z(net19856));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18622 (.I(_01691_),
    .Z(net18622));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19813 (.I(net19809),
    .Z(net19813));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21507 (.I(net21501),
    .Z(net21507));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19794 (.I(_14379_),
    .Z(net19794));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19786 (.I(_15833_[0]),
    .Z(net19786));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19793 (.I(_14379_),
    .Z(net19793));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19792 (.I(_14379_),
    .Z(net19792));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19791 (.I(net19788),
    .Z(net19791));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21506 (.I(net21501),
    .Z(net21506));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19843 (.I(net19840),
    .Z(net19843));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19809 (.I(_12912_),
    .Z(net19809));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19832 (.I(_11376_),
    .Z(net19832));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19831 (.I(_11376_),
    .Z(net19831));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19787 (.I(net19786),
    .Z(net19787));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19780 (.I(_14384_),
    .Z(net19780));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19812 (.I(net19811),
    .Z(net19812));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19804 (.I(net19802),
    .Z(net19804));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 place19799 (.I(net19798),
    .Z(net19799));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19815 (.I(net19814),
    .Z(net19815));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19788 (.I(_14379_),
    .Z(net19788));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19790 (.I(net19788),
    .Z(net19790));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19789 (.I(net19788),
    .Z(net19789));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place19798 (.I(_13647_),
    .Z(net19798));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19800 (.I(net417),
    .Z(net19800));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19797 (.I(net19796),
    .Z(net19797));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19796 (.I(_15842_[0]),
    .Z(net19796));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19830 (.I(_11376_),
    .Z(net19830));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21134 (.I(_07372_),
    .Z(net21134));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19814 (.I(net19809),
    .Z(net19814));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19803 (.I(net19802),
    .Z(net19803));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19829 (.I(_11376_),
    .Z(net19829));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19828 (.I(_11376_),
    .Z(net19828));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21505 (.I(net21501),
    .Z(net21505));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19801 (.I(net604),
    .Z(net19801));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21504 (.I(net21501),
    .Z(net21504));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19845 (.I(net19840),
    .Z(net19845));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18617 (.I(_01774_),
    .Z(net18617));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18618 (.I(net18617),
    .Z(net18618));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18605 (.I(_02367_),
    .Z(net18605));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20694 (.I(net20685),
    .Z(net20694));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19855 (.I(net19854),
    .Z(net19855));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19805 (.I(_15810_[0]),
    .Z(net19805));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19810 (.I(net19809),
    .Z(net19810));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19802 (.I(_13642_),
    .Z(net19802));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19807 (.I(net19806),
    .Z(net19807));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19824 (.I(net19823),
    .Z(net19824));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19854 (.I(_10556_),
    .Z(net19854));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19806 (.I(_15810_[0]),
    .Z(net19806));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19811 (.I(net19809),
    .Z(net19811));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19822 (.I(_12855_),
    .Z(net19822));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19808 (.I(_12912_),
    .Z(net19808));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20760 (.I(net20757),
    .Z(net20760));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19844 (.I(net19840),
    .Z(net19844));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18470 (.I(_05452_),
    .Z(net18470));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18473 (.I(_05421_),
    .Z(net18473));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19918 (.I(_06892_),
    .Z(net19918));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19858 (.I(net19857),
    .Z(net19858));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place19826 (.I(_11991_),
    .Z(net19826));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19825 (.I(_12046_),
    .Z(net19825));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20733 (.I(net20721),
    .Z(net20733));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20736 (.I(net20721),
    .Z(net20736));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20674 (.I(net20669),
    .Z(net20674));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19839 (.I(_11183_),
    .Z(net19839));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19838 (.I(net19837),
    .Z(net19838));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19916 (.I(_06892_),
    .Z(net19916));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18440 (.I(_06919_),
    .Z(net18440));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20232 (.I(_15239_),
    .Z(net20232));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19947 (.I(net19945),
    .Z(net19947));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19864 (.I(_10532_),
    .Z(net19864));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19863 (.I(_10532_),
    .Z(net19863));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19862 (.I(_10532_),
    .Z(net19862));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19861 (.I(_10532_),
    .Z(net19861));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19949 (.I(net19945),
    .Z(net19949));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19868 (.I(_10445_),
    .Z(net19868));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19835 (.I(net19834),
    .Z(net19835));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19837 (.I(_15714_[0]),
    .Z(net19837));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20574 (.I(_07717_),
    .Z(net20574));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19827 (.I(_11376_),
    .Z(net19827));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19833 (.I(_11242_),
    .Z(net19833));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place19834 (.I(_15705_[0]),
    .Z(net19834));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19836 (.I(_11236_),
    .Z(net19836));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19939 (.I(_05457_),
    .Z(net19939));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19867 (.I(net19866),
    .Z(net19867));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19938 (.I(_05457_),
    .Z(net19938));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19866 (.I(_10445_),
    .Z(net19866));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21081 (.I(_10378_),
    .Z(net21081));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19842 (.I(net19840),
    .Z(net19842));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19841 (.I(net19840),
    .Z(net19841));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19948 (.I(net19945),
    .Z(net19948));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19919 (.I(_06892_),
    .Z(net19919));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19950 (.I(_04650_),
    .Z(net19950));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place19840 (.I(_10572_),
    .Z(net19840));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19860 (.I(_10532_),
    .Z(net19860));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19937 (.I(_05457_),
    .Z(net19937));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19865 (.I(_10532_),
    .Z(net19865));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19920 (.I(_06892_),
    .Z(net19920));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19976 (.I(net19975),
    .Z(net19976));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19957 (.I(_03831_),
    .Z(net19957));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19961 (.I(net19957),
    .Z(net19961));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19953 (.I(_03959_),
    .Z(net19953));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19970 (.I(net19969),
    .Z(net19970));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19966 (.I(_03210_),
    .Z(net19966));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20253 (.I(net20252),
    .Z(net20253));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20252 (.I(net20248),
    .Z(net20252));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19900 (.I(_09179_),
    .Z(net19900));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19877 (.I(_09863_),
    .Z(net19877));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19935 (.I(_05457_),
    .Z(net19935));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19930 (.I(_06108_),
    .Z(net19930));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19869 (.I(_10440_),
    .Z(net19869));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19870 (.I(net19869),
    .Z(net19870));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19886 (.I(_09772_),
    .Z(net19886));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place19888 (.I(_09752_),
    .Z(net19888));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19885 (.I(_09783_),
    .Z(net19885));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19876 (.I(_09880_),
    .Z(net19876));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19929 (.I(net19928),
    .Z(net19929));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19928 (.I(_06108_),
    .Z(net19928));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19871 (.I(_10135_),
    .Z(net19871));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19907 (.I(_08645_),
    .Z(net19907));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19875 (.I(_09880_),
    .Z(net19875));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19874 (.I(_10046_),
    .Z(net19874));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19872 (.I(_10120_),
    .Z(net19872));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19896 (.I(_09288_),
    .Z(net19896));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19878 (.I(_09862_),
    .Z(net19878));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19965 (.I(_03210_),
    .Z(net19965));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21080 (.I(_10378_),
    .Z(net21080));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19873 (.I(_10081_),
    .Z(net19873));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20250 (.I(net20248),
    .Z(net20250));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19923 (.I(net19921),
    .Z(net19923));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19922 (.I(net19921),
    .Z(net19922));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19880 (.I(_09842_),
    .Z(net19880));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19884 (.I(_09793_),
    .Z(net19884));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19889 (.I(_09752_),
    .Z(net19889));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19879 (.I(_09842_),
    .Z(net19879));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19881 (.I(_09836_),
    .Z(net19881));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19882 (.I(_09817_),
    .Z(net19882));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19883 (.I(_09811_),
    .Z(net19883));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19915 (.I(net19914),
    .Z(net19915));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19887 (.I(_09752_),
    .Z(net19887));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19894 (.I(_09295_),
    .Z(net19894));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19890 (.I(_09378_),
    .Z(net19890));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19891 (.I(_09364_),
    .Z(net19891));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19903 (.I(_08764_),
    .Z(net19903));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19893 (.I(_09327_),
    .Z(net19893));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19892 (.I(_09347_),
    .Z(net19892));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19902 (.I(_08795_),
    .Z(net19902));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19898 (.I(_09192_),
    .Z(net19898));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19897 (.I(_09273_),
    .Z(net19897));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19899 (.I(_09179_),
    .Z(net19899));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19901 (.I(_09164_),
    .Z(net19901));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20249 (.I(net20248),
    .Z(net20249));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19921 (.I(_06761_),
    .Z(net19921));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19904 (.I(_08734_),
    .Z(net19904));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19912 (.I(_08112_),
    .Z(net19912));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19905 (.I(_08680_),
    .Z(net19905));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19906 (.I(_08662_),
    .Z(net19906));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19908 (.I(_08237_),
    .Z(net19908));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19911 (.I(_08214_),
    .Z(net19911));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19910 (.I(_08217_),
    .Z(net19910));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19909 (.I(_08217_),
    .Z(net19909));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20243 (.I(_14485_),
    .Z(net20243));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20210 (.I(net20205),
    .Z(net20210));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19969 (.I(_03174_),
    .Z(net19969));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19913 (.I(_06892_),
    .Z(net19913));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19964 (.I(_03210_),
    .Z(net19964));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place19925 (.I(_06717_),
    .Z(net19925));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19990 (.I(net19985),
    .Z(net19990));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20061 (.I(net20059),
    .Z(net20061));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19924 (.I(_06723_),
    .Z(net19924));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19989 (.I(net19985),
    .Z(net19989));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19956 (.I(net19953),
    .Z(net19956));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19946 (.I(net19945),
    .Z(net19946));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19932 (.I(_05457_),
    .Z(net19932));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19988 (.I(net19985),
    .Z(net19988));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19941 (.I(_05419_),
    .Z(net19941));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19940 (.I(_05419_),
    .Z(net19940));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19934 (.I(_05457_),
    .Z(net19934));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19955 (.I(net19953),
    .Z(net19955));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19954 (.I(net19953),
    .Z(net19954));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19931 (.I(_06023_),
    .Z(net19931));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19933 (.I(_05457_),
    .Z(net19933));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20073 (.I(_09877_),
    .Z(net20073));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19975 (.I(_03174_),
    .Z(net19975));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19974 (.I(net19969),
    .Z(net19974));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19944 (.I(_05260_),
    .Z(net19944));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20075 (.I(_09831_),
    .Z(net20075));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19958 (.I(net19957),
    .Z(net19958));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19960 (.I(net19957),
    .Z(net19960));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19952 (.I(_04567_),
    .Z(net19952));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19942 (.I(_05301_),
    .Z(net19942));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19943 (.I(_05265_),
    .Z(net19943));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20069 (.I(_09923_),
    .Z(net20069));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20064 (.I(_10383_),
    .Z(net20064));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19987 (.I(net19985),
    .Z(net19987));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19962 (.I(_03210_),
    .Z(net19962));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19963 (.I(_03210_),
    .Z(net19963));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19959 (.I(net19957),
    .Z(net19959));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19968 (.I(_03210_),
    .Z(net19968));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19967 (.I(net19966),
    .Z(net19967));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19945 (.I(_04650_),
    .Z(net19945));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place19986 (.I(net19985),
    .Z(net19986));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19973 (.I(net19969),
    .Z(net19973));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20124 (.I(_08585_),
    .Z(net20124));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20136 (.I(_08120_),
    .Z(net20136));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21079 (.I(_10378_),
    .Z(net21079));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21078 (.I(_10378_),
    .Z(net21078));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20033 (.I(net20032),
    .Z(net20033));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20032 (.I(_13739_),
    .Z(net20032));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19996 (.I(_02458_),
    .Z(net19996));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19995 (.I(net19991),
    .Z(net19995));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19972 (.I(net19971),
    .Z(net19972));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20114 (.I(_08679_),
    .Z(net20114));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20022 (.I(_14378_),
    .Z(net20022));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20389 (.I(_06872_),
    .Z(net20389));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20269 (.I(_12969_),
    .Z(net20269));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20236 (.I(net20234),
    .Z(net20236));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20012 (.I(net20009),
    .Z(net20012));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19971 (.I(net19969),
    .Z(net19971));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19994 (.I(net19991),
    .Z(net19994));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place19991 (.I(_02458_),
    .Z(net19991));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place19985 (.I(_03143_),
    .Z(net19985));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19993 (.I(net19991),
    .Z(net19993));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20390 (.I(_06872_),
    .Z(net20390));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20251 (.I(net20248),
    .Z(net20251));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19992 (.I(net19991),
    .Z(net19992));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20005 (.I(net20000),
    .Z(net20005));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20003 (.I(net20000),
    .Z(net20003));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19999 (.I(_01180_),
    .Z(net19999));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place19997 (.I(_02319_),
    .Z(net19997));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20004 (.I(net20000),
    .Z(net20004));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21077 (.I(net21076),
    .Z(net21077));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20241 (.I(_14485_),
    .Z(net20241));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20226 (.I(net20222),
    .Z(net20226));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20192 (.I(_04691_),
    .Z(net20192));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20183 (.I(_05358_),
    .Z(net20183));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20173 (.I(_06739_),
    .Z(net20173));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20225 (.I(net20222),
    .Z(net20225));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20167 (.I(net20163),
    .Z(net20167));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20016 (.I(_14458_),
    .Z(net20016));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20157 (.I(_15641_[0]),
    .Z(net20157));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20002 (.I(net20000),
    .Z(net20002));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20001 (.I(net20000),
    .Z(net20001));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19998 (.I(_01180_),
    .Z(net19998));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20011 (.I(net20009),
    .Z(net20011));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20006 (.I(_00877_),
    .Z(net20006));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20020 (.I(_14409_),
    .Z(net20020));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20208 (.I(net20205),
    .Z(net20208));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20350 (.I(net20349),
    .Z(net20350));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20030 (.I(_13739_),
    .Z(net20030));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20277 (.I(net20275),
    .Z(net20277));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20273 (.I(_12198_),
    .Z(net20273));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20019 (.I(_14458_),
    .Z(net20019));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20018 (.I(_14458_),
    .Z(net20018));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20000 (.I(_00968_),
    .Z(net20000));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20029 (.I(_13739_),
    .Z(net20029));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20028 (.I(_13739_),
    .Z(net20028));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20027 (.I(_13739_),
    .Z(net20027));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20010 (.I(net20009),
    .Z(net20010));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20060 (.I(net20059),
    .Z(net20060));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20015 (.I(_15116_),
    .Z(net20015));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20014 (.I(net20013),
    .Z(net20014));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20007 (.I(_00872_),
    .Z(net20007));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20013 (.I(_15121_),
    .Z(net20013));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20008 (.I(_00827_),
    .Z(net20008));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20017 (.I(_14458_),
    .Z(net20017));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20156 (.I(_15642_[0]),
    .Z(net20156));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20059 (.I(_10555_),
    .Z(net20059));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20049 (.I(_11352_),
    .Z(net20049));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20009 (.I(_15189_),
    .Z(net20009));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20048 (.I(_11352_),
    .Z(net20048));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20021 (.I(_14383_),
    .Z(net20021));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20031 (.I(_13739_),
    .Z(net20031));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20802 (.I(net20794),
    .Z(net20802));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20190 (.I(_04739_),
    .Z(net20190));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20268 (.I(_12969_),
    .Z(net20268));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20263 (.I(_13015_),
    .Z(net20263));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20026 (.I(net20025),
    .Z(net20026));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20037 (.I(_13106_),
    .Z(net20037));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20054 (.I(net20052),
    .Z(net20054));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20025 (.I(_13739_),
    .Z(net20025));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20034 (.I(_13695_),
    .Z(net20034));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20139 (.I(_08101_),
    .Z(net20139));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20207 (.I(net20205),
    .Z(net20207));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20023 (.I(_14336_),
    .Z(net20023));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20053 (.I(net20052),
    .Z(net20053));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20169 (.I(net20163),
    .Z(net20169));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20055 (.I(net20052),
    .Z(net20055));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20050 (.I(_11241_),
    .Z(net20050));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20046 (.I(net20045),
    .Z(net20046));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20042 (.I(_12114_),
    .Z(net20042));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20040 (.I(_12184_),
    .Z(net20040));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20041 (.I(net20040),
    .Z(net20041));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20024 (.I(_13739_),
    .Z(net20024));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20036 (.I(_13106_),
    .Z(net20036));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20035 (.I(_13106_),
    .Z(net20035));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20181 (.I(net20180),
    .Z(net20181));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20172 (.I(net20170),
    .Z(net20172));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20171 (.I(net20170),
    .Z(net20171));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20044 (.I(_12042_),
    .Z(net20044));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20043 (.I(_12050_),
    .Z(net20043));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20058 (.I(net20052),
    .Z(net20058));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20039 (.I(_12803_),
    .Z(net20039));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20038 (.I(_12851_),
    .Z(net20038));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20083 (.I(net20082),
    .Z(net20083));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20066 (.I(_10103_),
    .Z(net20066));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20047 (.I(_11352_),
    .Z(net20047));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20057 (.I(net20052),
    .Z(net20057));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20062 (.I(_10444_),
    .Z(net20062));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20164 (.I(net20163),
    .Z(net20164));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20163 (.I(_06815_),
    .Z(net20163));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20045 (.I(_11352_),
    .Z(net20045));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20063 (.I(_10439_),
    .Z(net20063));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20056 (.I(net20052),
    .Z(net20056));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20051 (.I(_11232_),
    .Z(net20051));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20363 (.I(_08040_),
    .Z(net20363));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20166 (.I(net20163),
    .Z(net20166));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20138 (.I(_08109_),
    .Z(net20138));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20077 (.I(_09809_),
    .Z(net20077));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20103 (.I(_09172_),
    .Z(net20103));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20100 (.I(_09224_),
    .Z(net20100));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20052 (.I(_10555_),
    .Z(net20052));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20125 (.I(_08579_),
    .Z(net20125));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20085 (.I(_09757_),
    .Z(net20085));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20143 (.I(_08070_),
    .Z(net20143));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20209 (.I(net20205),
    .Z(net20209));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20135 (.I(_08141_),
    .Z(net20135));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20222 (.I(_01008_),
    .Z(net20222));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20130 (.I(_08244_),
    .Z(net20130));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20065 (.I(_10134_),
    .Z(net20065));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20067 (.I(_10040_),
    .Z(net20067));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20165 (.I(net20163),
    .Z(net20165));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20068 (.I(_09976_),
    .Z(net20068));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20086 (.I(_09757_),
    .Z(net20086));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place20070 (.I(_09912_),
    .Z(net20070));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20162 (.I(_06874_),
    .Z(net20162));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20071 (.I(_09900_),
    .Z(net20071));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20072 (.I(_09885_),
    .Z(net20072));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20161 (.I(_06874_),
    .Z(net20161));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20082 (.I(_09779_),
    .Z(net20082));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20074 (.I(_09831_),
    .Z(net20074));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place20076 (.I(_09809_),
    .Z(net20076));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20079 (.I(_09794_),
    .Z(net20079));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20078 (.I(_09794_),
    .Z(net20078));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20080 (.I(_09782_),
    .Z(net20080));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20081 (.I(_09779_),
    .Z(net20081));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20084 (.I(_09771_),
    .Z(net20084));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20094 (.I(_09320_),
    .Z(net20094));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20145 (.I(net20144),
    .Z(net20145));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20089 (.I(_09456_),
    .Z(net20089));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20126 (.I(_08570_),
    .Z(net20126));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20087 (.I(_09751_),
    .Z(net20087));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20092 (.I(_09379_),
    .Z(net20092));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20088 (.I(_09740_),
    .Z(net20088));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20091 (.I(_09379_),
    .Z(net20091));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20129 (.I(_08257_),
    .Z(net20129));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20090 (.I(_09403_),
    .Z(net20090));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20096 (.I(_09294_),
    .Z(net20096));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20098 (.I(_09266_),
    .Z(net20098));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20095 (.I(_09320_),
    .Z(net20095));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20097 (.I(_09287_),
    .Z(net20097));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20093 (.I(_09320_),
    .Z(net20093));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20099 (.I(_09232_),
    .Z(net20099));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20113 (.I(_08706_),
    .Z(net20113));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20106 (.I(_08894_),
    .Z(net20106));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20105 (.I(_09159_),
    .Z(net20105));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20102 (.I(_09174_),
    .Z(net20102));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20101 (.I(_09178_),
    .Z(net20101));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20111 (.I(_08709_),
    .Z(net20111));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20104 (.I(_09162_),
    .Z(net20104));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20108 (.I(_08753_),
    .Z(net20108));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20116 (.I(_08644_),
    .Z(net20116));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20107 (.I(_08849_),
    .Z(net20107));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20110 (.I(_08726_),
    .Z(net20110));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20109 (.I(_08739_),
    .Z(net20109));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20112 (.I(_08706_),
    .Z(net20112));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20122 (.I(_08612_),
    .Z(net20122));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20117 (.I(_08644_),
    .Z(net20117));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20115 (.I(_08661_),
    .Z(net20115));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20118 (.I(_08634_),
    .Z(net20118));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20119 (.I(_08631_),
    .Z(net20119));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20120 (.I(_08628_),
    .Z(net20120));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20121 (.I(_08612_),
    .Z(net20121));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20123 (.I(_08600_),
    .Z(net20123));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20127 (.I(_08568_),
    .Z(net20127));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20224 (.I(net20222),
    .Z(net20224));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20128 (.I(_08317_),
    .Z(net20128));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20131 (.I(_08193_),
    .Z(net20131));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20133 (.I(_08149_),
    .Z(net20133));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20485 (.I(_09244_),
    .Z(net20485));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20479 (.I(_09278_),
    .Z(net20479));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20132 (.I(_08171_),
    .Z(net20132));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20154 (.I(_15648_[0]),
    .Z(net20154));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20150 (.I(_07990_),
    .Z(net20150));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20134 (.I(_08145_),
    .Z(net20134));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20137 (.I(_08111_),
    .Z(net20137));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20149 (.I(_08012_),
    .Z(net20149));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20140 (.I(_08096_),
    .Z(net20140));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20141 (.I(_08093_),
    .Z(net20141));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20142 (.I(_08087_),
    .Z(net20142));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20146 (.I(_08059_),
    .Z(net20146));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20144 (.I(_08067_),
    .Z(net20144));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20147 (.I(_08054_),
    .Z(net20147));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20168 (.I(net20163),
    .Z(net20168));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20153 (.I(_15651_[0]),
    .Z(net20153));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20148 (.I(_08015_),
    .Z(net20148));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20151 (.I(_07978_),
    .Z(net20151));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20158 (.I(_15641_[0]),
    .Z(net20158));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20481 (.I(_09278_),
    .Z(net20481));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20152 (.I(_15653_[0]),
    .Z(net20152));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20155 (.I(_15643_[0]),
    .Z(net20155));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20475 (.I(_09546_),
    .Z(net20475));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20170 (.I(_06757_),
    .Z(net20170));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20159 (.I(_15569_[0]),
    .Z(net20159));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20160 (.I(_15560_[0]),
    .Z(net20160));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20175 (.I(_06194_),
    .Z(net20175));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20177 (.I(_06019_),
    .Z(net20177));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20193 (.I(_04691_),
    .Z(net20193));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20191 (.I(_04691_),
    .Z(net20191));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20174 (.I(_06194_),
    .Z(net20174));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20176 (.I(_06187_),
    .Z(net20176));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20474 (.I(net20473),
    .Z(net20474));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20214 (.I(_02493_),
    .Z(net20214));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20413 (.I(net20412),
    .Z(net20413));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20182 (.I(_05358_),
    .Z(net20182));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20178 (.I(_06000_),
    .Z(net20178));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20405 (.I(_03848_),
    .Z(net20405));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20206 (.I(net20205),
    .Z(net20206));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20502 (.I(_09155_),
    .Z(net20502));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20473 (.I(_15639_[0]),
    .Z(net20473));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20179 (.I(_05514_),
    .Z(net20179));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20188 (.I(_04739_),
    .Z(net20188));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20184 (.I(_05330_),
    .Z(net20184));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20180 (.I(_05418_),
    .Z(net20180));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20189 (.I(_04739_),
    .Z(net20189));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20491 (.I(_09195_),
    .Z(net20491));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20488 (.I(_09204_),
    .Z(net20488));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20186 (.I(_05280_),
    .Z(net20186));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20550 (.I(net20542),
    .Z(net20550));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20185 (.I(_05297_),
    .Z(net20185));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place20471 (.I(net661),
    .Z(net20471));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20503 (.I(net20502),
    .Z(net20503));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20577 (.I(_07717_),
    .Z(net20577));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20204 (.I(_03257_),
    .Z(net20204));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20187 (.I(_04739_),
    .Z(net20187));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20194 (.I(_04563_),
    .Z(net20194));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20195 (.I(_04544_),
    .Z(net20195));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20199 (.I(_03325_),
    .Z(net20199));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20196 (.I(_04062_),
    .Z(net20196));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20212 (.I(net20211),
    .Z(net20212));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20399 (.I(_05275_),
    .Z(net20399));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place20198 (.I(_03791_),
    .Z(net20198));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20203 (.I(net20202),
    .Z(net20203));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20202 (.I(_03257_),
    .Z(net20202));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20197 (.I(_03827_),
    .Z(net20197));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20201 (.I(_03257_),
    .Z(net20201));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20213 (.I(_02493_),
    .Z(net20213));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20200 (.I(_03257_),
    .Z(net20200));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20211 (.I(_02561_),
    .Z(net20211));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20205 (.I(_03189_),
    .Z(net20205));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20242 (.I(_14485_),
    .Z(net20242));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20227 (.I(_00876_),
    .Z(net20227));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20422 (.I(_01712_),
    .Z(net20422));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20573 (.I(_07717_),
    .Z(net20573));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20220 (.I(_01740_),
    .Z(net20220));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20215 (.I(_02457_),
    .Z(net20215));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20395 (.I(_06142_),
    .Z(net20395));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18425 (.I(_15675_[0]),
    .Z(net18425));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20267 (.I(_12969_),
    .Z(net20267));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20266 (.I(_12969_),
    .Z(net20266));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20265 (.I(net20264),
    .Z(net20265));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20500 (.I(net20499),
    .Z(net20500));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20223 (.I(net20222),
    .Z(net20223));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20499 (.I(_09186_),
    .Z(net20499));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20388 (.I(_15544_[0]),
    .Z(net20388));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20216 (.I(_02456_),
    .Z(net20216));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20372 (.I(_15621_[0]),
    .Z(net20372));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20217 (.I(_02314_),
    .Z(net20217));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20415 (.I(net20412),
    .Z(net20415));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20259 (.I(net20258),
    .Z(net20259));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20343 (.I(_08220_),
    .Z(net20343));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20351 (.I(_08114_),
    .Z(net20351));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20360 (.I(_08044_),
    .Z(net20360));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20228 (.I(_00868_),
    .Z(net20228));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20219 (.I(_01740_),
    .Z(net20219));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20218 (.I(_01740_),
    .Z(net20218));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20374 (.I(_15617_[0]),
    .Z(net20374));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20221 (.I(_01596_),
    .Z(net20221));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20229 (.I(_00849_),
    .Z(net20229));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20248 (.I(_13738_),
    .Z(net20248));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20233 (.I(_15239_),
    .Z(net20233));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20235 (.I(net20234),
    .Z(net20235));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20237 (.I(_15112_),
    .Z(net20237));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20238 (.I(_15088_),
    .Z(net20238));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20230 (.I(_00825_),
    .Z(net20230));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20231 (.I(_15239_),
    .Z(net20231));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20234 (.I(_15120_),
    .Z(net20234));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20240 (.I(_14485_),
    .Z(net20240));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20239 (.I(_14485_),
    .Z(net20239));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20255 (.I(_13663_),
    .Z(net20255));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20244 (.I(_14382_),
    .Z(net20244));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20245 (.I(_14374_),
    .Z(net20245));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20246 (.I(_14357_),
    .Z(net20246));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18423 (.I(_15680_[0]),
    .Z(net18423));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18542 (.I(net18541),
    .Z(net18542));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20593 (.I(_07571_),
    .Z(net20593));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20271 (.I(net20270),
    .Z(net20271));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20247 (.I(_14334_),
    .Z(net20247));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20258 (.I(_13043_),
    .Z(net20258));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20260 (.I(net20258),
    .Z(net20260));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20256 (.I(_13597_),
    .Z(net20256));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20766 (.I(net20757),
    .Z(net20766));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20272 (.I(_12801_),
    .Z(net20272));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20601 (.I(_07571_),
    .Z(net20601));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20572 (.I(_07717_),
    .Z(net20572));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20276 (.I(net20275),
    .Z(net20276));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20362 (.I(_08040_),
    .Z(net20362));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20270 (.I(_12969_),
    .Z(net20270));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20257 (.I(_13043_),
    .Z(net20257));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20264 (.I(_12969_),
    .Z(net20264));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20275 (.I(_12160_),
    .Z(net20275));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18398 (.I(_15899_[0]),
    .Z(net18398));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18391 (.I(_15967_[0]),
    .Z(net18391));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18259 (.I(_13844_),
    .Z(net18259));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20274 (.I(_12160_),
    .Z(net20274));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20311 (.I(_09173_),
    .Z(net20311));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20319 (.I(_08783_),
    .Z(net20319));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20342 (.I(_08245_),
    .Z(net20342));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20278 (.I(_12012_),
    .Z(net20278));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20335 (.I(net20334),
    .Z(net20335));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20349 (.I(_08121_),
    .Z(net20349));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20344 (.I(_08168_),
    .Z(net20344));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20301 (.I(_09290_),
    .Z(net20301));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20334 (.I(_08592_),
    .Z(net20334));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20291 (.I(_09784_),
    .Z(net20291));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20279 (.I(_11209_),
    .Z(net20279));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20409 (.I(net20408),
    .Z(net20409));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20407 (.I(_03263_),
    .Z(net20407));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20394 (.I(_06734_),
    .Z(net20394));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20411 (.I(net20410),
    .Z(net20411));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20381 (.I(_15587_[0]),
    .Z(net20381));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20315 (.I(_09156_),
    .Z(net20315));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18258 (.I(_13851_),
    .Z(net18258));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20292 (.I(_09778_),
    .Z(net20292));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20288 (.I(_09813_),
    .Z(net20288));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20285 (.I(_09878_),
    .Z(net20285));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20283 (.I(_09965_),
    .Z(net20283));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20298 (.I(_09319_),
    .Z(net20298));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20280 (.I(_10443_),
    .Z(net20280));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20281 (.I(_10435_),
    .Z(net20281));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20286 (.I(_09870_),
    .Z(net20286));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20282 (.I(_10380_),
    .Z(net20282));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20289 (.I(_09813_),
    .Z(net20289));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20284 (.I(_09928_),
    .Z(net20284));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18262 (.I(_13836_),
    .Z(net18262));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20313 (.I(net20312),
    .Z(net20313));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20287 (.I(_09855_),
    .Z(net20287));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20290 (.I(_09784_),
    .Z(net20290));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20331 (.I(_08603_),
    .Z(net20331));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20293 (.I(_09768_),
    .Z(net20293));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20296 (.I(_09459_),
    .Z(net20296));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20299 (.I(_09305_),
    .Z(net20299));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20294 (.I(_09738_),
    .Z(net20294));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20295 (.I(_09578_),
    .Z(net20295));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18256 (.I(_13895_),
    .Z(net18256));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18254 (.I(_13903_),
    .Z(net18254));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20307 (.I(_09231_),
    .Z(net20307));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20312 (.I(_09165_),
    .Z(net20312));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20297 (.I(_09387_),
    .Z(net20297));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20300 (.I(_09293_),
    .Z(net20300));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20309 (.I(_09228_),
    .Z(net20309));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20302 (.I(_09261_),
    .Z(net20302));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20303 (.I(_09254_),
    .Z(net20303));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20304 (.I(_09242_),
    .Z(net20304));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20305 (.I(_09239_),
    .Z(net20305));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20306 (.I(_09231_),
    .Z(net20306));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20308 (.I(_09228_),
    .Z(net20308));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20310 (.I(_09219_),
    .Z(net20310));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18253 (.I(_13905_),
    .Z(net18253));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20314 (.I(_09161_),
    .Z(net20314));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20318 (.I(_08904_),
    .Z(net20318));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20316 (.I(_09069_),
    .Z(net20316));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20317 (.I(_09040_),
    .Z(net20317));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20325 (.I(_08660_),
    .Z(net20325));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place18315 (.I(net475),
    .Z(net18315));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20322 (.I(_08687_),
    .Z(net20322));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20321 (.I(_08687_),
    .Z(net20321));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20320 (.I(_08705_),
    .Z(net20320));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20340 (.I(net20339),
    .Z(net20340));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20323 (.I(_08682_),
    .Z(net20323));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20333 (.I(net20332),
    .Z(net20333));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20324 (.I(_08674_),
    .Z(net20324));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20326 (.I(_08633_),
    .Z(net20326));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20361 (.I(_08044_),
    .Z(net20361));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20327 (.I(_08625_),
    .Z(net20327));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20329 (.I(_08622_),
    .Z(net20329));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20328 (.I(_08622_),
    .Z(net20328));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20337 (.I(_08578_),
    .Z(net20337));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20332 (.I(_08599_),
    .Z(net20332));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20330 (.I(_08603_),
    .Z(net20330));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20336 (.I(_08584_),
    .Z(net20336));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20375 (.I(_15614_[0]),
    .Z(net20375));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place18314 (.I(_15738_[0]),
    .Z(net18314));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20338 (.I(_08569_),
    .Z(net20338));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20346 (.I(_08138_),
    .Z(net20346));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20348 (.I(_08121_),
    .Z(net20348));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18313 (.I(_12493_),
    .Z(net18313));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18311 (.I(_12919_),
    .Z(net18311));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20339 (.I(_08566_),
    .Z(net20339));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20341 (.I(_08353_),
    .Z(net20341));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20345 (.I(_08152_),
    .Z(net20345));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20347 (.I(_08121_),
    .Z(net20347));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20358 (.I(net20357),
    .Z(net20358));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20356 (.I(_08058_),
    .Z(net20356));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20353 (.I(_08100_),
    .Z(net20353));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20354 (.I(_08088_),
    .Z(net20354));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20352 (.I(_08100_),
    .Z(net20352));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20357 (.I(_08058_),
    .Z(net20357));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20355 (.I(_08066_),
    .Z(net20355));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20359 (.I(_08050_),
    .Z(net20359));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place18263 (.I(_13832_),
    .Z(net18263));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20369 (.I(_15635_[0]),
    .Z(net20369));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20383 (.I(_15585_[0]),
    .Z(net20383));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20385 (.I(_15580_[0]),
    .Z(net20385));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20364 (.I(_08037_),
    .Z(net20364));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20365 (.I(_08011_),
    .Z(net20365));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20367 (.I(_15657_[0]),
    .Z(net20367));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18308 (.I(_12972_),
    .Z(net18308));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20376 (.I(net20375),
    .Z(net20376));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18205 (.I(_15871_[0]),
    .Z(net18205));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20366 (.I(_07988_),
    .Z(net20366));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20368 (.I(_15655_[0]),
    .Z(net20368));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20370 (.I(_15633_[0]),
    .Z(net20370));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18198 (.I(_15386_),
    .Z(net18198));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18197 (.I(_15386_),
    .Z(net18197));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20386 (.I(_15553_[0]),
    .Z(net20386));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20371 (.I(_15623_[0]),
    .Z(net20371));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20384 (.I(_15583_[0]),
    .Z(net20384));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20373 (.I(_15619_[0]),
    .Z(net20373));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20377 (.I(_15612_[0]),
    .Z(net20377));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20378 (.I(_15603_[0]),
    .Z(net20378));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20379 (.I(_15601_[0]),
    .Z(net20379));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20380 (.I(_15589_[0]),
    .Z(net20380));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20382 (.I(_15587_[0]),
    .Z(net20382));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20393 (.I(_06866_),
    .Z(net20393));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20391 (.I(_06866_),
    .Z(net20391));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20387 (.I(_15546_[0]),
    .Z(net20387));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20587 (.I(_07630_),
    .Z(net20587));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20392 (.I(net20391),
    .Z(net20392));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20410 (.I(_03220_),
    .Z(net20410));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20498 (.I(_09186_),
    .Z(net20498));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20487 (.I(_09215_),
    .Z(net20487));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20401 (.I(_04539_),
    .Z(net20401));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20496 (.I(net20495),
    .Z(net20496));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20406 (.I(_03263_),
    .Z(net20406));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20586 (.I(_07630_),
    .Z(net20586));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20397 (.I(_05386_),
    .Z(net20397));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20396 (.I(_05995_),
    .Z(net20396));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20571 (.I(_07717_),
    .Z(net20571));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20400 (.I(_04690_),
    .Z(net20400));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20398 (.I(_05333_),
    .Z(net20398));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20425 (.I(_01018_),
    .Z(net20425));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20402 (.I(_03999_),
    .Z(net20402));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20403 (.I(net20402),
    .Z(net20403));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20404 (.I(_03852_),
    .Z(net20404));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20570 (.I(_07717_),
    .Z(net20570));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20424 (.I(_01018_),
    .Z(net20424));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20421 (.I(_01739_),
    .Z(net20421));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20417 (.I(_02422_),
    .Z(net20417));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20412 (.I(_02503_),
    .Z(net20412));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20408 (.I(_03220_),
    .Z(net20408));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20414 (.I(net20412),
    .Z(net20414));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20446 (.I(_09875_),
    .Z(net20446));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place20438 (.I(_13636_),
    .Z(net20438));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20419 (.I(_02360_),
    .Z(net20419));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20445 (.I(_11204_),
    .Z(net20445));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20420 (.I(_02356_),
    .Z(net20420));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20497 (.I(_09186_),
    .Z(net20497));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20428 (.I(_15288_),
    .Z(net20428));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20434 (.I(net20433),
    .Z(net20434));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20427 (.I(_15288_),
    .Z(net20427));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20423 (.I(_01638_),
    .Z(net20423));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20510 (.I(_08621_),
    .Z(net20510));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20426 (.I(_00844_),
    .Z(net20426));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place20472 (.I(net663),
    .Z(net20472));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20430 (.I(net20429),
    .Z(net20430));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20429 (.I(_15238_),
    .Z(net20429));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20440 (.I(_12314_),
    .Z(net20440));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20431 (.I(_14517_),
    .Z(net20431));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20433 (.I(_14483_),
    .Z(net20433));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20437 (.I(_14352_),
    .Z(net20437));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20452 (.I(_09838_),
    .Z(net20452));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20551 (.I(net20542),
    .Z(net20551));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20457 (.I(net20455),
    .Z(net20457));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20456 (.I(net20455),
    .Z(net20456));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20470 (.I(_09737_),
    .Z(net20470));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20549 (.I(net20542),
    .Z(net20549));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20447 (.I(net20446),
    .Z(net20447));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20448 (.I(_09854_),
    .Z(net20448));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20443 (.I(_12159_),
    .Z(net20443));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20444 (.I(_11388_),
    .Z(net20444));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20534 (.I(_08027_),
    .Z(net20534));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20564 (.I(_07717_),
    .Z(net20564));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20576 (.I(_07717_),
    .Z(net20576));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20501 (.I(_09186_),
    .Z(net20501));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20458 (.I(net20455),
    .Z(net20458));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20568 (.I(_07717_),
    .Z(net20568));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20569 (.I(net20568),
    .Z(net20569));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20493 (.I(_09186_),
    .Z(net20493));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20492 (.I(_09186_),
    .Z(net20492));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20449 (.I(_09847_),
    .Z(net20449));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20453 (.I(_09838_),
    .Z(net20453));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20553 (.I(net20542),
    .Z(net20553));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20454 (.I(_09827_),
    .Z(net20454));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20455 (.I(_09742_),
    .Z(net20455));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20552 (.I(net20542),
    .Z(net20552));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20567 (.I(_07717_),
    .Z(net20567));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20548 (.I(net20542),
    .Z(net20548));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20563 (.I(net20562),
    .Z(net20563));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20559 (.I(net20558),
    .Z(net20559));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18171 (.I(_01096_),
    .Z(net18171));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20480 (.I(net20479),
    .Z(net20480));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20478 (.I(_09279_),
    .Z(net20478));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20476 (.I(_09343_),
    .Z(net20476));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20477 (.I(_09343_),
    .Z(net20477));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18172 (.I(_01090_),
    .Z(net18172));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18164 (.I(_01194_),
    .Z(net18164));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18086 (.I(_04233_),
    .Z(net18086));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18083 (.I(_04598_),
    .Z(net18083));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18129 (.I(_02722_),
    .Z(net18129));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18118 (.I(_03351_),
    .Z(net18118));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18123 (.I(_03235_),
    .Z(net18123));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18126 (.I(_03235_),
    .Z(net18126));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18110 (.I(_03977_),
    .Z(net18110));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20484 (.I(_09249_),
    .Z(net20484));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20511 (.I(_08621_),
    .Z(net20511));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18081 (.I(_04657_),
    .Z(net18081));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place18080 (.I(_04660_),
    .Z(net18080));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20482 (.I(_09275_),
    .Z(net20482));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18079 (.I(_04663_),
    .Z(net18079));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18077 (.I(_04697_),
    .Z(net18077));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20483 (.I(_09249_),
    .Z(net20483));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20546 (.I(net20542),
    .Z(net20546));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20486 (.I(_09215_),
    .Z(net20486));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20538 (.I(_08006_),
    .Z(net20538));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20489 (.I(_09198_),
    .Z(net20489));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20495 (.I(_09186_),
    .Z(net20495));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20504 (.I(_08688_),
    .Z(net20504));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20494 (.I(_09186_),
    .Z(net20494));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20537 (.I(_08027_),
    .Z(net20537));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20547 (.I(net20542),
    .Z(net20547));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20518 (.I(net20517),
    .Z(net20518));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20505 (.I(net20504),
    .Z(net20505));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20536 (.I(_08027_),
    .Z(net20536));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20506 (.I(_08686_),
    .Z(net20506));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18075 (.I(net18074),
    .Z(net18075));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20535 (.I(net20534),
    .Z(net20535));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20507 (.I(_08654_),
    .Z(net20507));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18070 (.I(_04771_),
    .Z(net18070));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18069 (.I(_04774_),
    .Z(net18069));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18062 (.I(_04789_),
    .Z(net18062));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20610 (.I(net20608),
    .Z(net20610));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20596 (.I(_07571_),
    .Z(net20596));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20595 (.I(net20594),
    .Z(net20595));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20515 (.I(_08587_),
    .Z(net20515));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20508 (.I(_08642_),
    .Z(net20508));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20509 (.I(_08637_),
    .Z(net20509));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20528 (.I(_08048_),
    .Z(net20528));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20512 (.I(_08606_),
    .Z(net20512));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20516 (.I(_08587_),
    .Z(net20516));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20562 (.I(_07727_),
    .Z(net20562));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20527 (.I(_08048_),
    .Z(net20527));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20513 (.I(_08590_),
    .Z(net20513));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20558 (.I(_07727_),
    .Z(net20558));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20514 (.I(_08587_),
    .Z(net20514));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20517 (.I(_08577_),
    .Z(net20517));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20557 (.I(_07727_),
    .Z(net20557));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20544 (.I(net20542),
    .Z(net20544));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20554 (.I(_07976_),
    .Z(net20554));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20543 (.I(net20542),
    .Z(net20543));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20526 (.I(_08056_),
    .Z(net20526));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20524 (.I(_08084_),
    .Z(net20524));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20519 (.I(_08565_),
    .Z(net20519));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20520 (.I(_08201_),
    .Z(net20520));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20531 (.I(_08033_),
    .Z(net20531));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20521 (.I(_08162_),
    .Z(net20521));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20523 (.I(_08084_),
    .Z(net20523));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20529 (.I(_08038_),
    .Z(net20529));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20522 (.I(_08086_),
    .Z(net20522));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20525 (.I(_08056_),
    .Z(net20525));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20530 (.I(_08038_),
    .Z(net20530));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20561 (.I(_07727_),
    .Z(net20561));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20545 (.I(net20542),
    .Z(net20545));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20533 (.I(_08027_),
    .Z(net20533));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20532 (.I(_08027_),
    .Z(net20532));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20540 (.I(_07996_),
    .Z(net20540));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20539 (.I(_08006_),
    .Z(net20539));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20560 (.I(_07727_),
    .Z(net20560));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20541 (.I(_07993_),
    .Z(net20541));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20594 (.I(_07571_),
    .Z(net20594));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20600 (.I(net20599),
    .Z(net20600));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20556 (.I(_07976_),
    .Z(net20556));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20555 (.I(_07976_),
    .Z(net20555));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20599 (.I(_07571_),
    .Z(net20599));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20585 (.I(_07630_),
    .Z(net20585));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20542 (.I(_07984_),
    .Z(net20542));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20565 (.I(_07717_),
    .Z(net20565));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20575 (.I(_07717_),
    .Z(net20575));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20566 (.I(_07717_),
    .Z(net20566));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20584 (.I(_07630_),
    .Z(net20584));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20609 (.I(net20608),
    .Z(net20609));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18065 (.I(_04781_),
    .Z(net18065));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18059 (.I(_04852_),
    .Z(net18059));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18057 (.I(_04902_),
    .Z(net18057));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18068 (.I(_04774_),
    .Z(net18068));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18055 (.I(_04981_),
    .Z(net18055));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18054 (.I(_05324_),
    .Z(net18054));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18048 (.I(_05422_),
    .Z(net18048));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20621 (.I(_15574_[0]),
    .Z(net20621));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20583 (.I(_07630_),
    .Z(net20583));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20582 (.I(_07630_),
    .Z(net20582));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20581 (.I(net20580),
    .Z(net20581));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20579 (.I(_07630_),
    .Z(net20579));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20580 (.I(_07630_),
    .Z(net20580));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20616 (.I(_15608_[0]),
    .Z(net20616));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20673 (.I(net20669),
    .Z(net20673));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20672 (.I(net20669),
    .Z(net20672));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20597 (.I(_07571_),
    .Z(net20597));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20598 (.I(_07571_),
    .Z(net20598));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20636 (.I(_13322_),
    .Z(net20636));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20693 (.I(net20685),
    .Z(net20693));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20608 (.I(_07330_),
    .Z(net20608));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20607 (.I(_07330_),
    .Z(net20607));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20656 (.I(net20654),
    .Z(net20656));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20692 (.I(net20685),
    .Z(net20692));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20604 (.I(_07330_),
    .Z(net20604));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20603 (.I(_07330_),
    .Z(net20603));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20606 (.I(_07330_),
    .Z(net20606));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20605 (.I(_07330_),
    .Z(net20605));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20691 (.I(net20685),
    .Z(net20691));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20690 (.I(net20685),
    .Z(net20690));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20658 (.I(net20654),
    .Z(net20658));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20615 (.I(_15609_[0]),
    .Z(net20615));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20662 (.I(net20659),
    .Z(net20662));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20661 (.I(net20659),
    .Z(net20661));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20660 (.I(net20659),
    .Z(net20660));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20657 (.I(net20654),
    .Z(net20657));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20659 (.I(_09182_),
    .Z(net20659));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20649 (.I(_09762_),
    .Z(net20649));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20633 (.I(_13821_),
    .Z(net20633));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20732 (.I(net20721),
    .Z(net20732));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20625 (.I(_15539_[0]),
    .Z(net20625));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20731 (.I(net20721),
    .Z(net20731));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20735 (.I(net20721),
    .Z(net20735));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20689 (.I(net20685),
    .Z(net20689));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20648 (.I(_09762_),
    .Z(net20648));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20618 (.I(_15594_[0]),
    .Z(net20618));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20635 (.I(net20634),
    .Z(net20635));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18073 (.I(_04747_),
    .Z(net18073));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18045 (.I(_05431_),
    .Z(net18045));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20686 (.I(net20685),
    .Z(net20686));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20626 (.I(_06713_),
    .Z(net20626));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20685 (.I(_07706_),
    .Z(net20685));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20684 (.I(net20683),
    .Z(net20684));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20683 (.I(net20681),
    .Z(net20683));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20682 (.I(net20681),
    .Z(net20682));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20681 (.I(_07706_),
    .Z(net20681));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20671 (.I(net20669),
    .Z(net20671));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18044 (.I(_05434_),
    .Z(net18044));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20670 (.I(net20669),
    .Z(net20670));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20666 (.I(_08575_),
    .Z(net20666));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18043 (.I(_05471_),
    .Z(net18043));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18035 (.I(_06052_),
    .Z(net18035));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18031 (.I(_06200_),
    .Z(net18031));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18030 (.I(_06202_),
    .Z(net18030));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20619 (.I(_15575_[0]),
    .Z(net20619));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20617 (.I(_15607_[0]),
    .Z(net20617));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18022 (.I(_06784_),
    .Z(net18022));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18021 (.I(_06790_),
    .Z(net18021));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20631 (.I(_15286_),
    .Z(net20631));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20627 (.I(_05974_),
    .Z(net20627));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20620 (.I(_15574_[0]),
    .Z(net20620));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20622 (.I(_15573_[0]),
    .Z(net20622));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20680 (.I(net20669),
    .Z(net20680));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20623 (.I(_15541_[0]),
    .Z(net20623));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20624 (.I(_15540_[0]),
    .Z(net20624));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20628 (.I(_05970_),
    .Z(net20628));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20663 (.I(_08934_),
    .Z(net20663));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20630 (.I(_01016_),
    .Z(net20630));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20653 (.I(_09203_),
    .Z(net20653));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20632 (.I(_14515_),
    .Z(net20632));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17897 (.I(_13057_),
    .Z(net17897));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20651 (.I(net20650),
    .Z(net20651));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17894 (.I(_13075_),
    .Z(net17894));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20634 (.I(_13747_),
    .Z(net20634));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20647 (.I(_09762_),
    .Z(net20647));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20644 (.I(_10590_),
    .Z(net20644));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20650 (.I(_09369_),
    .Z(net20650));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20641 (.I(_11441_),
    .Z(net20641));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20637 (.I(_12256_),
    .Z(net20637));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20655 (.I(net20654),
    .Z(net20655));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20638 (.I(_12156_),
    .Z(net20638));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17892 (.I(_13093_),
    .Z(net17892));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17899 (.I(_13046_),
    .Z(net17899));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20643 (.I(_10590_),
    .Z(net20643));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20639 (.I(_12082_),
    .Z(net20639));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17889 (.I(_13183_),
    .Z(net17889));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17887 (.I(_13212_),
    .Z(net17887));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20640 (.I(_12071_),
    .Z(net20640));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20642 (.I(_10641_),
    .Z(net20642));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17901 (.I(_13021_),
    .Z(net17901));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20645 (.I(_10475_),
    .Z(net20645));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17886 (.I(_13370_),
    .Z(net17886));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17882 (.I(_13750_),
    .Z(net17882));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17943 (.I(_11399_),
    .Z(net17943));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20646 (.I(_09762_),
    .Z(net20646));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20654 (.I(_09182_),
    .Z(net20654));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20652 (.I(_09203_),
    .Z(net20652));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17835 (.I(_15295_),
    .Z(net17835));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17841 (.I(_15242_),
    .Z(net17841));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17927 (.I(_11774_),
    .Z(net17927));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17840 (.I(_15242_),
    .Z(net17840));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17839 (.I(_15242_),
    .Z(net17839));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17834 (.I(_15315_),
    .Z(net17834));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20730 (.I(net20721),
    .Z(net20730));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20702 (.I(net20701),
    .Z(net20702));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20734 (.I(net20721),
    .Z(net20734));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20697 (.I(_07697_),
    .Z(net20697));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20668 (.I(_07726_),
    .Z(net20668));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20669 (.I(_07716_),
    .Z(net20669));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20665 (.I(_08626_),
    .Z(net20665));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20664 (.I(_08653_),
    .Z(net20664));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20688 (.I(net20685),
    .Z(net20688));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20701 (.I(net20697),
    .Z(net20701));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17829 (.I(_15350_),
    .Z(net17829));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17742 (.I(_02644_),
    .Z(net17742));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20667 (.I(_08184_),
    .Z(net20667));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17827 (.I(_00906_),
    .Z(net17827));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17752 (.I(_02488_),
    .Z(net17752));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17750 (.I(_02525_),
    .Z(net17750));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17787 (.I(_01667_),
    .Z(net17787));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place17753 (.I(_02482_),
    .Z(net17753));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17795 (.I(_01212_),
    .Z(net17795));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17766 (.I(_01831_),
    .Z(net17766));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17764 (.I(_01880_),
    .Z(net17764));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17779 (.I(_01722_),
    .Z(net17779));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17763 (.I(_02345_),
    .Z(net17763));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17738 (.I(_02777_),
    .Z(net17738));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17728 (.I(_03273_),
    .Z(net17728));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17722 (.I(_03287_),
    .Z(net17722));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20699 (.I(net20697),
    .Z(net20699));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19094 (.I(net19082),
    .Z(net19094));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20698 (.I(net20697),
    .Z(net20698));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20687 (.I(net20685),
    .Z(net20687));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place19093 (.I(net19082),
    .Z(net19093));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20938 (.I(_13649_),
    .Z(net20938));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20759 (.I(net20757),
    .Z(net20759));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20758 (.I(net20757),
    .Z(net20758));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20700 (.I(net20697),
    .Z(net20700));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20756 (.I(_07586_),
    .Z(net20756));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20726 (.I(net20721),
    .Z(net20726));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20725 (.I(net20721),
    .Z(net20725));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20711 (.I(net20708),
    .Z(net20711));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20717 (.I(_07639_),
    .Z(net20717));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20729 (.I(net20721),
    .Z(net20729));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20763 (.I(net20757),
    .Z(net20763));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20755 (.I(net20748),
    .Z(net20755));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20719 (.I(_07639_),
    .Z(net20719));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20706 (.I(_15645_[0]),
    .Z(net20706));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20754 (.I(net20748),
    .Z(net20754));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20727 (.I(net20721),
    .Z(net20727));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20720 (.I(_07639_),
    .Z(net20720));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20705 (.I(_15645_[0]),
    .Z(net20705));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20716 (.I(_07639_),
    .Z(net20716));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17720 (.I(_03305_),
    .Z(net17720));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20724 (.I(net20721),
    .Z(net20724));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20753 (.I(net20748),
    .Z(net20753));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18094 (.I(net18093),
    .Z(net18094));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18093 (.I(_04079_),
    .Z(net18093));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20713 (.I(net20712),
    .Z(net20713));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20709 (.I(net20708),
    .Z(net20709));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20708 (.I(_07654_),
    .Z(net20708));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18019 (.I(_06836_),
    .Z(net18019));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18018 (.I(_06847_),
    .Z(net18018));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18635 (.I(net18634),
    .Z(net18635));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18831 (.I(net18813),
    .Z(net18831));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place20712 (.I(_07647_),
    .Z(net20712));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21070 (.I(net21068),
    .Z(net21070));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20728 (.I(net20721),
    .Z(net20728));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21069 (.I(net21068),
    .Z(net21069));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20932 (.I(_02316_),
    .Z(net20932));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20891 (.I(_12833_),
    .Z(net20891));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21068 (.I(_10378_),
    .Z(net21068));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20722 (.I(net20721),
    .Z(net20722));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20723 (.I(net20722),
    .Z(net20723));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20718 (.I(_07639_),
    .Z(net20718));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21037 (.I(net21036),
    .Z(net21037));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place20721 (.I(_07629_),
    .Z(net20721));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20752 (.I(net20748),
    .Z(net20752));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20740 (.I(_07622_),
    .Z(net20740));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20739 (.I(net20738),
    .Z(net20739));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20738 (.I(_07622_),
    .Z(net20738));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21030 (.I(_11965_),
    .Z(net21030));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20751 (.I(net20750),
    .Z(net20751));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20744 (.I(net20743),
    .Z(net20744));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20743 (.I(net20741),
    .Z(net20743));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20742 (.I(net20741),
    .Z(net20742));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20741 (.I(_15582_[0]),
    .Z(net20741));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20747 (.I(net20746),
    .Z(net20747));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21029 (.I(_11965_),
    .Z(net21029));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20774 (.I(_15616_[0]),
    .Z(net20774));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20773 (.I(_15616_[0]),
    .Z(net20773));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20787 (.I(net20782),
    .Z(net20787));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20955 (.I(_10545_),
    .Z(net20955));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18830 (.I(net18813),
    .Z(net18830));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20780 (.I(net20779),
    .Z(net20780));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20775 (.I(net20774),
    .Z(net20775));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20786 (.I(net20782),
    .Z(net20786));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20771 (.I(_07563_),
    .Z(net20771));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20770 (.I(_07563_),
    .Z(net20770));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20746 (.I(_15577_[0]),
    .Z(net20746));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20745 (.I(_15577_[0]),
    .Z(net20745));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20804 (.I(_01654_),
    .Z(net20804));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20785 (.I(net20782),
    .Z(net20785));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18017 (.I(_06849_),
    .Z(net18017));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20750 (.I(net20748),
    .Z(net20750));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20769 (.I(net20768),
    .Z(net20769));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18193 (.I(net18189),
    .Z(net18193));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18230 (.I(_14531_),
    .Z(net18230));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18203 (.I(net401),
    .Z(net18203));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21075 (.I(_10378_),
    .Z(net21075));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21074 (.I(_10378_),
    .Z(net21074));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21073 (.I(_10378_),
    .Z(net21073));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21072 (.I(_10378_),
    .Z(net21072));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20830 (.I(net20828),
    .Z(net20830));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20792 (.I(net20791),
    .Z(net20792));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20748 (.I(_07586_),
    .Z(net20748));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20749 (.I(net20748),
    .Z(net20749));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18192 (.I(net18189),
    .Z(net18192));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20772 (.I(_07563_),
    .Z(net20772));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20829 (.I(net20828),
    .Z(net20829));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20768 (.I(_07563_),
    .Z(net20768));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20767 (.I(_07563_),
    .Z(net20767));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20757 (.I(_07570_),
    .Z(net20757));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20784 (.I(net20782),
    .Z(net20784));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20861 (.I(net20859),
    .Z(net20861));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20798 (.I(net20794),
    .Z(net20798));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18829 (.I(net18828),
    .Z(net18829));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20828 (.I(_15571_[0]),
    .Z(net20828));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20826 (.I(net20823),
    .Z(net20826));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20776 (.I(_15611_[0]),
    .Z(net20776));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20779 (.I(_07536_),
    .Z(net20779));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20778 (.I(_07536_),
    .Z(net20778));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18202 (.I(net18201),
    .Z(net18202));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20855 (.I(net20848),
    .Z(net20855));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20801 (.I(net20794),
    .Z(net20801));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20800 (.I(net20794),
    .Z(net20800));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20799 (.I(net20794),
    .Z(net20799));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20790 (.I(net20788),
    .Z(net20790));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20854 (.I(net20848),
    .Z(net20854));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20808 (.I(net20807),
    .Z(net20808));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20777 (.I(_07536_),
    .Z(net20777));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18237 (.I(net18236),
    .Z(net18237));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20850 (.I(net20848),
    .Z(net20850));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20841 (.I(net20837),
    .Z(net20841));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20793 (.I(_15543_[0]),
    .Z(net20793));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20783 (.I(net20782),
    .Z(net20783));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20781 (.I(_07513_),
    .Z(net20781));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place20782 (.I(net20781),
    .Z(net20782));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20791 (.I(_15548_[0]),
    .Z(net20791));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20789 (.I(net20788),
    .Z(net20789));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20788 (.I(_07484_),
    .Z(net20788));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20807 (.I(_13072_),
    .Z(net20807));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20797 (.I(net20794),
    .Z(net20797));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20803 (.I(_02374_),
    .Z(net20803));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18828 (.I(net18813),
    .Z(net18828));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18196 (.I(_00581_),
    .Z(net18196));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18195 (.I(_00581_),
    .Z(net18195));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17838 (.I(_15295_),
    .Z(net17838));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20796 (.I(net20794),
    .Z(net20796));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20795 (.I(net20794),
    .Z(net20795));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20853 (.I(net20848),
    .Z(net20853));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place20794 (.I(_07319_),
    .Z(net20794));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17833 (.I(_15322_),
    .Z(net17833));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17826 (.I(_00911_),
    .Z(net17826));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21076 (.I(_10378_),
    .Z(net21076));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20812 (.I(_15606_[0]),
    .Z(net20812));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18191 (.I(net18189),
    .Z(net18191));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20805 (.I(_13820_),
    .Z(net20805));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20825 (.I(net20823),
    .Z(net20825));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20809 (.I(_11964_),
    .Z(net20809));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place18106 (.I(_03982_),
    .Z(net18106));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17712 (.I(_03373_),
    .Z(net17712));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20819 (.I(net20817),
    .Z(net20819));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20816 (.I(net20814),
    .Z(net20816));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20806 (.I(_13072_),
    .Z(net20806));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17715 (.I(net17713),
    .Z(net17715));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17692 (.I(_04177_),
    .Z(net17692));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17688 (.I(_04729_),
    .Z(net17688));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17654 (.I(_06053_),
    .Z(net17654));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17647 (.I(_06116_),
    .Z(net17647));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17640 (.I(_06203_),
    .Z(net17640));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20837 (.I(_07735_),
    .Z(net20837));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17646 (.I(_06123_),
    .Z(net17646));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17652 (.I(_06080_),
    .Z(net17652));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20815 (.I(net20814),
    .Z(net20815));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place20810 (.I(_09734_),
    .Z(net20810));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20840 (.I(net20837),
    .Z(net20840));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20813 (.I(_09153_),
    .Z(net20813));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20814 (.I(_09153_),
    .Z(net20814));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20852 (.I(net20848),
    .Z(net20852));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20818 (.I(net20817),
    .Z(net20818));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20811 (.I(_15606_[0]),
    .Z(net20811));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20817 (.I(_15605_[0]),
    .Z(net20817));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20851 (.I(net20848),
    .Z(net20851));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20839 (.I(net20837),
    .Z(net20839));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17699 (.I(net17698),
    .Z(net17699));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21103 (.I(_10338_),
    .Z(net21103));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17696 (.I(net611),
    .Z(net17696));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20827 (.I(_08564_),
    .Z(net20827));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20821 (.I(net20820),
    .Z(net20821));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20820 (.I(_15572_[0]),
    .Z(net20820));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20822 (.I(_15572_[0]),
    .Z(net20822));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20824 (.I(net20823),
    .Z(net20824));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20823 (.I(_08564_),
    .Z(net20823));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20832 (.I(_15538_[0]),
    .Z(net20832));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18190 (.I(net18189),
    .Z(net18190));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20836 (.I(net20834),
    .Z(net20836));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20831 (.I(net20828),
    .Z(net20831));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21503 (.I(net21501),
    .Z(net21503));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20925 (.I(_06719_),
    .Z(net20925));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20908 (.I(_11189_),
    .Z(net20908));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20881 (.I(net20880),
    .Z(net20881));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20835 (.I(net20834),
    .Z(net20835));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20834 (.I(_15537_[0]),
    .Z(net20834));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20879 (.I(_00811_),
    .Z(net20879));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20833 (.I(net20832),
    .Z(net20833));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20860 (.I(net20859),
    .Z(net20860));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20878 (.I(_00811_),
    .Z(net20878));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17890 (.I(_13101_),
    .Z(net17890));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17705 (.I(net17704),
    .Z(net17705));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17694 (.I(_04053_),
    .Z(net17694));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20877 (.I(_01560_),
    .Z(net20877));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17633 (.I(_06622_),
    .Z(net17633));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17645 (.I(_06176_),
    .Z(net17645));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20875 (.I(_01588_),
    .Z(net20875));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20864 (.I(net20863),
    .Z(net20864));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20838 (.I(net20837),
    .Z(net20838));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20856 (.I(_07619_),
    .Z(net20856));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20842 (.I(_07704_),
    .Z(net20842));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place20848 (.I(_07637_),
    .Z(net20848));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20843 (.I(_07695_),
    .Z(net20843));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21099 (.I(_10345_),
    .Z(net21099));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17638 (.I(_06224_),
    .Z(net17638));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17537 (.I(_13762_),
    .Z(net17537));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20844 (.I(_07679_),
    .Z(net20844));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20931 (.I(_03037_),
    .Z(net20931));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17541 (.I(_13210_),
    .Z(net17541));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20858 (.I(_00403_),
    .Z(net20858));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20845 (.I(_00394_),
    .Z(net20845));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20847 (.I(_07660_),
    .Z(net20847));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20846 (.I(_07666_),
    .Z(net20846));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20849 (.I(net20848),
    .Z(net20849));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21071 (.I(_10378_),
    .Z(net21071));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20857 (.I(_00404_),
    .Z(net20857));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20907 (.I(_11210_),
    .Z(net20907));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20862 (.I(_07560_),
    .Z(net20862));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20900 (.I(_12000_),
    .Z(net20900));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20899 (.I(_12024_),
    .Z(net20899));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20910 (.I(_11156_),
    .Z(net20910));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20897 (.I(_12080_),
    .Z(net20897));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20870 (.I(_02320_),
    .Z(net20870));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20866 (.I(_04546_),
    .Z(net20866));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20863 (.I(_07534_),
    .Z(net20863));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20887 (.I(_12889_),
    .Z(net20887));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17878 (.I(_13786_),
    .Z(net17878));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17888 (.I(_13187_),
    .Z(net17888));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place20859 (.I(_07578_),
    .Z(net20859));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place17698 (.I(_03974_),
    .Z(net17698));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21522 (.I(net21521),
    .Z(net21522));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21521 (.I(net21520),
    .Z(net21521));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20949 (.I(_11342_),
    .Z(net20949));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21502 (.I(net21501),
    .Z(net21502));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20873 (.I(_02281_),
    .Z(net20873));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17865 (.I(_14463_),
    .Z(net17865));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place20880 (.I(_00807_),
    .Z(net20880));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20865 (.I(_05281_),
    .Z(net20865));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20930 (.I(_03793_),
    .Z(net20930));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20872 (.I(_02281_),
    .Z(net20872));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20869 (.I(_02325_),
    .Z(net20869));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20867 (.I(_03022_),
    .Z(net20867));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20868 (.I(_03018_),
    .Z(net20868));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20871 (.I(_02285_),
    .Z(net20871));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20915 (.I(_10389_),
    .Z(net20915));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21514 (.I(_07705_),
    .Z(net21514));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21520 (.I(net21518),
    .Z(net21520));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20876 (.I(_01578_),
    .Z(net20876));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20895 (.I(_12770_),
    .Z(net20895));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20874 (.I(_01598_),
    .Z(net20874));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21098 (.I(_10357_),
    .Z(net21098));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20884 (.I(_14317_),
    .Z(net20884));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20890 (.I(_12867_),
    .Z(net20890));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place21097 (.I(_10360_),
    .Z(net21097));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20882 (.I(_15062_),
    .Z(net20882));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21519 (.I(net21518),
    .Z(net21519));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21517 (.I(net21515),
    .Z(net21517));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20885 (.I(_13587_),
    .Z(net20885));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20883 (.I(_14358_),
    .Z(net20883));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20892 (.I(_12809_),
    .Z(net20892));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20886 (.I(_13583_),
    .Z(net20886));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20888 (.I(_12885_),
    .Z(net20888));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20889 (.I(_12876_),
    .Z(net20889));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20901 (.I(_11973_),
    .Z(net20901));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20893 (.I(_12777_),
    .Z(net20893));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20894 (.I(_12774_),
    .Z(net20894));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20896 (.I(_12765_),
    .Z(net20896));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place20904 (.I(_11963_),
    .Z(net20904));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20898 (.I(_12076_),
    .Z(net20898));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20905 (.I(net20904),
    .Z(net20905));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21119 (.I(_07607_),
    .Z(net21119));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21516 (.I(net21515),
    .Z(net21516));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20902 (.I(_11969_),
    .Z(net20902));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20903 (.I(_11963_),
    .Z(net20903));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20906 (.I(_11215_),
    .Z(net20906));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20923 (.I(_07541_),
    .Z(net20923));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20928 (.I(_05266_),
    .Z(net20928));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20924 (.I(_06736_),
    .Z(net20924));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20922 (.I(_07559_),
    .Z(net20922));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20909 (.I(_11161_),
    .Z(net20909));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20920 (.I(net20919),
    .Z(net20920));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20911 (.I(_11152_),
    .Z(net20911));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20917 (.I(_10362_),
    .Z(net20917));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20912 (.I(_10515_),
    .Z(net20912));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20914 (.I(_10427_),
    .Z(net20914));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place20916 (.I(_10366_),
    .Z(net20916));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21530 (.I(_07276_),
    .Z(net21530));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20929 (.I(_04541_),
    .Z(net20929));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place20919 (.I(_10347_),
    .Z(net20919));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place20918 (.I(_10354_),
    .Z(net20918));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20921 (.I(_10342_),
    .Z(net20921));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20926 (.I(_06017_),
    .Z(net20926));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20927 (.I(_05277_),
    .Z(net20927));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17514 (.I(_15221_),
    .Z(net17514));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17511 (.I(_15227_),
    .Z(net17511));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21128 (.I(_07538_),
    .Z(net21128));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21425 (.I(net21424),
    .Z(net21425));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17507 (.I(_15310_),
    .Z(net17507));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21524 (.I(net21518),
    .Z(net21524));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20933 (.I(_01593_),
    .Z(net20933));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21523 (.I(net21518),
    .Z(net21523));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place21501 (.I(net21490),
    .Z(net21501));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21500 (.I(net21490),
    .Z(net21500));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21275 (.I(\sa31_sub[7] ),
    .Z(net21275));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21529 (.I(net21526),
    .Z(net21529));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21499 (.I(net21493),
    .Z(net21499));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20934 (.I(_01573_),
    .Z(net20934));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20937 (.I(_13652_),
    .Z(net20937));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17504 (.I(_00598_),
    .Z(net17504));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17499 (.I(_01029_),
    .Z(net17499));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20935 (.I(_15110_),
    .Z(net20935));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21409 (.I(\sa11_sr[1] ),
    .Z(net21409));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17498 (.I(_01041_),
    .Z(net17498));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20936 (.I(_14354_),
    .Z(net20936));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21527 (.I(net21526),
    .Z(net21527));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21526 (.I(_07276_),
    .Z(net21526));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21424 (.I(net21423),
    .Z(net21424));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21498 (.I(net21493),
    .Z(net21498));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21497 (.I(net21493),
    .Z(net21497));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20940 (.I(_12958_),
    .Z(net20940));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20939 (.I(_13007_),
    .Z(net20939));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20941 (.I(_12896_),
    .Z(net20941));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20943 (.I(_12840_),
    .Z(net20943));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17510 (.I(_15254_),
    .Z(net17510));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20944 (.I(_12831_),
    .Z(net20944));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20945 (.I(_12823_),
    .Z(net20945));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20946 (.I(_12151_),
    .Z(net20946));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20947 (.I(_12022_),
    .Z(net20947));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20964 (.I(_05261_),
    .Z(net20964));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20948 (.I(_11382_),
    .Z(net20948));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20951 (.I(_11304_),
    .Z(net20951));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21496 (.I(net21493),
    .Z(net21496));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20970 (.I(_01557_),
    .Z(net20970));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20950 (.I(_11339_),
    .Z(net20950));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20952 (.I(_11213_),
    .Z(net20952));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21495 (.I(net21493),
    .Z(net21495));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20953 (.I(_11206_),
    .Z(net20953));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20954 (.I(_11187_),
    .Z(net20954));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21542 (.I(net129),
    .Z(net21542));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21538 (.I(net21533),
    .Z(net21538));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20956 (.I(_10419_),
    .Z(net20956));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21494 (.I(net21493),
    .Z(net21494));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20957 (.I(_10416_),
    .Z(net20957));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20958 (.I(_10415_),
    .Z(net20958));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20959 (.I(_10395_),
    .Z(net20959));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20960 (.I(_07699_),
    .Z(net20960));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20962 (.I(_07682_),
    .Z(net20962));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20961 (.I(_07691_),
    .Z(net20961));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17495 (.I(net438),
    .Z(net17495));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21518 (.I(_07276_),
    .Z(net21518));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17494 (.I(_01087_),
    .Z(net17494));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21515 (.I(_07535_),
    .Z(net21515));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17480 (.I(_01720_),
    .Z(net17480));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17478 (.I(_01730_),
    .Z(net17478));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17486 (.I(_01325_),
    .Z(net17486));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17466 (.I(_01841_),
    .Z(net17466));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17442 (.I(_02779_),
    .Z(net17442));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21051 (.I(_10542_),
    .Z(net21051));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20965 (.I(_04530_),
    .Z(net20965));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20995 (.I(_12864_),
    .Z(net20995));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20963 (.I(_05329_),
    .Z(net20963));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20969 (.I(_01557_),
    .Z(net20969));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21525 (.I(_07276_),
    .Z(net21525));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21026 (.I(_11980_),
    .Z(net21026));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20966 (.I(_03773_),
    .Z(net20966));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21528 (.I(net21526),
    .Z(net21528));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21414 (.I(\sa10_sr[7] ),
    .Z(net21414));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20968 (.I(_02278_),
    .Z(net20968));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20973 (.I(_00826_),
    .Z(net20973));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20967 (.I(_03015_),
    .Z(net20967));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20971 (.I(_00918_),
    .Z(net20971));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21015 (.I(_12065_),
    .Z(net21015));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21306 (.I(\sa30_sr[3] ),
    .Z(net21306));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21012 (.I(_12761_),
    .Z(net21012));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20987 (.I(_13580_),
    .Z(net20987));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21021 (.I(_12006_),
    .Z(net21021));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20972 (.I(_00890_),
    .Z(net20972));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20976 (.I(_15064_),
    .Z(net20976));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20974 (.I(_00804_),
    .Z(net20974));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_35_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21017 (.I(_12025_),
    .Z(net21017));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20999 (.I(_12834_),
    .Z(net20999));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20975 (.I(_15075_),
    .Z(net20975));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20981 (.I(_14314_),
    .Z(net20981));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20977 (.I(_15059_),
    .Z(net20977));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20978 (.I(_14410_),
    .Z(net20978));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20997 (.I(_12839_),
    .Z(net20997));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20984 (.I(_13650_),
    .Z(net20984));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20979 (.I(_14400_),
    .Z(net20979));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21001 (.I(_12815_),
    .Z(net21001));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20980 (.I(_14335_),
    .Z(net20980));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21341 (.I(net21340),
    .Z(net21341));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20982 (.I(_13689_),
    .Z(net20982));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20983 (.I(_13653_),
    .Z(net20983));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21305 (.I(\sa30_sr[3] ),
    .Z(net21305));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20985 (.I(_13648_),
    .Z(net20985));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20986 (.I(_13598_),
    .Z(net20986));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20988 (.I(_13068_),
    .Z(net20988));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20989 (.I(_12955_),
    .Z(net20989));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20990 (.I(_12928_),
    .Z(net20990));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20991 (.I(_12882_),
    .Z(net20991));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20992 (.I(_12870_),
    .Z(net20992));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20993 (.I(_12868_),
    .Z(net20993));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21000 (.I(_12832_),
    .Z(net21000));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20994 (.I(_12864_),
    .Z(net20994));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20998 (.I(_12839_),
    .Z(net20998));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20996 (.I(_12841_),
    .Z(net20996));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21294 (.I(\sa30_sub[2] ),
    .Z(net21294));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21413 (.I(\sa10_sr[7] ),
    .Z(net21413));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21005 (.I(_12783_),
    .Z(net21005));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21003 (.I(_12790_),
    .Z(net21003));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21007 (.I(net21006),
    .Z(net21007));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21002 (.I(_12811_),
    .Z(net21002));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21004 (.I(_12783_),
    .Z(net21004));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place21006 (.I(_12780_),
    .Z(net21006));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21009 (.I(_12766_),
    .Z(net21009));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_30_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21008 (.I(_12768_),
    .Z(net21008));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21014 (.I(_12066_),
    .Z(net21014));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21543 (.I(net21542),
    .Z(net21543));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21010 (.I(_12762_),
    .Z(net21010));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21011 (.I(_12761_),
    .Z(net21011));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21013 (.I(_12148_),
    .Z(net21013));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21458 (.I(\sa01_sr[7] ),
    .Z(net21458));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21439 (.I(net21438),
    .Z(net21439));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21323 (.I(\sa21_sub[3] ),
    .Z(net21323));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21018 (.I(_12023_),
    .Z(net21018));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21016 (.I(_12032_),
    .Z(net21016));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21036 (.I(_11223_),
    .Z(net21036));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21019 (.I(_12021_),
    .Z(net21019));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21050 (.I(_10582_),
    .Z(net21050));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21042 (.I(_11190_),
    .Z(net21042));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place21060 (.I(_10396_),
    .Z(net21060));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21020 (.I(_12006_),
    .Z(net21020));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21022 (.I(_12002_),
    .Z(net21022));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21023 (.I(_11992_),
    .Z(net21023));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21025 (.I(_11980_),
    .Z(net21025));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21024 (.I(_11981_),
    .Z(net21024));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21027 (.I(_11978_),
    .Z(net21027));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21028 (.I(_11966_),
    .Z(net21028));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21031 (.I(_11960_),
    .Z(net21031));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21049 (.I(_11147_),
    .Z(net21049));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21032 (.I(_11959_),
    .Z(net21032));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21033 (.I(_11266_),
    .Z(net21033));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21040 (.I(_11212_),
    .Z(net21040));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21034 (.I(_11258_),
    .Z(net21034));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21039 (.I(_11214_),
    .Z(net21039));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21038 (.I(_11216_),
    .Z(net21038));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21035 (.I(_11250_),
    .Z(net21035));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21043 (.I(_11166_),
    .Z(net21043));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21041 (.I(_11194_),
    .Z(net21041));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21067 (.I(_10378_),
    .Z(net21067));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place21061 (.I(_10394_),
    .Z(net21061));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21044 (.I(_11165_),
    .Z(net21044));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21308 (.I(net21307),
    .Z(net21308));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21456 (.I(\sa02_sr[0] ),
    .Z(net21456));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place21045 (.I(_11158_),
    .Z(net21045));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21046 (.I(_11157_),
    .Z(net21046));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21047 (.I(_11149_),
    .Z(net21047));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21048 (.I(_11148_),
    .Z(net21048));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21488 (.I(net21482),
    .Z(net21488));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21056 (.I(net21055),
    .Z(net21056));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21065 (.I(net21064),
    .Z(net21065));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21052 (.I(_10512_),
    .Z(net21052));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17437 (.I(_03148_),
    .Z(net17437));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17462 (.I(_01917_),
    .Z(net17462));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21053 (.I(_10458_),
    .Z(net21053));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21054 (.I(_10450_),
    .Z(net21054));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21055 (.I(_10425_),
    .Z(net21055));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21057 (.I(_10420_),
    .Z(net21057));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21058 (.I(_10417_),
    .Z(net21058));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21313 (.I(\sa30_sr[0] ),
    .Z(net21313));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21064 (.I(_10378_),
    .Z(net21064));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21059 (.I(_10414_),
    .Z(net21059));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21063 (.I(_10382_),
    .Z(net21063));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place21062 (.I(_10391_),
    .Z(net21062));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21066 (.I(_10378_),
    .Z(net21066));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21309 (.I(\sa30_sr[2] ),
    .Z(net21309));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21487 (.I(net21486),
    .Z(net21487));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17452 (.I(_02598_),
    .Z(net17452));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17651 (.I(net490),
    .Z(net17651));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17425 (.I(_03249_),
    .Z(net17425));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21105 (.I(_07908_),
    .Z(net21105));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21100 (.I(_10343_),
    .Z(net21100));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21123 (.I(_07562_),
    .Z(net21123));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17641 (.I(_06203_),
    .Z(net17641));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17639 (.I(_06210_),
    .Z(net17639));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17636 (.I(_06224_),
    .Z(net17636));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17426 (.I(_03245_),
    .Z(net17426));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17634 (.I(_06455_),
    .Z(net17634));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer39 (.I(net19205),
    .Z(net426));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17632 (.I(_06818_),
    .Z(net17632));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17566 (.I(_11708_),
    .Z(net17566));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17562 (.I(_12177_),
    .Z(net17562));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17447 (.I(_02700_),
    .Z(net17447));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17438 (.I(_03148_),
    .Z(net17438));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17435 (.I(net17433),
    .Z(net17435));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17563 (.I(_12177_),
    .Z(net17563));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17444 (.I(_02767_),
    .Z(net17444));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17557 (.I(_12264_),
    .Z(net17557));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17615 (.I(_07018_),
    .Z(net17615));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17440 (.I(_03086_),
    .Z(net17440));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17439 (.I(_03086_),
    .Z(net17439));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17569 (.I(_11532_),
    .Z(net17569));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17455 (.I(_02536_),
    .Z(net17455));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17553 (.I(_12279_),
    .Z(net17553));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17474 (.I(_01750_),
    .Z(net17474));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17477 (.I(_01744_),
    .Z(net17477));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17458 (.I(_02037_),
    .Z(net17458));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17558 (.I(_12264_),
    .Z(net17558));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17551 (.I(_12452_),
    .Z(net17551));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17481 (.I(_01718_),
    .Z(net17481));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17476 (.I(_01744_),
    .Z(net17476));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17631 (.I(_06818_),
    .Z(net17631));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17554 (.I(_12279_),
    .Z(net17554));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17556 (.I(_12276_),
    .Z(net17556));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17550 (.I(_12990_),
    .Z(net17550));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17549 (.I(_12998_),
    .Z(net17549));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21112 (.I(_07689_),
    .Z(net21112));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21104 (.I(_07913_),
    .Z(net21104));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21101 (.I(_10339_),
    .Z(net21101));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21102 (.I(_10338_),
    .Z(net21102));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17427 (.I(_03245_),
    .Z(net17427));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21111 (.I(_07692_),
    .Z(net21111));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21106 (.I(_07874_),
    .Z(net21106));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21107 (.I(_07869_),
    .Z(net21107));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21108 (.I(_07828_),
    .Z(net21108));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21109 (.I(_07782_),
    .Z(net21109));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21110 (.I(_07696_),
    .Z(net21110));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17420 (.I(_03276_),
    .Z(net17420));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17414 (.I(_03385_),
    .Z(net17414));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21120 (.I(_07604_),
    .Z(net21120));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21116 (.I(_07621_),
    .Z(net21116));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21121 (.I(_07599_),
    .Z(net21121));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21113 (.I(_07675_),
    .Z(net21113));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21114 (.I(_07672_),
    .Z(net21114));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21115 (.I(_07624_),
    .Z(net21115));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21117 (.I(_07616_),
    .Z(net21117));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21118 (.I(_07615_),
    .Z(net21118));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21131 (.I(_07464_),
    .Z(net21131));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21272 (.I(\sa32_sub[0] ),
    .Z(net21272));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17419 (.I(_03288_),
    .Z(net17419));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21122 (.I(_07565_),
    .Z(net21122));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21124 (.I(_07556_),
    .Z(net21124));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21249 (.I(\u0.subword[17] ),
    .Z(net21249));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21244 (.I(\u0.subword[9] ),
    .Z(net21244));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21138 (.I(\u0.tmp_w[3] ),
    .Z(net21138));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21126 (.I(_07548_),
    .Z(net21126));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21266 (.I(\sa32_sub[3] ),
    .Z(net21266));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21125 (.I(_07555_),
    .Z(net21125));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21129 (.I(_07531_),
    .Z(net21129));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place21535 (.I(net21533),
    .Z(net21535));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21130 (.I(_07491_),
    .Z(net21130));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21127 (.I(_07539_),
    .Z(net21127));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21534 (.I(net21533),
    .Z(net21534));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21532 (.I(net21531),
    .Z(net21532));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21133 (.I(_07448_),
    .Z(net21133));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21132 (.I(_07463_),
    .Z(net21132));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21531 (.I(net129),
    .Z(net21531));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21135 (.I(_07243_),
    .Z(net21135));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21136 (.I(\u0.tmp_w[9] ),
    .Z(net21136));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21137 (.I(\u0.tmp_w[8] ),
    .Z(net21137));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21139 (.I(\u0.tmp_w[2] ),
    .Z(net21139));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21140 (.I(\u0.tmp_w[29] ),
    .Z(net21140));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21165 (.I(\u0.w[2][28] ),
    .Z(net21165));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21141 (.I(\u0.tmp_w[28] ),
    .Z(net21141));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21149 (.I(\u0.tmp_w[18] ),
    .Z(net21149));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21142 (.I(\u0.tmp_w[27] ),
    .Z(net21142));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21143 (.I(\u0.tmp_w[26] ),
    .Z(net21143));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21144 (.I(\u0.tmp_w[25] ),
    .Z(net21144));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21145 (.I(\u0.tmp_w[24] ),
    .Z(net21145));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21146 (.I(\u0.tmp_w[20] ),
    .Z(net21146));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21147 (.I(\u0.tmp_w[1] ),
    .Z(net21147));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21179 (.I(\u0.w[2][11] ),
    .Z(net21179));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21148 (.I(\u0.tmp_w[19] ),
    .Z(net21148));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21150 (.I(\u0.tmp_w[17] ),
    .Z(net21150));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21151 (.I(\u0.tmp_w[16] ),
    .Z(net21151));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21152 (.I(\u0.tmp_w[12] ),
    .Z(net21152));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21153 (.I(\u0.tmp_w[11] ),
    .Z(net21153));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21154 (.I(\u0.tmp_w[10] ),
    .Z(net21154));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21155 (.I(\u0.tmp_w[0] ),
    .Z(net21155));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21156 (.I(\u0.w[2][9] ),
    .Z(net21156));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21157 (.I(\u0.w[2][8] ),
    .Z(net21157));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21158 (.I(\u0.w[2][5] ),
    .Z(net21158));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21159 (.I(\u0.w[2][4] ),
    .Z(net21159));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21160 (.I(\u0.w[2][3] ),
    .Z(net21160));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21161 (.I(\u0.w[2][31] ),
    .Z(net21161));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21162 (.I(\u0.w[2][30] ),
    .Z(net21162));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21163 (.I(\u0.w[2][2] ),
    .Z(net21163));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21164 (.I(\u0.w[2][29] ),
    .Z(net21164));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21166 (.I(\u0.w[2][27] ),
    .Z(net21166));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21167 (.I(\u0.w[2][26] ),
    .Z(net21167));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21168 (.I(net665),
    .Z(net21168));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21169 (.I(net684),
    .Z(net21169));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21170 (.I(\u0.w[2][21] ),
    .Z(net21170));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21171 (.I(\u0.w[2][20] ),
    .Z(net21171));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21172 (.I(\u0.w[2][1] ),
    .Z(net21172));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21173 (.I(\u0.w[2][19] ),
    .Z(net21173));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21174 (.I(\u0.w[2][18] ),
    .Z(net21174));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21175 (.I(\u0.w[2][17] ),
    .Z(net21175));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21176 (.I(\u0.w[2][16] ),
    .Z(net21176));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21260 (.I(\sa32_sub[7] ),
    .Z(net21260));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21177 (.I(\u0.w[2][13] ),
    .Z(net21177));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21178 (.I(\u0.w[2][12] ),
    .Z(net21178));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21180 (.I(\u0.w[2][10] ),
    .Z(net21180));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21181 (.I(\u0.w[2][0] ),
    .Z(net21181));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21182 (.I(\u0.w[1][9] ),
    .Z(net21182));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21183 (.I(\u0.w[1][8] ),
    .Z(net21183));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21184 (.I(\u0.w[1][7] ),
    .Z(net21184));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21185 (.I(\u0.w[1][6] ),
    .Z(net21185));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21186 (.I(\u0.w[1][5] ),
    .Z(net21186));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21187 (.I(\u0.w[1][4] ),
    .Z(net21187));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21188 (.I(\u0.w[1][3] ),
    .Z(net21188));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21189 (.I(\u0.w[1][2] ),
    .Z(net21189));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21190 (.I(\u0.w[1][29] ),
    .Z(net21190));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21191 (.I(\u0.w[1][28] ),
    .Z(net21191));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21227 (.I(\u0.w[0][19] ),
    .Z(net21227));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21192 (.I(\u0.w[1][27] ),
    .Z(net21192));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21193 (.I(\u0.w[1][26] ),
    .Z(net21193));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21194 (.I(\u0.w[1][25] ),
    .Z(net21194));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21195 (.I(\u0.w[1][24] ),
    .Z(net21195));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21196 (.I(\u0.w[1][22] ),
    .Z(net21196));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21197 (.I(\u0.w[1][21] ),
    .Z(net21197));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21198 (.I(\u0.w[1][20] ),
    .Z(net21198));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21199 (.I(\u0.w[1][1] ),
    .Z(net21199));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21200 (.I(\u0.w[1][19] ),
    .Z(net21200));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21201 (.I(\u0.w[1][18] ),
    .Z(net21201));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21202 (.I(\u0.w[1][17] ),
    .Z(net21202));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21203 (.I(\u0.w[1][16] ),
    .Z(net21203));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21211 (.I(net21210),
    .Z(net21211));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21204 (.I(\u0.w[1][13] ),
    .Z(net21204));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21213 (.I(\u0.w[0][4] ),
    .Z(net21213));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21205 (.I(\u0.w[1][12] ),
    .Z(net21205));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21206 (.I(\u0.w[1][11] ),
    .Z(net21206));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21207 (.I(\u0.w[1][10] ),
    .Z(net21207));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21208 (.I(\u0.w[1][0] ),
    .Z(net21208));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21209 (.I(\u0.w[0][9] ),
    .Z(net21209));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21210 (.I(\u0.w[0][8] ),
    .Z(net21210));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21212 (.I(\u0.w[0][5] ),
    .Z(net21212));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21264 (.I(\sa32_sub[4] ),
    .Z(net21264));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21214 (.I(\u0.w[0][3] ),
    .Z(net21214));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21215 (.I(\u0.w[0][31] ),
    .Z(net21215));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21216 (.I(\u0.w[0][30] ),
    .Z(net21216));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21217 (.I(\u0.w[0][2] ),
    .Z(net21217));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21218 (.I(\u0.w[0][29] ),
    .Z(net21218));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21219 (.I(\u0.w[0][28] ),
    .Z(net21219));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21220 (.I(\u0.w[0][27] ),
    .Z(net21220));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21221 (.I(\u0.w[0][26] ),
    .Z(net21221));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21222 (.I(\u0.w[0][25] ),
    .Z(net21222));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21223 (.I(\u0.w[0][24] ),
    .Z(net21223));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21224 (.I(\u0.w[0][21] ),
    .Z(net21224));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21225 (.I(\u0.w[0][20] ),
    .Z(net21225));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21533 (.I(net21531),
    .Z(net21533));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21226 (.I(\u0.w[0][1] ),
    .Z(net21226));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21228 (.I(\u0.w[0][18] ),
    .Z(net21228));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21229 (.I(\u0.w[0][17] ),
    .Z(net21229));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21230 (.I(\u0.w[0][16] ),
    .Z(net21230));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21231 (.I(\u0.w[0][14] ),
    .Z(net21231));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21232 (.I(\u0.w[0][13] ),
    .Z(net21232));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21233 (.I(\u0.w[0][12] ),
    .Z(net21233));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21234 (.I(\u0.w[0][11] ),
    .Z(net21234));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21235 (.I(\u0.w[0][10] ),
    .Z(net21235));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21236 (.I(\u0.w[0][0] ),
    .Z(net21236));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21237 (.I(\u0.subword[3] ),
    .Z(net21237));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21238 (.I(\u0.subword[2] ),
    .Z(net21238));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21293 (.I(\sa30_sub[2] ),
    .Z(net21293));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21404 (.I(\sa11_sr[6] ),
    .Z(net21404));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21239 (.I(\u0.subword[1] ),
    .Z(net21239));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21240 (.I(\u0.subword[0] ),
    .Z(net21240));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21241 (.I(\u0.subword[12] ),
    .Z(net21241));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21242 (.I(\u0.subword[11] ),
    .Z(net21242));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21267 (.I(\sa32_sub[2] ),
    .Z(net21267));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21243 (.I(\u0.subword[10] ),
    .Z(net21243));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21245 (.I(\u0.subword[8] ),
    .Z(net21245));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21246 (.I(\u0.subword[21] ),
    .Z(net21246));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21247 (.I(\u0.subword[20] ),
    .Z(net21247));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21248 (.I(\u0.subword[19] ),
    .Z(net21248));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21259 (.I(\sa32_sub[7] ),
    .Z(net21259));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21250 (.I(\u0.subword[16] ),
    .Z(net21250));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21251 (.I(\u0.subword[27] ),
    .Z(net21251));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21252 (.I(\u0.subword[26] ),
    .Z(net21252));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21253 (.I(\u0.subword[25] ),
    .Z(net21253));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17410 (.I(_03714_),
    .Z(net17410));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21254 (.I(\u0.subword[24] ),
    .Z(net21254));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21255 (.I(\u0.r0.out[26] ),
    .Z(net21255));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21256 (.I(\u0.r0.out[25] ),
    .Z(net21256));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21257 (.I(\u0.r0.out[24] ),
    .Z(net21257));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17408 (.I(_03882_),
    .Z(net17408));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21258 (.I(\sa32_sub[7] ),
    .Z(net21258));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21261 (.I(\sa32_sub[6] ),
    .Z(net21261));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21262 (.I(\sa32_sub[5] ),
    .Z(net21262));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17403 (.I(_04147_),
    .Z(net17403));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17429 (.I(net17428),
    .Z(net17429));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17409 (.I(net17408),
    .Z(net17409));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17394 (.I(_04342_),
    .Z(net17394));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17336 (.I(_12227_),
    .Z(net17336));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17337 (.I(_12227_),
    .Z(net17337));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17334 (.I(_12237_),
    .Z(net17334));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17333 (.I(_12237_),
    .Z(net17333));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17328 (.I(_12290_),
    .Z(net17328));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17327 (.I(_12295_),
    .Z(net17327));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17325 (.I(_12354_),
    .Z(net17325));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_25_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17357 (.I(_11297_),
    .Z(net17357));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17310 (.I(_14817_),
    .Z(net17310));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17302 (.I(_15246_),
    .Z(net17302));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_28_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17298 (.I(_15290_),
    .Z(net17298));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17295 (.I(_15345_),
    .Z(net17295));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21322 (.I(\sa21_sub[3] ),
    .Z(net21322));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17506 (.I(_15375_),
    .Z(net17506));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21311 (.I(\sa30_sr[1] ),
    .Z(net21311));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21286 (.I(\sa30_sub[7] ),
    .Z(net21286));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21276 (.I(\sa31_sub[6] ),
    .Z(net21276));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21287 (.I(\sa30_sub[7] ),
    .Z(net21287));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21263 (.I(\sa32_sub[4] ),
    .Z(net21263));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21270 (.I(net21269),
    .Z(net21270));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21265 (.I(\sa32_sub[3] ),
    .Z(net21265));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21268 (.I(\sa32_sub[2] ),
    .Z(net21268));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21269 (.I(\sa32_sub[1] ),
    .Z(net21269));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21280 (.I(\sa31_sub[3] ),
    .Z(net21280));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21271 (.I(\sa32_sub[0] ),
    .Z(net21271));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21274 (.I(\sa31_sub[7] ),
    .Z(net21274));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21273 (.I(\sa31_sub[7] ),
    .Z(net21273));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17503 (.I(net17502),
    .Z(net17503));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21363 (.I(\sa20_sr[6] ),
    .Z(net21363));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21282 (.I(\sa31_sub[2] ),
    .Z(net21282));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21277 (.I(\sa31_sub[5] ),
    .Z(net21277));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21375 (.I(\sa10_sub[7] ),
    .Z(net21375));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21278 (.I(\sa31_sub[4] ),
    .Z(net21278));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21281 (.I(\sa31_sub[2] ),
    .Z(net21281));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21279 (.I(\sa31_sub[3] ),
    .Z(net21279));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21299 (.I(\sa30_sr[7] ),
    .Z(net21299));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21283 (.I(\sa31_sub[1] ),
    .Z(net21283));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21300 (.I(net21299),
    .Z(net21300));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21284 (.I(\sa31_sub[0] ),
    .Z(net21284));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21541 (.I(net21540),
    .Z(net21541));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21285 (.I(\sa30_sub[7] ),
    .Z(net21285));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21296 (.I(\sa30_sub[1] ),
    .Z(net21296));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21288 (.I(\sa30_sub[6] ),
    .Z(net21288));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21302 (.I(\sa30_sr[4] ),
    .Z(net21302));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21289 (.I(\sa30_sub[5] ),
    .Z(net21289));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21540 (.I(net21531),
    .Z(net21540));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21290 (.I(\sa30_sub[4] ),
    .Z(net21290));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21303 (.I(\sa30_sr[4] ),
    .Z(net21303));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21292 (.I(\sa30_sub[2] ),
    .Z(net21292));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21291 (.I(\sa30_sub[3] ),
    .Z(net21291));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21353 (.I(\sa21_sr[3] ),
    .Z(net21353));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21295 (.I(\sa30_sub[1] ),
    .Z(net21295));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21297 (.I(\sa30_sub[0] ),
    .Z(net21297));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21298 (.I(\sa30_sr[7] ),
    .Z(net21298));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21301 (.I(\sa30_sr[5] ),
    .Z(net21301));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17501 (.I(_00981_),
    .Z(net17501));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21348 (.I(\sa21_sr[6] ),
    .Z(net21348));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21537 (.I(net21535),
    .Z(net21537));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21345 (.I(\sa20_sub[0] ),
    .Z(net21345));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21307 (.I(\sa30_sr[2] ),
    .Z(net21307));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21304 (.I(\sa30_sr[3] ),
    .Z(net21304));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21318 (.I(\sa21_sub[5] ),
    .Z(net21318));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place21310 (.I(\sa30_sr[1] ),
    .Z(net21310));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21342 (.I(\sa20_sub[1] ),
    .Z(net21342));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21312 (.I(\sa30_sr[0] ),
    .Z(net21312));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21314 (.I(\sa21_sub[7] ),
    .Z(net21314));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21315 (.I(\sa21_sub[7] ),
    .Z(net21315));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21316 (.I(\sa21_sub[6] ),
    .Z(net21316));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21319 (.I(\sa21_sub[5] ),
    .Z(net21319));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21317 (.I(\sa21_sub[5] ),
    .Z(net21317));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21320 (.I(\sa21_sub[4] ),
    .Z(net21320));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21334 (.I(\sa20_sub[7] ),
    .Z(net21334));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21331 (.I(\sa21_sub[0] ),
    .Z(net21331));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21328 (.I(\sa21_sub[1] ),
    .Z(net21328));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17314 (.I(_14469_),
    .Z(net17314));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21321 (.I(\sa21_sub[3] ),
    .Z(net21321));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17313 (.I(_14469_),
    .Z(net17313));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21536 (.I(net21535),
    .Z(net21536));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21325 (.I(\sa21_sub[2] ),
    .Z(net21325));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21324 (.I(\sa21_sub[2] ),
    .Z(net21324));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21326 (.I(\sa21_sub[1] ),
    .Z(net21326));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21327 (.I(\sa21_sub[1] ),
    .Z(net21327));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21329 (.I(\sa21_sub[0] ),
    .Z(net21329));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place21330 (.I(\sa21_sub[0] ),
    .Z(net21330));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21333 (.I(\sa20_sub[7] ),
    .Z(net21333));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21332 (.I(\sa20_sub[7] ),
    .Z(net21332));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place21493 (.I(net21490),
    .Z(net21493));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21340 (.I(\sa20_sub[2] ),
    .Z(net21340));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21335 (.I(\sa20_sub[6] ),
    .Z(net21335));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21356 (.I(\sa21_sr[2] ),
    .Z(net21356));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21336 (.I(\sa20_sub[5] ),
    .Z(net21336));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer189 (.I(\sa02_sr[0] ),
    .Z(net649));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21337 (.I(\sa20_sub[4] ),
    .Z(net21337));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17500 (.I(_00981_),
    .Z(net17500));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21338 (.I(\sa20_sub[3] ),
    .Z(net21338));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21339 (.I(\sa20_sub[2] ),
    .Z(net21339));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17320 (.I(_12999_),
    .Z(net17320));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21343 (.I(\sa20_sub[1] ),
    .Z(net21343));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21347 (.I(net21346),
    .Z(net21347));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21344 (.I(\sa20_sub[0] ),
    .Z(net21344));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21346 (.I(\sa21_sr[7] ),
    .Z(net21346));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21365 (.I(\sa20_sr[3] ),
    .Z(net21365));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21492 (.I(net21490),
    .Z(net21492));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21351 (.I(\sa21_sr[4] ),
    .Z(net21351));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21349 (.I(net21348),
    .Z(net21349));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17294 (.I(_15376_),
    .Z(net17294));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21350 (.I(\sa21_sr[5] ),
    .Z(net21350));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17293 (.I(_15376_),
    .Z(net17293));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17281 (.I(_01813_),
    .Z(net17281));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21366 (.I(\sa20_sr[3] ),
    .Z(net21366));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21355 (.I(\sa21_sr[2] ),
    .Z(net21355));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21352 (.I(\sa21_sr[3] ),
    .Z(net21352));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21360 (.I(net21359),
    .Z(net21360));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21354 (.I(\sa21_sr[2] ),
    .Z(net21354));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21358 (.I(\sa21_sr[1] ),
    .Z(net21358));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21357 (.I(\sa21_sr[1] ),
    .Z(net21357));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21394 (.I(net21393),
    .Z(net21394));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21359 (.I(\sa21_sr[0] ),
    .Z(net21359));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21361 (.I(\sa20_sr[7] ),
    .Z(net21361));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21362 (.I(\sa20_sr[7] ),
    .Z(net21362));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place21372 (.I(net21371),
    .Z(net21372));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place21371 (.I(\sa20_sr[0] ),
    .Z(net21371));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17289 (.I(_00559_),
    .Z(net17289));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21401 (.I(\sa11_sr[7] ),
    .Z(net21401));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21364 (.I(\sa20_sr[4] ),
    .Z(net21364));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21389 (.I(net21387),
    .Z(net21389));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21380 (.I(\sa10_sub[2] ),
    .Z(net21380));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21374 (.I(\sa10_sub[7] ),
    .Z(net21374));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21403 (.I(net21402),
    .Z(net21403));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21368 (.I(\sa20_sr[1] ),
    .Z(net21368));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21367 (.I(\sa20_sr[2] ),
    .Z(net21367));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place21370 (.I(\sa20_sr[0] ),
    .Z(net21370));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21369 (.I(\sa20_sr[0] ),
    .Z(net21369));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21402 (.I(net21401),
    .Z(net21402));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21373 (.I(\sa10_sub[7] ),
    .Z(net21373));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21385 (.I(net21384),
    .Z(net21385));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21381 (.I(\sa10_sub[2] ),
    .Z(net21381));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21376 (.I(\sa10_sub[6] ),
    .Z(net21376));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21386 (.I(\sa12_sr[7] ),
    .Z(net21386));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21377 (.I(\sa10_sub[5] ),
    .Z(net21377));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21378 (.I(\sa10_sub[4] ),
    .Z(net21378));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21379 (.I(\sa10_sub[3] ),
    .Z(net21379));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21411 (.I(net21410),
    .Z(net21411));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21382 (.I(\sa10_sub[1] ),
    .Z(net21382));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21395 (.I(\sa12_sr[2] ),
    .Z(net21395));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21383 (.I(\sa10_sub[0] ),
    .Z(net21383));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21388 (.I(net21387),
    .Z(net21388));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place21384 (.I(\sa12_sr[7] ),
    .Z(net21384));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21387 (.I(\sa12_sr[6] ),
    .Z(net21387));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21390 (.I(\sa12_sr[4] ),
    .Z(net21390));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21391 (.I(\sa12_sr[3] ),
    .Z(net21391));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21392 (.I(\sa12_sr[3] ),
    .Z(net21392));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21466 (.I(\sa01_sr[1] ),
    .Z(net21466));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21393 (.I(\sa12_sr[2] ),
    .Z(net21393));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21396 (.I(\sa12_sr[1] ),
    .Z(net21396));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21399 (.I(\sa12_sr[0] ),
    .Z(net21399));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21397 (.I(\sa12_sr[1] ),
    .Z(net21397));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21398 (.I(\sa12_sr[0] ),
    .Z(net21398));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21400 (.I(\sa11_sr[7] ),
    .Z(net21400));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21491 (.I(net21490),
    .Z(net21491));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_29_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21429 (.I(net21428),
    .Z(net21429));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21405 (.I(\sa11_sr[5] ),
    .Z(net21405));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21408 (.I(\sa11_sr[2] ),
    .Z(net21408));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place21427 (.I(\sa10_sr[1] ),
    .Z(net21427));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21406 (.I(\sa11_sr[4] ),
    .Z(net21406));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21423 (.I(\sa10_sr[2] ),
    .Z(net21423));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21417 (.I(\sa10_sr[5] ),
    .Z(net21417));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21416 (.I(\sa10_sr[6] ),
    .Z(net21416));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21407 (.I(\sa11_sr[3] ),
    .Z(net21407));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place21428 (.I(\sa10_sr[1] ),
    .Z(net21428));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21412 (.I(net21410),
    .Z(net21412));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21410 (.I(\sa11_sr[0] ),
    .Z(net21410));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21436 (.I(\sa03_sr[7] ),
    .Z(net21436));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21415 (.I(\sa10_sr[7] ),
    .Z(net21415));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21420 (.I(\sa10_sr[3] ),
    .Z(net21420));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21430 (.I(\sa10_sr[0] ),
    .Z(net21430));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21419 (.I(\sa10_sr[3] ),
    .Z(net21419));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21418 (.I(\sa10_sr[4] ),
    .Z(net21418));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21435 (.I(net21433),
    .Z(net21435));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place21432 (.I(\sa10_sr[0] ),
    .Z(net21432));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21422 (.I(\sa10_sr[2] ),
    .Z(net21422));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21421 (.I(net21420),
    .Z(net21421));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21426 (.I(\sa10_sr[1] ),
    .Z(net21426));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21431 (.I(net21430),
    .Z(net21431));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21433 (.I(\sa03_sr[7] ),
    .Z(net21433));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21434 (.I(net21433),
    .Z(net21434));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21450 (.I(\sa02_sr[3] ),
    .Z(net21450));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place21490 (.I(ld_r),
    .Z(net21490));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21489 (.I(net21488),
    .Z(net21489));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21446 (.I(\sa02_sr[7] ),
    .Z(net21446));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21437 (.I(\sa03_sr[4] ),
    .Z(net21437));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21438 (.I(\sa03_sr[3] ),
    .Z(net21438));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21445 (.I(net21444),
    .Z(net21445));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place21442 (.I(\sa03_sr[1] ),
    .Z(net21442));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21440 (.I(\sa03_sr[2] ),
    .Z(net21440));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21441 (.I(\sa03_sr[1] ),
    .Z(net21441));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17362 (.I(_07016_),
    .Z(net17362));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21443 (.I(\sa03_sr[0] ),
    .Z(net21443));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17433 (.I(_03156_),
    .Z(net17433));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21444 (.I(\sa02_sr[7] ),
    .Z(net21444));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21447 (.I(\sa02_sr[6] ),
    .Z(net21447));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place21486 (.I(net21482),
    .Z(net21486));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21457 (.I(net649),
    .Z(net21457));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21449 (.I(\sa02_sr[4] ),
    .Z(net21449));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21448 (.I(\sa02_sr[4] ),
    .Z(net21448));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21464 (.I(\sa01_sr[2] ),
    .Z(net21464));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21452 (.I(\sa02_sr[2] ),
    .Z(net21452));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21485 (.I(net21482),
    .Z(net21485));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21451 (.I(\sa02_sr[2] ),
    .Z(net21451));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21455 (.I(net21454),
    .Z(net21455));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21453 (.I(\sa02_sr[1] ),
    .Z(net21453));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place21454 (.I(\sa02_sr[0] ),
    .Z(net21454));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21484 (.I(net21482),
    .Z(net21484));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21459 (.I(net21458),
    .Z(net21459));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21465 (.I(\sa01_sr[2] ),
    .Z(net21465));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21460 (.I(\sa01_sr[5] ),
    .Z(net21460));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17363 (.I(_06957_),
    .Z(net17363));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21469 (.I(\sa01_sr[0] ),
    .Z(net21469));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21480 (.I(\sa00_sr[0] ),
    .Z(net21480));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21461 (.I(\sa01_sr[4] ),
    .Z(net21461));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17280 (.I(_01819_),
    .Z(net17280));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17278 (.I(_01826_),
    .Z(net17278));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17360 (.I(_07054_),
    .Z(net17360));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21471 (.I(\sa00_sr[7] ),
    .Z(net21471));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21462 (.I(\sa01_sr[3] ),
    .Z(net21462));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21463 (.I(\sa01_sr[2] ),
    .Z(net21463));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21468 (.I(\sa01_sr[0] ),
    .Z(net21468));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21467 (.I(\sa01_sr[0] ),
    .Z(net21467));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21476 (.I(\sa00_sr[2] ),
    .Z(net21476));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21470 (.I(\sa00_sr[7] ),
    .Z(net21470));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17423 (.I(_03267_),
    .Z(net17423));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21479 (.I(\sa00_sr[1] ),
    .Z(net21479));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21472 (.I(\sa00_sr[5] ),
    .Z(net21472));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21478 (.I(net21477),
    .Z(net21478));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21473 (.I(\sa00_sr[4] ),
    .Z(net21473));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21475 (.I(\sa00_sr[2] ),
    .Z(net21475));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21474 (.I(\sa00_sr[3] ),
    .Z(net21474));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17393 (.I(_04351_),
    .Z(net17393));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17376 (.I(_06205_),
    .Z(net17376));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17368 (.I(_06574_),
    .Z(net17368));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17367 (.I(_06819_),
    .Z(net17367));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17364 (.I(_06889_),
    .Z(net17364));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place21477 (.I(\sa00_sr[1] ),
    .Z(net21477));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21481 (.I(\sa00_sr[0] ),
    .Z(net21481));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17365 (.I(_06877_),
    .Z(net17365));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21483 (.I(net21482),
    .Z(net21483));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21482 (.I(ld_r),
    .Z(net21482));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21544 (.I(net21542),
    .Z(net21544));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_32_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17487 (.I(_01290_),
    .Z(net17487));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17513 (.I(net17512),
    .Z(net17513));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17407 (.I(_03904_),
    .Z(net17407));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17432 (.I(_03169_),
    .Z(net17432));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17321 (.I(_12633_),
    .Z(net17321));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17200 (.I(_15268_),
    .Z(net17200));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place21539 (.I(net21538),
    .Z(net21539));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17249 (.I(_03493_),
    .Z(net17249));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17275 (.I(_01859_),
    .Z(net17275));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place17225 (.I(net17224),
    .Z(net17225));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17273 (.I(_01908_),
    .Z(net17273));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17319 (.I(_13161_),
    .Z(net17319));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17318 (.I(_13188_),
    .Z(net17318));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17245 (.I(_03572_),
    .Z(net17245));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17247 (.I(_03528_),
    .Z(net17247));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place17271 (.I(_01993_),
    .Z(net17271));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17265 (.I(_02842_),
    .Z(net17265));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17323 (.I(_12505_),
    .Z(net17323));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17322 (.I(_12505_),
    .Z(net17322));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17269 (.I(_02428_),
    .Z(net17269));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17268 (.I(_02563_),
    .Z(net17268));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17324 (.I(_12354_),
    .Z(net17324));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17331 (.I(_12238_),
    .Z(net17331));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17326 (.I(_12332_),
    .Z(net17326));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17210 (.I(_01860_),
    .Z(net17210));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17316 (.I(_14465_),
    .Z(net17316));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17251 (.I(_03430_),
    .Z(net17251));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17218 (.I(_15176_),
    .Z(net17218));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17223 (.I(_12511_),
    .Z(net17223));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17208 (.I(_01955_),
    .Z(net17208));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17204 (.I(_03654_),
    .Z(net17204));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place17224 (.I(_12509_),
    .Z(net17224));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17279 (.I(_01819_),
    .Z(net17279));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17221 (.I(_12665_),
    .Z(net17221));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17274 (.I(_01878_),
    .Z(net17274));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17272 (.I(_01928_),
    .Z(net17272));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17199 (.I(_01747_),
    .Z(net17199));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17267 (.I(_02609_),
    .Z(net17267));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17260 (.I(_03157_),
    .Z(net17260));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17258 (.I(_03268_),
    .Z(net17258));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17257 (.I(_03294_),
    .Z(net17257));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17214 (.I(_00553_),
    .Z(net17214));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17256 (.I(_03317_),
    .Z(net17256));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17211 (.I(_01802_),
    .Z(net17211));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place17202 (.I(_12550_),
    .Z(net17202));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17286 (.I(_01690_),
    .Z(net17286));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17240 (.I(_04251_),
    .Z(net17240));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17226 (.I(_12458_),
    .Z(net17226));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17263 (.I(_02849_),
    .Z(net17263));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17212 (.I(_00565_),
    .Z(net17212));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17254 (.I(_03371_),
    .Z(net17254));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17231 (.I(_11712_),
    .Z(net17231));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17207 (.I(_03158_),
    .Z(net17207));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17217 (.I(_15267_),
    .Z(net17217));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17213 (.I(_00563_),
    .Z(net17213));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17209 (.I(_01909_),
    .Z(net17209));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place17222 (.I(_12534_),
    .Z(net17222));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20714 (.I(_07639_),
    .Z(net20714));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20710 (.I(net20708),
    .Z(net20710));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20715 (.I(_07639_),
    .Z(net20715));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20707 (.I(_15645_[0]),
    .Z(net20707));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20704 (.I(net20703),
    .Z(net20704));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place20703 (.I(net660),
    .Z(net20703));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18306 (.I(_12974_),
    .Z(net18306));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18827 (.I(net18813),
    .Z(net18827));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18826 (.I(net18813),
    .Z(net18826));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18790 (.I(_14414_),
    .Z(net18790));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18789 (.I(net18786),
    .Z(net18789));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18307 (.I(_12972_),
    .Z(net18307));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18456 (.I(_06166_),
    .Z(net18456));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18471 (.I(_05440_),
    .Z(net18471));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18477 (.I(_05392_),
    .Z(net18477));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18480 (.I(_05391_),
    .Z(net18480));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18513 (.I(_04098_),
    .Z(net18513));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18515 (.I(_04049_),
    .Z(net18515));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18516 (.I(_03985_),
    .Z(net18516));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18519 (.I(_03976_),
    .Z(net18519));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18521 (.I(_03976_),
    .Z(net18521));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18520 (.I(_03976_),
    .Z(net18520));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18525 (.I(_03928_),
    .Z(net18525));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18533 (.I(net18532),
    .Z(net18533));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18532 (.I(_03891_),
    .Z(net18532));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18599 (.I(net691),
    .Z(net18599));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18598 (.I(net18586),
    .Z(net18598));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18557 (.I(net18549),
    .Z(net18557));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18556 (.I(net18549),
    .Z(net18556));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18555 (.I(net18549),
    .Z(net18555));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18554 (.I(net18549),
    .Z(net18554));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18553 (.I(net18549),
    .Z(net18553));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18552 (.I(net18549),
    .Z(net18552));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18551 (.I(net18549),
    .Z(net18551));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18550 (.I(net18549),
    .Z(net18550));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place18549 (.I(_03860_),
    .Z(net18549));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18821 (.I(net18820),
    .Z(net18821));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18811 (.I(net18806),
    .Z(net18811));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place18812 (.I(net18806),
    .Z(net18812));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18859 (.I(net18854),
    .Z(net18859));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18858 (.I(net18854),
    .Z(net18858));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18857 (.I(net18854),
    .Z(net18857));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18856 (.I(net18854),
    .Z(net18856));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18855 (.I(net18854),
    .Z(net18855));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18835 (.I(net18834),
    .Z(net18835));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18832 (.I(_13296_),
    .Z(net18832));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18922 (.I(net18919),
    .Z(net18922));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place18921 (.I(net18919),
    .Z(net18921));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place18249 (.I(_14435_),
    .Z(net18249));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19157 (.I(net19155),
    .Z(net19157));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19158 (.I(net19155),
    .Z(net19158));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place19159 (.I(net19155),
    .Z(net19159));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20461 (.I(_09742_),
    .Z(net20461));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20462 (.I(net20461),
    .Z(net20462));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20463 (.I(net20461),
    .Z(net20463));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20464 (.I(net20461),
    .Z(net20464));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place20465 (.I(_09742_),
    .Z(net20465));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20466 (.I(net20465),
    .Z(net20466));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20467 (.I(net20465),
    .Z(net20467));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20468 (.I(net20465),
    .Z(net20468));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20469 (.I(net20465),
    .Z(net20469));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20589 (.I(_07630_),
    .Z(net20589));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place20590 (.I(_07630_),
    .Z(net20590));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20591 (.I(net20590),
    .Z(net20591));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place20592 (.I(_07630_),
    .Z(net20592));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21083 (.I(_10378_),
    .Z(net21083));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21084 (.I(_10378_),
    .Z(net21084));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21085 (.I(net21084),
    .Z(net21085));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21086 (.I(_10378_),
    .Z(net21086));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21087 (.I(_10378_),
    .Z(net21087));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21088 (.I(net21087),
    .Z(net21088));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21089 (.I(_10378_),
    .Z(net21089));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21090 (.I(net21089),
    .Z(net21090));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21091 (.I(_10378_),
    .Z(net21091));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place21092 (.I(net21091),
    .Z(net21092));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place21093 (.I(_10378_),
    .Z(net21093));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21094 (.I(_10378_),
    .Z(net21094));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place21095 (.I(_10378_),
    .Z(net21095));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_36_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_37_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_39_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_42_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_43_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_45_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_49_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_53_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_54_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_57_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_58_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_61_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_64_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_67_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_71_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_75_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_77_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_81_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_82_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_86_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_91_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_96_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_102_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_106_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_111_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_111_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_123_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_123_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_125_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_126_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_127_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_130_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_130_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_138_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_139_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_141_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_141_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_142_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_143_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_143_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_144_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_150_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_152_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_154_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_154_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_159_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_159_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_160_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_160_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_161_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_161_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_166_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_167_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_168_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_168_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_169_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_169_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_178_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_185_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_185_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_191_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_205_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_205_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_206_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_206_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_207_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_207_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_209_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_221_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_223_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_223_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_231_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_239_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_239_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_241_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_246_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_246_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_249_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_249_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_250_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_250_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_252_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_252_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_254_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_254_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_257_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_257_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_270_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_270_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_273_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_273_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_277_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_277_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_283_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_283_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_289_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_289_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_290_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_290_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_301_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_301_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_303_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_303_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_313_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_315_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_315_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_318_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_318_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_349_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_349_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_352_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_352_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_354_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_354_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_355_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_355_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_358_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_358_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_362_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_362_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_363_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_363_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_369_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_369_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_370_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_370_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_372_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_372_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_376_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_376_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_377_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_377_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_378_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_378_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_382_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_382_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_385_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_385_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_389_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_389_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_390_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_390_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_394_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_394_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_399_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_399_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_410_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_410_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_411_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_411_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_412_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_412_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_413_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_413_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_415_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_415_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_417_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_417_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_423_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_423_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_424_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_424_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_425_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_425_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_431_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_431_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_0__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_1__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_2__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_3__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_4__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_5__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_6__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_7__f_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_8__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_9__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_10__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_11__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_12__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_13__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_14__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_15__f_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_16__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_17__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_18__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_19__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_20__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_21__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_22__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_23__f_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_24__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_25__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_26__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_27__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_28__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_29__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_30__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_5_31__f_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload0 (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload1 (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload2 (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload3 (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload4 (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload5 (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload6 (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload7 (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload8 (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload9 (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload10 (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 clkload11 (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload12 (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload13 (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload14 (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload15 (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload16 (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload17 (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload18 (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload19 (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload20 (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload21 (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload22 (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload23 (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload24 (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload25 (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload26 (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload27 (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload28 (.I(clknet_leaf_410_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload29 (.I(clknet_leaf_411_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload30 (.I(clknet_leaf_412_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload31 (.I(clknet_leaf_413_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload32 (.I(clknet_leaf_415_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload33 (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload34 (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload35 (.I(clknet_leaf_370_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload36 (.I(clknet_leaf_372_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload37 (.I(clknet_leaf_377_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload38 (.I(clknet_leaf_378_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload39 (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload40 (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload41 (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload42 (.I(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload43 (.I(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload44 (.I(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload45 (.I(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload46 (.I(clknet_leaf_141_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload47 (.I(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload48 (.I(clknet_leaf_143_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload49 (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload50 (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload51 (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload52 (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload53 (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload54 (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload55 (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload56 (.I(clknet_leaf_159_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload57 (.I(clknet_leaf_277_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload58 (.I(clknet_leaf_289_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload59 (.I(clknet_leaf_205_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload60 (.I(clknet_leaf_206_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload61 (.I(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload62 (.I(clknet_leaf_246_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer1 (.I(_16169_[0]),
    .Z(net388));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2 (.I(_15935_[0]),
    .Z(net389));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer3 (.I(_00971_),
    .Z(net390));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer4 (.I(_16178_[0]),
    .Z(net391));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer5 (.I(_06929_),
    .Z(net392));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer6 (.I(_06818_),
    .Z(net393));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer134 (.I(_13706_),
    .Z(net526));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer8 (.I(_13642_),
    .Z(net395));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer9 (.I(net19241),
    .Z(net396));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer10 (.I(_16178_[0]),
    .Z(net397));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer11 (.I(_11993_),
    .Z(net398));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer12 (.I(_15866_[0]),
    .Z(net399));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer13 (.I(net18200),
    .Z(net400));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer14 (.I(net18200),
    .Z(net401));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer15 (.I(_15868_[0]),
    .Z(net402));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer16 (.I(_16038_[0]),
    .Z(net403));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer17 (.I(_16038_[0]),
    .Z(net404));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer18 (.I(_16038_[0]),
    .Z(net405));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer19 (.I(_15871_[0]),
    .Z(net406));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer20 (.I(_13782_),
    .Z(net407));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer21 (.I(_13782_),
    .Z(net408));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer22 (.I(net17698),
    .Z(net409));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 rebuffer23 (.I(_13796_),
    .Z(net410));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer24 (.I(net630),
    .Z(net411));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer25 (.I(_15337_),
    .Z(net412));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer26 (.I(_15337_),
    .Z(net413));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer27 (.I(_12814_),
    .Z(net414));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer28 (.I(_16176_[0]),
    .Z(net415));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer29 (.I(net19798),
    .Z(net416));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer30 (.I(net19798),
    .Z(net417));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer31 (.I(_03974_),
    .Z(net418));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone40 (.I(net19204),
    .Z(net427));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer41 (.I(_01106_),
    .Z(net428));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer43 (.I(net19242),
    .Z(net430));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer52 (.I(_06817_),
    .Z(net439));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer53 (.I(_07181_),
    .Z(net440));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer54 (.I(_15971_[0]),
    .Z(net441));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer55 (.I(_15971_[0]),
    .Z(net442));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer56 (.I(net689),
    .Z(net443));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer57 (.I(_02410_),
    .Z(net444));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer58 (.I(_02534_),
    .Z(net445));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer59 (.I(_02534_),
    .Z(net446));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer60 (.I(_02605_),
    .Z(net447));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer61 (.I(_02605_),
    .Z(net448));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone62 (.I(_02367_),
    .Z(net449));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone63 (.I(_02367_),
    .Z(net450));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer75 (.I(net17701),
    .Z(net462));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer79 (.I(_01730_),
    .Z(net466));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer80 (.I(_15940_[0]),
    .Z(net467));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer81 (.I(_01722_),
    .Z(net468));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer82 (.I(_01568_),
    .Z(net469));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer84 (.I(_03881_),
    .Z(net471));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer86 (.I(_06963_),
    .Z(net473));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer87 (.I(_06963_),
    .Z(net474));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer88 (.I(_15738_[0]),
    .Z(net475));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer98 (.I(_11997_),
    .Z(net485));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer99 (.I(_11997_),
    .Z(net486));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer100 (.I(_12227_),
    .Z(net487));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer101 (.I(_12227_),
    .Z(net488));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer102 (.I(_06123_),
    .Z(net489));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer103 (.I(_06085_),
    .Z(net490));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer104 (.I(_06199_),
    .Z(net491));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer105 (.I(net17804),
    .Z(net492));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 rebuffer107 (.I(_15673_[0]),
    .Z(net494));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer108 (.I(_15682_[0]),
    .Z(net495));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer109 (.I(_15682_[0]),
    .Z(net496));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer110 (.I(net19425),
    .Z(net497));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer112 (.I(_10622_),
    .Z(net499));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer113 (.I(_10537_),
    .Z(net500));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer114 (.I(_15674_[0]),
    .Z(net501));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer115 (.I(_15679_[0]),
    .Z(net502));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer116 (.I(net20918),
    .Z(net503));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer117 (.I(net21097),
    .Z(net504));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer118 (.I(net19400),
    .Z(net505));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer119 (.I(net19400),
    .Z(net506));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer120 (.I(net19400),
    .Z(net507));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer130 (.I(net18958),
    .Z(net517));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer131 (.I(net18958),
    .Z(net518));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer132 (.I(net18958),
    .Z(net519));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer133 (.I(_06931_),
    .Z(net520));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 clone134 (.A1(net19462),
    .A2(net519),
    .ZN(net521));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer141 (.I(net527),
    .Z(net528));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer144 (.I(_04024_),
    .Z(net531));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer145 (.I(_13052_),
    .Z(net532));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer146 (.I(_13052_),
    .Z(net533));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer147 (.I(_09793_),
    .Z(net534));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer148 (.I(_09849_),
    .Z(net535));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold149 (.I(key[123]),
    .Z(net536));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold150 (.I(key[120]),
    .Z(net537));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold151 (.I(key[121]),
    .Z(net538));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold152 (.I(key[122]),
    .Z(net539));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold153 (.I(key[117]),
    .Z(net540));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold154 (.I(key[60]),
    .Z(net541));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold155 (.I(key[47]),
    .Z(net542));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold156 (.I(text_in[112]),
    .Z(net543));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold157 (.I(key[35]),
    .Z(net544));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold158 (.I(key[57]),
    .Z(net545));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold159 (.I(key[126]),
    .Z(net546));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold160 (.I(key[56]),
    .Z(net547));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold161 (.I(key[99]),
    .Z(net548));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold162 (.I(key[59]),
    .Z(net549));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold163 (.I(key[46]),
    .Z(net550));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold164 (.I(key[63]),
    .Z(net551));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold165 (.I(key[32]),
    .Z(net552));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold166 (.I(key[110]),
    .Z(net553));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold167 (.I(key[96]),
    .Z(net554));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold168 (.I(text_in[95]),
    .Z(net555));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold169 (.I(text_in[55]),
    .Z(net556));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold170 (.I(text_in[94]),
    .Z(net557));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold171 (.I(text_in[67]),
    .Z(net558));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold172 (.I(text_in[65]),
    .Z(net559));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold173 (.I(rst),
    .Z(net560));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold174 (.I(text_in[91]),
    .Z(net561));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold175 (.I(key[109]),
    .Z(net562));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold176 (.I(text_in[97]),
    .Z(net563));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold177 (.I(text_in[96]),
    .Z(net564));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold178 (.I(key[125]),
    .Z(net565));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold179 (.I(key[103]),
    .Z(net566));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold180 (.I(text_in[11]),
    .Z(net567));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold181 (.I(key[53]),
    .Z(net568));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold182 (.I(key[48]),
    .Z(net569));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold183 (.I(key[44]),
    .Z(net570));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold184 (.I(text_in[72]),
    .Z(net571));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold185 (.I(key[54]),
    .Z(net572));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold186 (.I(text_in[100]),
    .Z(net573));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold187 (.I(text_in[113]),
    .Z(net574));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold188 (.I(text_in[71]),
    .Z(net575));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold189 (.I(key[41]),
    .Z(net576));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold190 (.I(text_in[76]),
    .Z(net577));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold191 (.I(text_in[84]),
    .Z(net578));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold192 (.I(text_in[73]),
    .Z(net579));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold193 (.I(key[43]),
    .Z(net580));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold194 (.I(key[111]),
    .Z(net581));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold195 (.I(key[55]),
    .Z(net582));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold196 (.I(text_in[74]),
    .Z(net583));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold197 (.I(key[50]),
    .Z(net584));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold198 (.I(key[127]),
    .Z(net585));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold199 (.I(key[62]),
    .Z(net586));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold200 (.I(key[49]),
    .Z(net587));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold201 (.I(key[124]),
    .Z(net588));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold202 (.I(text_in[82]),
    .Z(net589));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold203 (.I(text_in[81]),
    .Z(net590));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold204 (.I(text_in[86]),
    .Z(net591));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold205 (.I(text_in[15]),
    .Z(net592));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold206 (.I(text_in[85]),
    .Z(net593));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold207 (.I(text_in[87]),
    .Z(net594));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold208 (.I(text_in[5]),
    .Z(net595));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold209 (.I(text_in[90]),
    .Z(net596));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold210 (.I(text_in[78]),
    .Z(net597));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold211 (.I(text_in[10]),
    .Z(net598));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold212 (.I(text_in[89]),
    .Z(net599));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold213 (.I(text_in[13]),
    .Z(net600));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold214 (.I(text_in[117]),
    .Z(net601));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold215 (.I(text_in[24]),
    .Z(net602));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer7 (.I(_12821_),
    .Z(net419));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer35 (.I(_15872_[0]),
    .Z(net423));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer46 (.I(net18318),
    .Z(net435));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer47 (.I(_12133_),
    .Z(net436));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer49 (.I(_01062_),
    .Z(net438));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer50 (.I(_01029_),
    .Z(net451));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer51 (.I(_01029_),
    .Z(net452));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer62 (.I(_00905_),
    .Z(net453));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer63 (.I(_15124_),
    .Z(net454));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer70 (.I(_16172_[0]),
    .Z(net461));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer71 (.I(_06709_),
    .Z(net463));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer72 (.I(_01963_),
    .Z(net464));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer73 (.I(net17767),
    .Z(net470));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer74 (.I(_01674_),
    .Z(net472));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer76 (.I(net18445),
    .Z(net476));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer77 (.I(_06908_),
    .Z(net477));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer83 (.I(_16043_[0]),
    .Z(net478));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer94 (.I(_04724_),
    .Z(net493));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer95 (.I(_04994_),
    .Z(net508));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer96 (.I(_16074_[0]),
    .Z(net509));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer97 (.I(net19609),
    .Z(net510));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer106 (.I(net19610),
    .Z(net511));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer121 (.I(_16082_[0]),
    .Z(net512));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer122 (.I(_04700_),
    .Z(net513));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer123 (.I(_04660_),
    .Z(net514));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer124 (.I(_03881_),
    .Z(net515));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer127 (.I(net18080),
    .Z(net523));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer128 (.I(_12267_),
    .Z(net524));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer129 (.I(_13826_),
    .Z(net525));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer135 (.I(_15804_[0]),
    .Z(net529));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer136 (.I(_13845_),
    .Z(net530));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer137 (.I(_13845_),
    .Z(net603));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer138 (.I(_15801_[0]),
    .Z(net604));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer139 (.I(net21432),
    .Z(net605));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer151 (.I(_03988_),
    .Z(net611));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer152 (.I(net18102),
    .Z(net612));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer153 (.I(net18102),
    .Z(net613));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer154 (.I(net18102),
    .Z(net614));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer155 (.I(net18102),
    .Z(net615));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer156 (.I(_04024_),
    .Z(net616));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer157 (.I(net17704),
    .Z(net617));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer158 (.I(_03903_),
    .Z(net618));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer159 (.I(net19242),
    .Z(net619));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer170 (.I(_13796_),
    .Z(net630));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer171 (.I(_13796_),
    .Z(net631));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer174 (.I(_13847_),
    .Z(net634));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer175 (.I(_13786_),
    .Z(net635));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 rebuffer176 (.I(_15813_[0]),
    .Z(net636));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer177 (.I(_13968_),
    .Z(net637));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone181 (.I(net18318),
    .Z(net641));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone182 (.A1(net19331),
    .A2(net645),
    .ZN(net642));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer183 (.I(net644),
    .Z(net643));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 clone184 (.A1(net19334),
    .A2(net435),
    .A3(net19330),
    .ZN(net644));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone185 (.I(net657),
    .Z(net645));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer186 (.I(_12128_),
    .Z(net646));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone187 (.I(_12128_),
    .Z(net647));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 clone188 (.I(_12212_),
    .Z(net648));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer190 (.I(_15431_),
    .Z(net650));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer191 (.I(_15874_[0]),
    .Z(net651));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer192 (.I(_04662_),
    .Z(net652));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer193 (.I(_04701_),
    .Z(net653));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer194 (.I(_12226_),
    .Z(net654));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer195 (.I(_12174_),
    .Z(net655));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer196 (.I(_15737_[0]),
    .Z(net656));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer197 (.I(net18315),
    .Z(net657));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer199 (.I(net19888),
    .Z(net659));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer200 (.I(_15650_[0]),
    .Z(net660));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer201 (.I(_15640_[0]),
    .Z(net661));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer202 (.I(_09884_),
    .Z(net662));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer203 (.I(net20471),
    .Z(net663));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer204 (.I(net20472),
    .Z(net664));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer205 (.I(\u0.w[2][25] ),
    .Z(net665));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer206 (.I(_15645_[0]),
    .Z(net666));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer208 (.I(net17902),
    .Z(net668));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer209 (.I(net17902),
    .Z(net669));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer220 (.I(_01750_),
    .Z(net680));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer221 (.I(_12140_),
    .Z(net681));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer222 (.I(_12293_),
    .Z(net682));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer223 (.I(_09915_),
    .Z(net683));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer224 (.I(\u0.w[2][24] ),
    .Z(net684));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer227 (.I(_15976_[0]),
    .Z(net687));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer228 (.I(_02428_),
    .Z(net688));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer229 (.I(net21347),
    .Z(net689));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer230 (.I(_02309_),
    .Z(net690));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone231 (.I(net693),
    .Z(net691));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone232 (.I(_02391_),
    .Z(net692));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer233 (.I(_02391_),
    .Z(net693));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_1 (.I(key[0]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_2 (.I(key[100]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_3 (.I(key[101]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_4 (.I(key[102]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_5 (.I(key[102]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_6 (.I(key[121]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_7 (.I(key[123]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_8 (.I(key[125]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_9 (.I(key[126]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_10 (.I(key[15]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_11 (.I(key[1]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_12 (.I(key[22]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_13 (.I(key[2]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_14 (.I(key[30]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_15 (.I(key[33]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_16 (.I(key[33]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_17 (.I(key[35]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_18 (.I(key[35]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_19 (.I(key[43]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_20 (.I(key[58]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_21 (.I(key[62]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_22 (.I(key[69]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_23 (.I(key[80]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_24 (.I(key[85]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_25 (.I(key[87]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_26 (.I(key[91]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_27 (.I(key[93]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_28 (.I(key[97]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_29 (.I(rst));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_30 (.I(text_in[100]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_31 (.I(text_in[109]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_32 (.I(text_in[109]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_33 (.I(text_in[117]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_34 (.I(text_in[118]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_35 (.I(text_in[118]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_36 (.I(text_in[119]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_37 (.I(text_in[119]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_38 (.I(text_in[120]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_39 (.I(text_in[120]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_40 (.I(text_in[124]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_41 (.I(text_in[126]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_42 (.I(text_in[126]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_43 (.I(text_in[3]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_44 (.I(text_in[52]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_45 (.I(text_in[52]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_46 (.I(text_in[79]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_47 (.I(text_in[91]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_48 (.I(text_in[94]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_49 (.I(text_in[95]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_50 (.I(key[58]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_51 (.I(text_in[113]));
 gf180mcu_fd_sc_mcu9t5v0__antenna ANTENNA_52 (.I(text_in[13]));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_2169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_2201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_2205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_2166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_2194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_2203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_2147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_2181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_2209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_2170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_2185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_2140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_2212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_2179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_2211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_2139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_2145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_2165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_2197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_2213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_2210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_2214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_2199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_2200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_2124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_2125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_2121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_2129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_2128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_2127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_2131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_2135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_2126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_2122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_2130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_2132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_235_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_235_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_235_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_235_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_235_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_236_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_236_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_236_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_236_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_236_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_236_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_237_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_237_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_237_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_237_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_237_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_238_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_238_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_238_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_238_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_238_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_238_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_239_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_239_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_239_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_239_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_239_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_240_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_240_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_240_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_240_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_240_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_240_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_241_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_241_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_241_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_241_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_241_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_242_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_242_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_242_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_242_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_242_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_242_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_243_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_243_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_243_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_243_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_243_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_244_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_244_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_244_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_244_2152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_244_2216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_244_2220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_245_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_2120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_245_2138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_245_2202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_245_2218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_245_2220 ();
endmodule
