module riscv (clk,
    memread,
    memwrite,
    reset,
    suspend,
    aluout,
    instr,
    pc,
    readdata,
    writedata);
 input clk;
 output memread;
 output memwrite;
 input reset;
 output suspend;
 output [31:0] aluout;
 input [31:0] instr;
 output [31:0] pc;
 input [31:0] readdata;
 output [31:0] writedata;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_79_clk;
 wire net480;
 wire net513;
 wire net510;
 wire net543;
 wire net542;
 wire net509;
 wire net490;
 wire net489;
 wire net486;
 wire net484;
 wire net483;
 wire net545;
 wire net479;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_18_clk;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire _01029_;
 wire _01030_;
 wire clknet_6_46__leaf_clk;
 wire _01032_;
 wire _01033_;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire _01036_;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire _01045_;
 wire clknet_6_39__leaf_clk;
 wire _01047_;
 wire _01048_;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire _01052_;
 wire _01053_;
 wire clknet_6_35__leaf_clk;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire clknet_6_34__leaf_clk;
 wire _01060_;
 wire clknet_6_33__leaf_clk;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire clknet_6_32__leaf_clk;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire _01073_;
 wire _01074_;
 wire clknet_6_27__leaf_clk;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire clknet_6_26__leaf_clk;
 wire _01081_;
 wire _01082_;
 wire clknet_6_25__leaf_clk;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire _01092_;
 wire clknet_6_22__leaf_clk;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire clknet_6_21__leaf_clk;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire clknet_6_20__leaf_clk;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire _01122_;
 wire _01123_;
 wire clknet_6_17__leaf_clk;
 wire _01125_;
 wire _01126_;
 wire clknet_6_16__leaf_clk;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire _01140_;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire _01144_;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire _01147_;
 wire _01148_;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire _01154_;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_4_15_0_clk;
 wire _01160_;
 wire _01161_;
 wire clknet_4_14_0_clk;
 wire clknet_4_13_0_clk;
 wire _01164_;
 wire _01165_;
 wire clknet_4_12_0_clk;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire clknet_4_11_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_7_0_clk;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire clknet_4_6_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_4_0_clk;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire clknet_4_3_0_clk;
 wire _01189_;
 wire clknet_4_2_0_clk;
 wire _01191_;
 wire clknet_4_1_0_clk;
 wire clknet_4_0_0_clk;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire clknet_0_clk;
 wire clknet_leaf_712_clk;
 wire clknet_leaf_711_clk;
 wire clknet_leaf_705_clk;
 wire clknet_leaf_704_clk;
 wire clknet_leaf_702_clk;
 wire _01205_;
 wire _01206_;
 wire clknet_leaf_700_clk;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire clknet_leaf_698_clk;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire clknet_leaf_697_clk;
 wire clknet_leaf_694_clk;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire clknet_leaf_693_clk;
 wire clknet_leaf_692_clk;
 wire clknet_leaf_689_clk;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire clknet_leaf_687_clk;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire clknet_leaf_685_clk;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire clknet_leaf_684_clk;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire clknet_leaf_682_clk;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire clknet_leaf_680_clk;
 wire _01290_;
 wire clknet_leaf_679_clk;
 wire clknet_leaf_678_clk;
 wire _01293_;
 wire _01294_;
 wire clknet_leaf_675_clk;
 wire _01296_;
 wire _01297_;
 wire clknet_leaf_673_clk;
 wire clknet_leaf_670_clk;
 wire _01300_;
 wire clknet_leaf_668_clk;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire clknet_leaf_665_clk;
 wire clknet_leaf_664_clk;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire clknet_leaf_662_clk;
 wire clknet_leaf_658_clk;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire clknet_leaf_657_clk;
 wire clknet_leaf_656_clk;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire clknet_leaf_655_clk;
 wire clknet_leaf_654_clk;
 wire clknet_leaf_652_clk;
 wire _01329_;
 wire clknet_leaf_651_clk;
 wire clknet_leaf_649_clk;
 wire clknet_leaf_647_clk;
 wire _01333_;
 wire _01334_;
 wire clknet_leaf_645_clk;
 wire clknet_leaf_642_clk;
 wire clknet_leaf_641_clk;
 wire _01338_;
 wire _01339_;
 wire clknet_leaf_640_clk;
 wire clknet_leaf_639_clk;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire clknet_leaf_638_clk;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire clknet_leaf_637_clk;
 wire clknet_leaf_633_clk;
 wire clknet_leaf_632_clk;
 wire _01356_;
 wire clknet_leaf_631_clk;
 wire clknet_leaf_630_clk;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire clknet_leaf_629_clk;
 wire clknet_leaf_628_clk;
 wire _01365_;
 wire _01366_;
 wire clknet_leaf_626_clk;
 wire _01368_;
 wire clknet_leaf_624_clk;
 wire _01370_;
 wire clknet_leaf_623_clk;
 wire clknet_leaf_622_clk;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire clknet_leaf_618_clk;
 wire clknet_leaf_616_clk;
 wire _01380_;
 wire clknet_leaf_614_clk;
 wire clknet_leaf_611_clk;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire clknet_leaf_609_clk;
 wire _01387_;
 wire _01388_;
 wire clknet_leaf_608_clk;
 wire clknet_leaf_598_clk;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire clknet_leaf_597_clk;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire clknet_leaf_596_clk;
 wire _01409_;
 wire clknet_leaf_595_clk;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire clknet_leaf_592_clk;
 wire clknet_leaf_591_clk;
 wire clknet_leaf_590_clk;
 wire clknet_leaf_588_clk;
 wire _01420_;
 wire _01421_;
 wire clknet_leaf_587_clk;
 wire clknet_leaf_584_clk;
 wire _01424_;
 wire _01425_;
 wire clknet_leaf_581_clk;
 wire clknet_leaf_578_clk;
 wire clknet_leaf_572_clk;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire clknet_leaf_570_clk;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire clknet_leaf_569_clk;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire clknet_leaf_562_clk;
 wire clknet_leaf_561_clk;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire clknet_leaf_557_clk;
 wire clknet_leaf_546_clk;
 wire _01457_;
 wire _01458_;
 wire clknet_leaf_545_clk;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire clknet_leaf_536_clk;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire clknet_leaf_534_clk;
 wire clknet_leaf_533_clk;
 wire clknet_leaf_530_clk;
 wire _01484_;
 wire _01485_;
 wire clknet_leaf_528_clk;
 wire _01487_;
 wire _01488_;
 wire clknet_leaf_526_clk;
 wire _01490_;
 wire _01491_;
 wire clknet_leaf_516_clk;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire clknet_leaf_515_clk;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire clknet_leaf_513_clk;
 wire _01514_;
 wire _01515_;
 wire clknet_leaf_509_clk;
 wire clknet_leaf_507_clk;
 wire _01518_;
 wire clknet_leaf_505_clk;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire clknet_leaf_502_clk;
 wire clknet_leaf_497_clk;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire clknet_leaf_496_clk;
 wire clknet_leaf_494_clk;
 wire clknet_leaf_493_clk;
 wire _01539_;
 wire _01540_;
 wire clknet_leaf_492_clk;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire clknet_leaf_491_clk;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire clknet_leaf_488_clk;
 wire clknet_leaf_486_clk;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire clknet_leaf_484_clk;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire clknet_leaf_481_clk;
 wire _01582_;
 wire _01583_;
 wire clknet_leaf_473_clk;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire clknet_leaf_469_clk;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire clknet_leaf_468_clk;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire clknet_leaf_459_clk;
 wire clknet_leaf_458_clk;
 wire clknet_leaf_457_clk;
 wire clknet_leaf_456_clk;
 wire clknet_leaf_454_clk;
 wire _01609_;
 wire _01610_;
 wire clknet_leaf_452_clk;
 wire clknet_leaf_449_clk;
 wire _01613_;
 wire _01614_;
 wire clknet_leaf_448_clk;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire clknet_leaf_446_clk;
 wire clknet_leaf_442_clk;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire clknet_leaf_441_clk;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire clknet_leaf_438_clk;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire clknet_leaf_436_clk;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire clknet_leaf_432_clk;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire clknet_leaf_427_clk;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire clknet_leaf_425_clk;
 wire _01685_;
 wire _01686_;
 wire clknet_leaf_424_clk;
 wire clknet_leaf_423_clk;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire clknet_leaf_421_clk;
 wire _01699_;
 wire clknet_leaf_419_clk;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire clknet_leaf_418_clk;
 wire clknet_leaf_413_clk;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire clknet_leaf_411_clk;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire clknet_leaf_408_clk;
 wire _01757_;
 wire _01758_;
 wire clknet_leaf_404_clk;
 wire clknet_leaf_403_clk;
 wire clknet_leaf_396_clk;
 wire _01762_;
 wire clknet_leaf_394_clk;
 wire _01764_;
 wire _01765_;
 wire clknet_leaf_393_clk;
 wire _01767_;
 wire _01768_;
 wire clknet_leaf_390_clk;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire clknet_leaf_383_clk;
 wire clknet_leaf_380_clk;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire clknet_leaf_375_clk;
 wire _01811_;
 wire clknet_leaf_374_clk;
 wire clknet_leaf_372_clk;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire clknet_leaf_370_clk;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire clknet_leaf_369_clk;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire clknet_leaf_366_clk;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire clknet_leaf_365_clk;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire clknet_leaf_358_clk;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire clknet_leaf_349_clk;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire clknet_leaf_348_clk;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire clknet_leaf_333_clk;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire clknet_leaf_330_clk;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire clknet_leaf_328_clk;
 wire clknet_leaf_326_clk;
 wire clknet_leaf_324_clk;
 wire _02049_;
 wire _02050_;
 wire clknet_leaf_319_clk;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire clknet_leaf_316_clk;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire clknet_leaf_315_clk;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire clknet_leaf_313_clk;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire clknet_leaf_310_clk;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_307_clk;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_294_clk;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_284_clk;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_282_clk;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire clknet_leaf_280_clk;
 wire _02896_;
 wire clknet_leaf_277_clk;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire clknet_leaf_276_clk;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_270_clk;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_267_clk;
 wire _02918_;
 wire _02919_;
 wire clknet_leaf_264_clk;
 wire _02921_;
 wire _02922_;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_253_clk;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire clknet_leaf_246_clk;
 wire _02929_;
 wire clknet_leaf_238_clk;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire clknet_leaf_231_clk;
 wire _02936_;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_228_clk;
 wire _02939_;
 wire clknet_leaf_224_clk;
 wire _02941_;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_220_clk;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire clknet_leaf_205_clk;
 wire _02948_;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_198_clk;
 wire _02951_;
 wire _02952_;
 wire clknet_leaf_195_clk;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_193_clk;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire clknet_leaf_192_clk;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_187_clk;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire clknet_leaf_185_clk;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_175_clk;
 wire _03068_;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_173_clk;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire clknet_leaf_172_clk;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire clknet_leaf_171_clk;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire clknet_leaf_170_clk;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_163_clk;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire clknet_leaf_161_clk;
 wire _03112_;
 wire _03113_;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_153_clk;
 wire _03116_;
 wire clknet_leaf_150_clk;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire clknet_leaf_145_clk;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire clknet_leaf_143_clk;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire clknet_leaf_141_clk;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_137_clk;
 wire _03200_;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_134_clk;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire clknet_leaf_131_clk;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_126_clk;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire clknet_leaf_125_clk;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire clknet_leaf_121_clk;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire clknet_leaf_118_clk;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire clknet_leaf_117_clk;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire clknet_leaf_116_clk;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_112_clk;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_14_clk;
 wire net478;
 wire _04018_;
 wire _04019_;
 wire net527;
 wire _04021_;
 wire clknet_leaf_11_clk;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire clknet_leaf_6_clk;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire clknet_leaf_0_clk;
 wire net529;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire clknet_leaf_12_clk;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire net528;
 wire _04068_;
 wire _04069_;
 wire clknet_leaf_3_clk;
 wire net516;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire clknet_leaf_2_clk;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire net548;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire net522;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire net526;
 wire _04105_;
 wire _04106_;
 wire net520;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire net519;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire net518;
 wire net551;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire net544;
 wire net541;
 wire _04155_;
 wire net525;
 wire net537;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire net540;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire net515;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire net521;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire net514;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire net534;
 wire net533;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire net523;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire net524;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire net511;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire net539;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire net536;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire net508;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire net507;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire net535;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire net530;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire net538;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire net506;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire net505;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire net532;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire net512;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire net531;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire net504;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire net550;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire net503;
 wire _04499_;
 wire _04500_;
 wire net502;
 wire net549;
 wire net501;
 wire net495;
 wire _04505_;
 wire net494;
 wire _04507_;
 wire net493;
 wire net492;
 wire _04510_;
 wire _04511_;
 wire net491;
 wire _04513_;
 wire _04514_;
 wire net496;
 wire net498;
 wire _04517_;
 wire _04518_;
 wire net499;
 wire net500;
 wire _04521_;
 wire _04522_;
 wire net547;
 wire _04524_;
 wire net517;
 wire _04526_;
 wire net488;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire net477;
 wire net482;
 wire _04537_;
 wire clknet_leaf_26_clk;
 wire _04539_;
 wire net497;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire clknet_leaf_27_clk;
 wire _04554_;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_42_clk;
 wire _04557_;
 wire clknet_leaf_56_clk;
 wire _04559_;
 wire net546;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire clknet_leaf_58_clk;
 wire net487;
 wire _04575_;
 wire clknet_leaf_60_clk;
 wire _04577_;
 wire clknet_leaf_64_clk;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire net485;
 wire clknet_leaf_65_clk;
 wire _04593_;
 wire clknet_leaf_67_clk;
 wire _04595_;
 wire clknet_leaf_68_clk;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire clknet_leaf_73_clk;
 wire _04611_;
 wire clknet_leaf_74_clk;
 wire _04613_;
 wire clknet_leaf_75_clk;
 wire _04615_;
 wire clknet_leaf_76_clk;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire clknet_leaf_13_clk;
 wire _04628_;
 wire net481;
 wire _04630_;
 wire clknet_leaf_78_clk;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire clknet_leaf_25_clk;
 wire _04643_;
 wire _04645_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04658_;
 wire _04660_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04671_;
 wire _04680_;
 wire _04682_;
 wire _04688_;
 wire _04691_;
 wire _04692_;
 wire _04695_;
 wire _04700_;
 wire _04704_;
 wire _04709_;
 wire _04711_;
 wire _04713_;
 wire _04714_;
 wire _04718_;
 wire _04720_;
 wire _04723_;
 wire _04725_;
 wire _04728_;
 wire _04731_;
 wire _04733_;
 wire _04735_;
 wire _04737_;
 wire _04738_;
 wire _04741_;
 wire _04743_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04755_;
 wire _04757_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04770_;
 wire _04772_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04786_;
 wire _04788_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04802_;
 wire _04804_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04817_;
 wire _04819_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04833_;
 wire _04835_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04850_;
 wire _04852_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04864_;
 wire _04873_;
 wire _04875_;
 wire _04881_;
 wire net65;
 wire _04884_;
 wire net64;
 wire net63;
 wire _04887_;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire _04892_;
 wire _04893_;
 wire net58;
 wire net57;
 wire net56;
 wire _04897_;
 wire _04898_;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire _04903_;
 wire net51;
 wire _04905_;
 wire net50;
 wire _04907_;
 wire net49;
 wire net48;
 wire net47;
 wire _04911_;
 wire net46;
 wire _04913_;
 wire net45;
 wire net44;
 wire _04916_;
 wire net43;
 wire _04918_;
 wire _04919_;
 wire net42;
 wire net41;
 wire _04922_;
 wire _04923_;
 wire net40;
 wire net39;
 wire _04926_;
 wire _04927_;
 wire net38;
 wire _04929_;
 wire net37;
 wire _04931_;
 wire net36;
 wire _04933_;
 wire _04934_;
 wire net35;
 wire net34;
 wire _04937_;
 wire net33;
 wire _04939_;
 wire net32;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire net31;
 wire net30;
 wire _04953_;
 wire net29;
 wire _04955_;
 wire net28;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire net27;
 wire net26;
 wire _04969_;
 wire net25;
 wire _04971_;
 wire net24;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire net23;
 wire _04984_;
 wire net22;
 wire _04986_;
 wire net21;
 wire _04988_;
 wire net20;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire net19;
 wire _05000_;
 wire net18;
 wire _05002_;
 wire net17;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire net16;
 wire _05014_;
 wire net15;
 wire _05016_;
 wire net14;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire net13;
 wire _05029_;
 wire net12;
 wire _05031_;
 wire net11;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire net10;
 wire net9;
 wire _05045_;
 wire net8;
 wire _05047_;
 wire net7;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire net6;
 wire net5;
 wire _05063_;
 wire net4;
 wire _05065_;
 wire net3;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire net2;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire net1;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_688_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_681_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_465_clk;
 wire clknet_leaf_430_clk;
 wire clknet_leaf_385_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_360_clk;
 wire clknet_leaf_351_clk;
 wire clknet_leaf_334_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_237_clk;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire \dp.ISRmux.d0[10] ;
 wire \dp.ISRmux.d0[11] ;
 wire \dp.ISRmux.d0[12] ;
 wire \dp.ISRmux.d0[13] ;
 wire \dp.ISRmux.d0[14] ;
 wire \dp.ISRmux.d0[15] ;
 wire \dp.ISRmux.d0[16] ;
 wire \dp.ISRmux.d0[17] ;
 wire \dp.ISRmux.d0[18] ;
 wire \dp.ISRmux.d0[19] ;
 wire \dp.ISRmux.d0[20] ;
 wire \dp.ISRmux.d0[21] ;
 wire \dp.ISRmux.d0[22] ;
 wire \dp.ISRmux.d0[23] ;
 wire \dp.ISRmux.d0[24] ;
 wire \dp.ISRmux.d0[25] ;
 wire \dp.ISRmux.d0[26] ;
 wire \dp.ISRmux.d0[27] ;
 wire \dp.ISRmux.d0[28] ;
 wire \dp.ISRmux.d0[29] ;
 wire \dp.ISRmux.d0[2] ;
 wire \dp.ISRmux.d0[30] ;
 wire \dp.ISRmux.d0[31] ;
 wire \dp.ISRmux.d0[3] ;
 wire \dp.ISRmux.d0[4] ;
 wire \dp.ISRmux.d0[5] ;
 wire \dp.ISRmux.d0[6] ;
 wire \dp.ISRmux.d0[7] ;
 wire \dp.ISRmux.d0[8] ;
 wire \dp.ISRmux.d0[9] ;
 wire \dp.rf.rf[0][0] ;
 wire \dp.rf.rf[0][10] ;
 wire \dp.rf.rf[0][11] ;
 wire \dp.rf.rf[0][12] ;
 wire \dp.rf.rf[0][13] ;
 wire \dp.rf.rf[0][14] ;
 wire \dp.rf.rf[0][15] ;
 wire \dp.rf.rf[0][16] ;
 wire \dp.rf.rf[0][17] ;
 wire \dp.rf.rf[0][18] ;
 wire \dp.rf.rf[0][19] ;
 wire \dp.rf.rf[0][1] ;
 wire \dp.rf.rf[0][20] ;
 wire \dp.rf.rf[0][21] ;
 wire \dp.rf.rf[0][22] ;
 wire \dp.rf.rf[0][23] ;
 wire \dp.rf.rf[0][24] ;
 wire \dp.rf.rf[0][25] ;
 wire \dp.rf.rf[0][26] ;
 wire \dp.rf.rf[0][27] ;
 wire \dp.rf.rf[0][28] ;
 wire \dp.rf.rf[0][29] ;
 wire \dp.rf.rf[0][2] ;
 wire \dp.rf.rf[0][30] ;
 wire \dp.rf.rf[0][31] ;
 wire \dp.rf.rf[0][3] ;
 wire \dp.rf.rf[0][4] ;
 wire \dp.rf.rf[0][5] ;
 wire \dp.rf.rf[0][6] ;
 wire \dp.rf.rf[0][7] ;
 wire \dp.rf.rf[0][8] ;
 wire \dp.rf.rf[0][9] ;
 wire \dp.rf.rf[10][0] ;
 wire \dp.rf.rf[10][10] ;
 wire \dp.rf.rf[10][11] ;
 wire \dp.rf.rf[10][12] ;
 wire \dp.rf.rf[10][13] ;
 wire \dp.rf.rf[10][14] ;
 wire \dp.rf.rf[10][15] ;
 wire \dp.rf.rf[10][16] ;
 wire \dp.rf.rf[10][17] ;
 wire \dp.rf.rf[10][18] ;
 wire \dp.rf.rf[10][19] ;
 wire \dp.rf.rf[10][1] ;
 wire \dp.rf.rf[10][20] ;
 wire \dp.rf.rf[10][21] ;
 wire \dp.rf.rf[10][22] ;
 wire \dp.rf.rf[10][23] ;
 wire \dp.rf.rf[10][24] ;
 wire \dp.rf.rf[10][25] ;
 wire \dp.rf.rf[10][26] ;
 wire \dp.rf.rf[10][27] ;
 wire \dp.rf.rf[10][28] ;
 wire \dp.rf.rf[10][29] ;
 wire \dp.rf.rf[10][2] ;
 wire \dp.rf.rf[10][30] ;
 wire \dp.rf.rf[10][31] ;
 wire \dp.rf.rf[10][3] ;
 wire \dp.rf.rf[10][4] ;
 wire \dp.rf.rf[10][5] ;
 wire \dp.rf.rf[10][6] ;
 wire \dp.rf.rf[10][7] ;
 wire \dp.rf.rf[10][8] ;
 wire \dp.rf.rf[10][9] ;
 wire \dp.rf.rf[11][0] ;
 wire \dp.rf.rf[11][10] ;
 wire \dp.rf.rf[11][11] ;
 wire \dp.rf.rf[11][12] ;
 wire \dp.rf.rf[11][13] ;
 wire \dp.rf.rf[11][14] ;
 wire \dp.rf.rf[11][15] ;
 wire \dp.rf.rf[11][16] ;
 wire \dp.rf.rf[11][17] ;
 wire \dp.rf.rf[11][18] ;
 wire \dp.rf.rf[11][19] ;
 wire \dp.rf.rf[11][1] ;
 wire \dp.rf.rf[11][20] ;
 wire \dp.rf.rf[11][21] ;
 wire \dp.rf.rf[11][22] ;
 wire \dp.rf.rf[11][23] ;
 wire \dp.rf.rf[11][24] ;
 wire \dp.rf.rf[11][25] ;
 wire \dp.rf.rf[11][26] ;
 wire \dp.rf.rf[11][27] ;
 wire \dp.rf.rf[11][28] ;
 wire \dp.rf.rf[11][29] ;
 wire \dp.rf.rf[11][2] ;
 wire \dp.rf.rf[11][30] ;
 wire \dp.rf.rf[11][31] ;
 wire \dp.rf.rf[11][3] ;
 wire \dp.rf.rf[11][4] ;
 wire \dp.rf.rf[11][5] ;
 wire \dp.rf.rf[11][6] ;
 wire \dp.rf.rf[11][7] ;
 wire \dp.rf.rf[11][8] ;
 wire \dp.rf.rf[11][9] ;
 wire \dp.rf.rf[12][0] ;
 wire \dp.rf.rf[12][10] ;
 wire \dp.rf.rf[12][11] ;
 wire \dp.rf.rf[12][12] ;
 wire \dp.rf.rf[12][13] ;
 wire \dp.rf.rf[12][14] ;
 wire \dp.rf.rf[12][15] ;
 wire \dp.rf.rf[12][16] ;
 wire \dp.rf.rf[12][17] ;
 wire \dp.rf.rf[12][18] ;
 wire \dp.rf.rf[12][19] ;
 wire \dp.rf.rf[12][1] ;
 wire \dp.rf.rf[12][20] ;
 wire \dp.rf.rf[12][21] ;
 wire \dp.rf.rf[12][22] ;
 wire \dp.rf.rf[12][23] ;
 wire \dp.rf.rf[12][24] ;
 wire \dp.rf.rf[12][25] ;
 wire \dp.rf.rf[12][26] ;
 wire \dp.rf.rf[12][27] ;
 wire \dp.rf.rf[12][28] ;
 wire \dp.rf.rf[12][29] ;
 wire \dp.rf.rf[12][2] ;
 wire \dp.rf.rf[12][30] ;
 wire \dp.rf.rf[12][31] ;
 wire \dp.rf.rf[12][3] ;
 wire \dp.rf.rf[12][4] ;
 wire \dp.rf.rf[12][5] ;
 wire \dp.rf.rf[12][6] ;
 wire \dp.rf.rf[12][7] ;
 wire \dp.rf.rf[12][8] ;
 wire \dp.rf.rf[12][9] ;
 wire \dp.rf.rf[13][0] ;
 wire \dp.rf.rf[13][10] ;
 wire \dp.rf.rf[13][11] ;
 wire \dp.rf.rf[13][12] ;
 wire \dp.rf.rf[13][13] ;
 wire \dp.rf.rf[13][14] ;
 wire \dp.rf.rf[13][15] ;
 wire \dp.rf.rf[13][16] ;
 wire \dp.rf.rf[13][17] ;
 wire \dp.rf.rf[13][18] ;
 wire \dp.rf.rf[13][19] ;
 wire \dp.rf.rf[13][1] ;
 wire \dp.rf.rf[13][20] ;
 wire \dp.rf.rf[13][21] ;
 wire \dp.rf.rf[13][22] ;
 wire \dp.rf.rf[13][23] ;
 wire \dp.rf.rf[13][24] ;
 wire \dp.rf.rf[13][25] ;
 wire \dp.rf.rf[13][26] ;
 wire \dp.rf.rf[13][27] ;
 wire \dp.rf.rf[13][28] ;
 wire \dp.rf.rf[13][29] ;
 wire \dp.rf.rf[13][2] ;
 wire \dp.rf.rf[13][30] ;
 wire \dp.rf.rf[13][31] ;
 wire \dp.rf.rf[13][3] ;
 wire \dp.rf.rf[13][4] ;
 wire \dp.rf.rf[13][5] ;
 wire \dp.rf.rf[13][6] ;
 wire \dp.rf.rf[13][7] ;
 wire \dp.rf.rf[13][8] ;
 wire \dp.rf.rf[13][9] ;
 wire \dp.rf.rf[14][0] ;
 wire \dp.rf.rf[14][10] ;
 wire \dp.rf.rf[14][11] ;
 wire \dp.rf.rf[14][12] ;
 wire \dp.rf.rf[14][13] ;
 wire \dp.rf.rf[14][14] ;
 wire \dp.rf.rf[14][15] ;
 wire \dp.rf.rf[14][16] ;
 wire \dp.rf.rf[14][17] ;
 wire \dp.rf.rf[14][18] ;
 wire \dp.rf.rf[14][19] ;
 wire \dp.rf.rf[14][1] ;
 wire \dp.rf.rf[14][20] ;
 wire \dp.rf.rf[14][21] ;
 wire \dp.rf.rf[14][22] ;
 wire \dp.rf.rf[14][23] ;
 wire \dp.rf.rf[14][24] ;
 wire \dp.rf.rf[14][25] ;
 wire \dp.rf.rf[14][26] ;
 wire \dp.rf.rf[14][27] ;
 wire \dp.rf.rf[14][28] ;
 wire \dp.rf.rf[14][29] ;
 wire \dp.rf.rf[14][2] ;
 wire \dp.rf.rf[14][30] ;
 wire \dp.rf.rf[14][31] ;
 wire \dp.rf.rf[14][3] ;
 wire \dp.rf.rf[14][4] ;
 wire \dp.rf.rf[14][5] ;
 wire \dp.rf.rf[14][6] ;
 wire \dp.rf.rf[14][7] ;
 wire \dp.rf.rf[14][8] ;
 wire \dp.rf.rf[14][9] ;
 wire \dp.rf.rf[15][0] ;
 wire \dp.rf.rf[15][10] ;
 wire \dp.rf.rf[15][11] ;
 wire \dp.rf.rf[15][12] ;
 wire \dp.rf.rf[15][13] ;
 wire \dp.rf.rf[15][14] ;
 wire \dp.rf.rf[15][15] ;
 wire \dp.rf.rf[15][16] ;
 wire \dp.rf.rf[15][17] ;
 wire \dp.rf.rf[15][18] ;
 wire \dp.rf.rf[15][19] ;
 wire \dp.rf.rf[15][1] ;
 wire \dp.rf.rf[15][20] ;
 wire \dp.rf.rf[15][21] ;
 wire \dp.rf.rf[15][22] ;
 wire \dp.rf.rf[15][23] ;
 wire \dp.rf.rf[15][24] ;
 wire \dp.rf.rf[15][25] ;
 wire \dp.rf.rf[15][26] ;
 wire \dp.rf.rf[15][27] ;
 wire \dp.rf.rf[15][28] ;
 wire \dp.rf.rf[15][29] ;
 wire \dp.rf.rf[15][2] ;
 wire \dp.rf.rf[15][30] ;
 wire \dp.rf.rf[15][31] ;
 wire \dp.rf.rf[15][3] ;
 wire \dp.rf.rf[15][4] ;
 wire \dp.rf.rf[15][5] ;
 wire \dp.rf.rf[15][6] ;
 wire \dp.rf.rf[15][7] ;
 wire \dp.rf.rf[15][8] ;
 wire \dp.rf.rf[15][9] ;
 wire \dp.rf.rf[16][0] ;
 wire \dp.rf.rf[16][10] ;
 wire \dp.rf.rf[16][11] ;
 wire \dp.rf.rf[16][12] ;
 wire \dp.rf.rf[16][13] ;
 wire \dp.rf.rf[16][14] ;
 wire \dp.rf.rf[16][15] ;
 wire \dp.rf.rf[16][16] ;
 wire \dp.rf.rf[16][17] ;
 wire \dp.rf.rf[16][18] ;
 wire \dp.rf.rf[16][19] ;
 wire \dp.rf.rf[16][1] ;
 wire \dp.rf.rf[16][20] ;
 wire \dp.rf.rf[16][21] ;
 wire \dp.rf.rf[16][22] ;
 wire \dp.rf.rf[16][23] ;
 wire \dp.rf.rf[16][24] ;
 wire \dp.rf.rf[16][25] ;
 wire \dp.rf.rf[16][26] ;
 wire \dp.rf.rf[16][27] ;
 wire \dp.rf.rf[16][28] ;
 wire \dp.rf.rf[16][29] ;
 wire \dp.rf.rf[16][2] ;
 wire \dp.rf.rf[16][30] ;
 wire \dp.rf.rf[16][31] ;
 wire \dp.rf.rf[16][3] ;
 wire \dp.rf.rf[16][4] ;
 wire \dp.rf.rf[16][5] ;
 wire \dp.rf.rf[16][6] ;
 wire \dp.rf.rf[16][7] ;
 wire \dp.rf.rf[16][8] ;
 wire \dp.rf.rf[16][9] ;
 wire \dp.rf.rf[17][0] ;
 wire \dp.rf.rf[17][10] ;
 wire \dp.rf.rf[17][11] ;
 wire \dp.rf.rf[17][12] ;
 wire \dp.rf.rf[17][13] ;
 wire \dp.rf.rf[17][14] ;
 wire \dp.rf.rf[17][15] ;
 wire \dp.rf.rf[17][16] ;
 wire \dp.rf.rf[17][17] ;
 wire \dp.rf.rf[17][18] ;
 wire \dp.rf.rf[17][19] ;
 wire \dp.rf.rf[17][1] ;
 wire \dp.rf.rf[17][20] ;
 wire \dp.rf.rf[17][21] ;
 wire \dp.rf.rf[17][22] ;
 wire \dp.rf.rf[17][23] ;
 wire \dp.rf.rf[17][24] ;
 wire \dp.rf.rf[17][25] ;
 wire \dp.rf.rf[17][26] ;
 wire \dp.rf.rf[17][27] ;
 wire \dp.rf.rf[17][28] ;
 wire \dp.rf.rf[17][29] ;
 wire \dp.rf.rf[17][2] ;
 wire \dp.rf.rf[17][30] ;
 wire \dp.rf.rf[17][31] ;
 wire \dp.rf.rf[17][3] ;
 wire \dp.rf.rf[17][4] ;
 wire \dp.rf.rf[17][5] ;
 wire \dp.rf.rf[17][6] ;
 wire \dp.rf.rf[17][7] ;
 wire \dp.rf.rf[17][8] ;
 wire \dp.rf.rf[17][9] ;
 wire \dp.rf.rf[18][0] ;
 wire \dp.rf.rf[18][10] ;
 wire \dp.rf.rf[18][11] ;
 wire \dp.rf.rf[18][12] ;
 wire \dp.rf.rf[18][13] ;
 wire \dp.rf.rf[18][14] ;
 wire \dp.rf.rf[18][15] ;
 wire \dp.rf.rf[18][16] ;
 wire \dp.rf.rf[18][17] ;
 wire \dp.rf.rf[18][18] ;
 wire \dp.rf.rf[18][19] ;
 wire \dp.rf.rf[18][1] ;
 wire \dp.rf.rf[18][20] ;
 wire \dp.rf.rf[18][21] ;
 wire \dp.rf.rf[18][22] ;
 wire \dp.rf.rf[18][23] ;
 wire \dp.rf.rf[18][24] ;
 wire \dp.rf.rf[18][25] ;
 wire \dp.rf.rf[18][26] ;
 wire \dp.rf.rf[18][27] ;
 wire \dp.rf.rf[18][28] ;
 wire \dp.rf.rf[18][29] ;
 wire \dp.rf.rf[18][2] ;
 wire \dp.rf.rf[18][30] ;
 wire \dp.rf.rf[18][31] ;
 wire \dp.rf.rf[18][3] ;
 wire \dp.rf.rf[18][4] ;
 wire \dp.rf.rf[18][5] ;
 wire \dp.rf.rf[18][6] ;
 wire \dp.rf.rf[18][7] ;
 wire \dp.rf.rf[18][8] ;
 wire \dp.rf.rf[18][9] ;
 wire \dp.rf.rf[19][0] ;
 wire \dp.rf.rf[19][10] ;
 wire \dp.rf.rf[19][11] ;
 wire \dp.rf.rf[19][12] ;
 wire \dp.rf.rf[19][13] ;
 wire \dp.rf.rf[19][14] ;
 wire \dp.rf.rf[19][15] ;
 wire \dp.rf.rf[19][16] ;
 wire \dp.rf.rf[19][17] ;
 wire \dp.rf.rf[19][18] ;
 wire \dp.rf.rf[19][19] ;
 wire \dp.rf.rf[19][1] ;
 wire \dp.rf.rf[19][20] ;
 wire \dp.rf.rf[19][21] ;
 wire \dp.rf.rf[19][22] ;
 wire \dp.rf.rf[19][23] ;
 wire \dp.rf.rf[19][24] ;
 wire \dp.rf.rf[19][25] ;
 wire \dp.rf.rf[19][26] ;
 wire \dp.rf.rf[19][27] ;
 wire \dp.rf.rf[19][28] ;
 wire \dp.rf.rf[19][29] ;
 wire \dp.rf.rf[19][2] ;
 wire \dp.rf.rf[19][30] ;
 wire \dp.rf.rf[19][31] ;
 wire \dp.rf.rf[19][3] ;
 wire \dp.rf.rf[19][4] ;
 wire \dp.rf.rf[19][5] ;
 wire \dp.rf.rf[19][6] ;
 wire \dp.rf.rf[19][7] ;
 wire \dp.rf.rf[19][8] ;
 wire \dp.rf.rf[19][9] ;
 wire \dp.rf.rf[1][0] ;
 wire \dp.rf.rf[1][10] ;
 wire \dp.rf.rf[1][11] ;
 wire \dp.rf.rf[1][12] ;
 wire \dp.rf.rf[1][13] ;
 wire \dp.rf.rf[1][14] ;
 wire \dp.rf.rf[1][15] ;
 wire \dp.rf.rf[1][16] ;
 wire \dp.rf.rf[1][17] ;
 wire \dp.rf.rf[1][18] ;
 wire \dp.rf.rf[1][19] ;
 wire \dp.rf.rf[1][1] ;
 wire \dp.rf.rf[1][20] ;
 wire \dp.rf.rf[1][21] ;
 wire \dp.rf.rf[1][22] ;
 wire \dp.rf.rf[1][23] ;
 wire \dp.rf.rf[1][24] ;
 wire \dp.rf.rf[1][25] ;
 wire \dp.rf.rf[1][26] ;
 wire \dp.rf.rf[1][27] ;
 wire \dp.rf.rf[1][28] ;
 wire \dp.rf.rf[1][29] ;
 wire \dp.rf.rf[1][2] ;
 wire \dp.rf.rf[1][30] ;
 wire \dp.rf.rf[1][31] ;
 wire \dp.rf.rf[1][3] ;
 wire \dp.rf.rf[1][4] ;
 wire \dp.rf.rf[1][5] ;
 wire \dp.rf.rf[1][6] ;
 wire \dp.rf.rf[1][7] ;
 wire \dp.rf.rf[1][8] ;
 wire \dp.rf.rf[1][9] ;
 wire \dp.rf.rf[20][0] ;
 wire \dp.rf.rf[20][10] ;
 wire \dp.rf.rf[20][11] ;
 wire \dp.rf.rf[20][12] ;
 wire \dp.rf.rf[20][13] ;
 wire \dp.rf.rf[20][14] ;
 wire \dp.rf.rf[20][15] ;
 wire \dp.rf.rf[20][16] ;
 wire \dp.rf.rf[20][17] ;
 wire \dp.rf.rf[20][18] ;
 wire \dp.rf.rf[20][19] ;
 wire \dp.rf.rf[20][1] ;
 wire \dp.rf.rf[20][20] ;
 wire \dp.rf.rf[20][21] ;
 wire \dp.rf.rf[20][22] ;
 wire \dp.rf.rf[20][23] ;
 wire \dp.rf.rf[20][24] ;
 wire \dp.rf.rf[20][25] ;
 wire \dp.rf.rf[20][26] ;
 wire \dp.rf.rf[20][27] ;
 wire \dp.rf.rf[20][28] ;
 wire \dp.rf.rf[20][29] ;
 wire \dp.rf.rf[20][2] ;
 wire \dp.rf.rf[20][30] ;
 wire \dp.rf.rf[20][31] ;
 wire \dp.rf.rf[20][3] ;
 wire \dp.rf.rf[20][4] ;
 wire \dp.rf.rf[20][5] ;
 wire \dp.rf.rf[20][6] ;
 wire \dp.rf.rf[20][7] ;
 wire \dp.rf.rf[20][8] ;
 wire \dp.rf.rf[20][9] ;
 wire \dp.rf.rf[21][0] ;
 wire \dp.rf.rf[21][10] ;
 wire \dp.rf.rf[21][11] ;
 wire \dp.rf.rf[21][12] ;
 wire \dp.rf.rf[21][13] ;
 wire \dp.rf.rf[21][14] ;
 wire \dp.rf.rf[21][15] ;
 wire \dp.rf.rf[21][16] ;
 wire \dp.rf.rf[21][17] ;
 wire \dp.rf.rf[21][18] ;
 wire \dp.rf.rf[21][19] ;
 wire \dp.rf.rf[21][1] ;
 wire \dp.rf.rf[21][20] ;
 wire \dp.rf.rf[21][21] ;
 wire \dp.rf.rf[21][22] ;
 wire \dp.rf.rf[21][23] ;
 wire \dp.rf.rf[21][24] ;
 wire \dp.rf.rf[21][25] ;
 wire \dp.rf.rf[21][26] ;
 wire \dp.rf.rf[21][27] ;
 wire \dp.rf.rf[21][28] ;
 wire \dp.rf.rf[21][29] ;
 wire \dp.rf.rf[21][2] ;
 wire \dp.rf.rf[21][30] ;
 wire \dp.rf.rf[21][31] ;
 wire \dp.rf.rf[21][3] ;
 wire \dp.rf.rf[21][4] ;
 wire \dp.rf.rf[21][5] ;
 wire \dp.rf.rf[21][6] ;
 wire \dp.rf.rf[21][7] ;
 wire \dp.rf.rf[21][8] ;
 wire \dp.rf.rf[21][9] ;
 wire \dp.rf.rf[22][0] ;
 wire \dp.rf.rf[22][10] ;
 wire \dp.rf.rf[22][11] ;
 wire \dp.rf.rf[22][12] ;
 wire \dp.rf.rf[22][13] ;
 wire \dp.rf.rf[22][14] ;
 wire \dp.rf.rf[22][15] ;
 wire \dp.rf.rf[22][16] ;
 wire \dp.rf.rf[22][17] ;
 wire \dp.rf.rf[22][18] ;
 wire \dp.rf.rf[22][19] ;
 wire \dp.rf.rf[22][1] ;
 wire \dp.rf.rf[22][20] ;
 wire \dp.rf.rf[22][21] ;
 wire \dp.rf.rf[22][22] ;
 wire \dp.rf.rf[22][23] ;
 wire \dp.rf.rf[22][24] ;
 wire \dp.rf.rf[22][25] ;
 wire \dp.rf.rf[22][26] ;
 wire \dp.rf.rf[22][27] ;
 wire \dp.rf.rf[22][28] ;
 wire \dp.rf.rf[22][29] ;
 wire \dp.rf.rf[22][2] ;
 wire \dp.rf.rf[22][30] ;
 wire \dp.rf.rf[22][31] ;
 wire \dp.rf.rf[22][3] ;
 wire \dp.rf.rf[22][4] ;
 wire \dp.rf.rf[22][5] ;
 wire \dp.rf.rf[22][6] ;
 wire \dp.rf.rf[22][7] ;
 wire \dp.rf.rf[22][8] ;
 wire \dp.rf.rf[22][9] ;
 wire \dp.rf.rf[23][0] ;
 wire \dp.rf.rf[23][10] ;
 wire \dp.rf.rf[23][11] ;
 wire \dp.rf.rf[23][12] ;
 wire \dp.rf.rf[23][13] ;
 wire \dp.rf.rf[23][14] ;
 wire \dp.rf.rf[23][15] ;
 wire \dp.rf.rf[23][16] ;
 wire \dp.rf.rf[23][17] ;
 wire \dp.rf.rf[23][18] ;
 wire \dp.rf.rf[23][19] ;
 wire \dp.rf.rf[23][1] ;
 wire \dp.rf.rf[23][20] ;
 wire \dp.rf.rf[23][21] ;
 wire \dp.rf.rf[23][22] ;
 wire \dp.rf.rf[23][23] ;
 wire \dp.rf.rf[23][24] ;
 wire \dp.rf.rf[23][25] ;
 wire \dp.rf.rf[23][26] ;
 wire \dp.rf.rf[23][27] ;
 wire \dp.rf.rf[23][28] ;
 wire \dp.rf.rf[23][29] ;
 wire \dp.rf.rf[23][2] ;
 wire \dp.rf.rf[23][30] ;
 wire \dp.rf.rf[23][31] ;
 wire \dp.rf.rf[23][3] ;
 wire \dp.rf.rf[23][4] ;
 wire \dp.rf.rf[23][5] ;
 wire \dp.rf.rf[23][6] ;
 wire \dp.rf.rf[23][7] ;
 wire \dp.rf.rf[23][8] ;
 wire \dp.rf.rf[23][9] ;
 wire \dp.rf.rf[24][0] ;
 wire \dp.rf.rf[24][10] ;
 wire \dp.rf.rf[24][11] ;
 wire \dp.rf.rf[24][12] ;
 wire \dp.rf.rf[24][13] ;
 wire \dp.rf.rf[24][14] ;
 wire \dp.rf.rf[24][15] ;
 wire \dp.rf.rf[24][16] ;
 wire \dp.rf.rf[24][17] ;
 wire \dp.rf.rf[24][18] ;
 wire \dp.rf.rf[24][19] ;
 wire \dp.rf.rf[24][1] ;
 wire \dp.rf.rf[24][20] ;
 wire \dp.rf.rf[24][21] ;
 wire \dp.rf.rf[24][22] ;
 wire \dp.rf.rf[24][23] ;
 wire \dp.rf.rf[24][24] ;
 wire \dp.rf.rf[24][25] ;
 wire \dp.rf.rf[24][26] ;
 wire \dp.rf.rf[24][27] ;
 wire \dp.rf.rf[24][28] ;
 wire \dp.rf.rf[24][29] ;
 wire \dp.rf.rf[24][2] ;
 wire \dp.rf.rf[24][30] ;
 wire \dp.rf.rf[24][31] ;
 wire \dp.rf.rf[24][3] ;
 wire \dp.rf.rf[24][4] ;
 wire \dp.rf.rf[24][5] ;
 wire \dp.rf.rf[24][6] ;
 wire \dp.rf.rf[24][7] ;
 wire \dp.rf.rf[24][8] ;
 wire \dp.rf.rf[24][9] ;
 wire \dp.rf.rf[25][0] ;
 wire \dp.rf.rf[25][10] ;
 wire \dp.rf.rf[25][11] ;
 wire \dp.rf.rf[25][12] ;
 wire \dp.rf.rf[25][13] ;
 wire \dp.rf.rf[25][14] ;
 wire \dp.rf.rf[25][15] ;
 wire \dp.rf.rf[25][16] ;
 wire \dp.rf.rf[25][17] ;
 wire \dp.rf.rf[25][18] ;
 wire \dp.rf.rf[25][19] ;
 wire \dp.rf.rf[25][1] ;
 wire \dp.rf.rf[25][20] ;
 wire \dp.rf.rf[25][21] ;
 wire \dp.rf.rf[25][22] ;
 wire \dp.rf.rf[25][23] ;
 wire \dp.rf.rf[25][24] ;
 wire \dp.rf.rf[25][25] ;
 wire \dp.rf.rf[25][26] ;
 wire \dp.rf.rf[25][27] ;
 wire \dp.rf.rf[25][28] ;
 wire \dp.rf.rf[25][29] ;
 wire \dp.rf.rf[25][2] ;
 wire \dp.rf.rf[25][30] ;
 wire \dp.rf.rf[25][31] ;
 wire \dp.rf.rf[25][3] ;
 wire \dp.rf.rf[25][4] ;
 wire \dp.rf.rf[25][5] ;
 wire \dp.rf.rf[25][6] ;
 wire \dp.rf.rf[25][7] ;
 wire \dp.rf.rf[25][8] ;
 wire \dp.rf.rf[25][9] ;
 wire \dp.rf.rf[26][0] ;
 wire \dp.rf.rf[26][10] ;
 wire \dp.rf.rf[26][11] ;
 wire \dp.rf.rf[26][12] ;
 wire \dp.rf.rf[26][13] ;
 wire \dp.rf.rf[26][14] ;
 wire \dp.rf.rf[26][15] ;
 wire \dp.rf.rf[26][16] ;
 wire \dp.rf.rf[26][17] ;
 wire \dp.rf.rf[26][18] ;
 wire \dp.rf.rf[26][19] ;
 wire \dp.rf.rf[26][1] ;
 wire \dp.rf.rf[26][20] ;
 wire \dp.rf.rf[26][21] ;
 wire \dp.rf.rf[26][22] ;
 wire \dp.rf.rf[26][23] ;
 wire \dp.rf.rf[26][24] ;
 wire \dp.rf.rf[26][25] ;
 wire \dp.rf.rf[26][26] ;
 wire \dp.rf.rf[26][27] ;
 wire \dp.rf.rf[26][28] ;
 wire \dp.rf.rf[26][29] ;
 wire \dp.rf.rf[26][2] ;
 wire \dp.rf.rf[26][30] ;
 wire \dp.rf.rf[26][31] ;
 wire \dp.rf.rf[26][3] ;
 wire \dp.rf.rf[26][4] ;
 wire \dp.rf.rf[26][5] ;
 wire \dp.rf.rf[26][6] ;
 wire \dp.rf.rf[26][7] ;
 wire \dp.rf.rf[26][8] ;
 wire \dp.rf.rf[26][9] ;
 wire \dp.rf.rf[27][0] ;
 wire \dp.rf.rf[27][10] ;
 wire \dp.rf.rf[27][11] ;
 wire \dp.rf.rf[27][12] ;
 wire \dp.rf.rf[27][13] ;
 wire \dp.rf.rf[27][14] ;
 wire \dp.rf.rf[27][15] ;
 wire \dp.rf.rf[27][16] ;
 wire \dp.rf.rf[27][17] ;
 wire \dp.rf.rf[27][18] ;
 wire \dp.rf.rf[27][19] ;
 wire \dp.rf.rf[27][1] ;
 wire \dp.rf.rf[27][20] ;
 wire \dp.rf.rf[27][21] ;
 wire \dp.rf.rf[27][22] ;
 wire \dp.rf.rf[27][23] ;
 wire \dp.rf.rf[27][24] ;
 wire \dp.rf.rf[27][25] ;
 wire \dp.rf.rf[27][26] ;
 wire \dp.rf.rf[27][27] ;
 wire \dp.rf.rf[27][28] ;
 wire \dp.rf.rf[27][29] ;
 wire \dp.rf.rf[27][2] ;
 wire \dp.rf.rf[27][30] ;
 wire \dp.rf.rf[27][31] ;
 wire \dp.rf.rf[27][3] ;
 wire \dp.rf.rf[27][4] ;
 wire \dp.rf.rf[27][5] ;
 wire \dp.rf.rf[27][6] ;
 wire \dp.rf.rf[27][7] ;
 wire \dp.rf.rf[27][8] ;
 wire \dp.rf.rf[27][9] ;
 wire \dp.rf.rf[28][0] ;
 wire \dp.rf.rf[28][10] ;
 wire \dp.rf.rf[28][11] ;
 wire \dp.rf.rf[28][12] ;
 wire \dp.rf.rf[28][13] ;
 wire \dp.rf.rf[28][14] ;
 wire \dp.rf.rf[28][15] ;
 wire \dp.rf.rf[28][16] ;
 wire \dp.rf.rf[28][17] ;
 wire \dp.rf.rf[28][18] ;
 wire \dp.rf.rf[28][19] ;
 wire \dp.rf.rf[28][1] ;
 wire \dp.rf.rf[28][20] ;
 wire \dp.rf.rf[28][21] ;
 wire \dp.rf.rf[28][22] ;
 wire \dp.rf.rf[28][23] ;
 wire \dp.rf.rf[28][24] ;
 wire \dp.rf.rf[28][25] ;
 wire \dp.rf.rf[28][26] ;
 wire \dp.rf.rf[28][27] ;
 wire \dp.rf.rf[28][28] ;
 wire \dp.rf.rf[28][29] ;
 wire \dp.rf.rf[28][2] ;
 wire \dp.rf.rf[28][30] ;
 wire \dp.rf.rf[28][31] ;
 wire \dp.rf.rf[28][3] ;
 wire \dp.rf.rf[28][4] ;
 wire \dp.rf.rf[28][5] ;
 wire \dp.rf.rf[28][6] ;
 wire \dp.rf.rf[28][7] ;
 wire \dp.rf.rf[28][8] ;
 wire \dp.rf.rf[28][9] ;
 wire \dp.rf.rf[29][0] ;
 wire \dp.rf.rf[29][10] ;
 wire \dp.rf.rf[29][11] ;
 wire \dp.rf.rf[29][12] ;
 wire \dp.rf.rf[29][13] ;
 wire \dp.rf.rf[29][14] ;
 wire \dp.rf.rf[29][15] ;
 wire \dp.rf.rf[29][16] ;
 wire \dp.rf.rf[29][17] ;
 wire \dp.rf.rf[29][18] ;
 wire \dp.rf.rf[29][19] ;
 wire \dp.rf.rf[29][1] ;
 wire \dp.rf.rf[29][20] ;
 wire \dp.rf.rf[29][21] ;
 wire \dp.rf.rf[29][22] ;
 wire \dp.rf.rf[29][23] ;
 wire \dp.rf.rf[29][24] ;
 wire \dp.rf.rf[29][25] ;
 wire \dp.rf.rf[29][26] ;
 wire \dp.rf.rf[29][27] ;
 wire \dp.rf.rf[29][28] ;
 wire \dp.rf.rf[29][29] ;
 wire \dp.rf.rf[29][2] ;
 wire \dp.rf.rf[29][30] ;
 wire \dp.rf.rf[29][31] ;
 wire \dp.rf.rf[29][3] ;
 wire \dp.rf.rf[29][4] ;
 wire \dp.rf.rf[29][5] ;
 wire \dp.rf.rf[29][6] ;
 wire \dp.rf.rf[29][7] ;
 wire \dp.rf.rf[29][8] ;
 wire \dp.rf.rf[29][9] ;
 wire \dp.rf.rf[2][0] ;
 wire \dp.rf.rf[2][10] ;
 wire \dp.rf.rf[2][11] ;
 wire \dp.rf.rf[2][12] ;
 wire \dp.rf.rf[2][13] ;
 wire \dp.rf.rf[2][14] ;
 wire \dp.rf.rf[2][15] ;
 wire \dp.rf.rf[2][16] ;
 wire \dp.rf.rf[2][17] ;
 wire \dp.rf.rf[2][18] ;
 wire \dp.rf.rf[2][19] ;
 wire \dp.rf.rf[2][1] ;
 wire \dp.rf.rf[2][20] ;
 wire \dp.rf.rf[2][21] ;
 wire \dp.rf.rf[2][22] ;
 wire \dp.rf.rf[2][23] ;
 wire \dp.rf.rf[2][24] ;
 wire \dp.rf.rf[2][25] ;
 wire \dp.rf.rf[2][26] ;
 wire \dp.rf.rf[2][27] ;
 wire \dp.rf.rf[2][28] ;
 wire \dp.rf.rf[2][29] ;
 wire \dp.rf.rf[2][2] ;
 wire \dp.rf.rf[2][30] ;
 wire \dp.rf.rf[2][31] ;
 wire \dp.rf.rf[2][3] ;
 wire \dp.rf.rf[2][4] ;
 wire \dp.rf.rf[2][5] ;
 wire \dp.rf.rf[2][6] ;
 wire \dp.rf.rf[2][7] ;
 wire \dp.rf.rf[2][8] ;
 wire \dp.rf.rf[2][9] ;
 wire \dp.rf.rf[30][0] ;
 wire \dp.rf.rf[30][10] ;
 wire \dp.rf.rf[30][11] ;
 wire \dp.rf.rf[30][12] ;
 wire \dp.rf.rf[30][13] ;
 wire \dp.rf.rf[30][14] ;
 wire \dp.rf.rf[30][15] ;
 wire \dp.rf.rf[30][16] ;
 wire \dp.rf.rf[30][17] ;
 wire \dp.rf.rf[30][18] ;
 wire \dp.rf.rf[30][19] ;
 wire \dp.rf.rf[30][1] ;
 wire \dp.rf.rf[30][20] ;
 wire \dp.rf.rf[30][21] ;
 wire \dp.rf.rf[30][22] ;
 wire \dp.rf.rf[30][23] ;
 wire \dp.rf.rf[30][24] ;
 wire \dp.rf.rf[30][25] ;
 wire \dp.rf.rf[30][26] ;
 wire \dp.rf.rf[30][27] ;
 wire \dp.rf.rf[30][28] ;
 wire \dp.rf.rf[30][29] ;
 wire \dp.rf.rf[30][2] ;
 wire \dp.rf.rf[30][30] ;
 wire \dp.rf.rf[30][31] ;
 wire \dp.rf.rf[30][3] ;
 wire \dp.rf.rf[30][4] ;
 wire \dp.rf.rf[30][5] ;
 wire \dp.rf.rf[30][6] ;
 wire \dp.rf.rf[30][7] ;
 wire \dp.rf.rf[30][8] ;
 wire \dp.rf.rf[30][9] ;
 wire \dp.rf.rf[31][0] ;
 wire \dp.rf.rf[31][10] ;
 wire \dp.rf.rf[31][11] ;
 wire \dp.rf.rf[31][12] ;
 wire \dp.rf.rf[31][13] ;
 wire \dp.rf.rf[31][14] ;
 wire \dp.rf.rf[31][15] ;
 wire \dp.rf.rf[31][16] ;
 wire \dp.rf.rf[31][17] ;
 wire \dp.rf.rf[31][18] ;
 wire \dp.rf.rf[31][19] ;
 wire \dp.rf.rf[31][1] ;
 wire \dp.rf.rf[31][20] ;
 wire \dp.rf.rf[31][21] ;
 wire \dp.rf.rf[31][22] ;
 wire \dp.rf.rf[31][23] ;
 wire \dp.rf.rf[31][24] ;
 wire \dp.rf.rf[31][25] ;
 wire \dp.rf.rf[31][26] ;
 wire \dp.rf.rf[31][27] ;
 wire \dp.rf.rf[31][28] ;
 wire \dp.rf.rf[31][29] ;
 wire \dp.rf.rf[31][2] ;
 wire \dp.rf.rf[31][30] ;
 wire \dp.rf.rf[31][31] ;
 wire \dp.rf.rf[31][3] ;
 wire \dp.rf.rf[31][4] ;
 wire \dp.rf.rf[31][5] ;
 wire \dp.rf.rf[31][6] ;
 wire \dp.rf.rf[31][7] ;
 wire \dp.rf.rf[31][8] ;
 wire \dp.rf.rf[31][9] ;
 wire \dp.rf.rf[3][0] ;
 wire \dp.rf.rf[3][10] ;
 wire \dp.rf.rf[3][11] ;
 wire \dp.rf.rf[3][12] ;
 wire \dp.rf.rf[3][13] ;
 wire \dp.rf.rf[3][14] ;
 wire \dp.rf.rf[3][15] ;
 wire \dp.rf.rf[3][16] ;
 wire \dp.rf.rf[3][17] ;
 wire \dp.rf.rf[3][18] ;
 wire \dp.rf.rf[3][19] ;
 wire \dp.rf.rf[3][1] ;
 wire \dp.rf.rf[3][20] ;
 wire \dp.rf.rf[3][21] ;
 wire \dp.rf.rf[3][22] ;
 wire \dp.rf.rf[3][23] ;
 wire \dp.rf.rf[3][24] ;
 wire \dp.rf.rf[3][25] ;
 wire \dp.rf.rf[3][26] ;
 wire \dp.rf.rf[3][27] ;
 wire \dp.rf.rf[3][28] ;
 wire \dp.rf.rf[3][29] ;
 wire \dp.rf.rf[3][2] ;
 wire \dp.rf.rf[3][30] ;
 wire \dp.rf.rf[3][31] ;
 wire \dp.rf.rf[3][3] ;
 wire \dp.rf.rf[3][4] ;
 wire \dp.rf.rf[3][5] ;
 wire \dp.rf.rf[3][6] ;
 wire \dp.rf.rf[3][7] ;
 wire \dp.rf.rf[3][8] ;
 wire \dp.rf.rf[3][9] ;
 wire \dp.rf.rf[4][0] ;
 wire \dp.rf.rf[4][10] ;
 wire \dp.rf.rf[4][11] ;
 wire \dp.rf.rf[4][12] ;
 wire \dp.rf.rf[4][13] ;
 wire \dp.rf.rf[4][14] ;
 wire \dp.rf.rf[4][15] ;
 wire \dp.rf.rf[4][16] ;
 wire \dp.rf.rf[4][17] ;
 wire \dp.rf.rf[4][18] ;
 wire \dp.rf.rf[4][19] ;
 wire \dp.rf.rf[4][1] ;
 wire \dp.rf.rf[4][20] ;
 wire \dp.rf.rf[4][21] ;
 wire \dp.rf.rf[4][22] ;
 wire \dp.rf.rf[4][23] ;
 wire \dp.rf.rf[4][24] ;
 wire \dp.rf.rf[4][25] ;
 wire \dp.rf.rf[4][26] ;
 wire \dp.rf.rf[4][27] ;
 wire \dp.rf.rf[4][28] ;
 wire \dp.rf.rf[4][29] ;
 wire \dp.rf.rf[4][2] ;
 wire \dp.rf.rf[4][30] ;
 wire \dp.rf.rf[4][31] ;
 wire \dp.rf.rf[4][3] ;
 wire \dp.rf.rf[4][4] ;
 wire \dp.rf.rf[4][5] ;
 wire \dp.rf.rf[4][6] ;
 wire \dp.rf.rf[4][7] ;
 wire \dp.rf.rf[4][8] ;
 wire \dp.rf.rf[4][9] ;
 wire \dp.rf.rf[5][0] ;
 wire \dp.rf.rf[5][10] ;
 wire \dp.rf.rf[5][11] ;
 wire \dp.rf.rf[5][12] ;
 wire \dp.rf.rf[5][13] ;
 wire \dp.rf.rf[5][14] ;
 wire \dp.rf.rf[5][15] ;
 wire \dp.rf.rf[5][16] ;
 wire \dp.rf.rf[5][17] ;
 wire \dp.rf.rf[5][18] ;
 wire \dp.rf.rf[5][19] ;
 wire \dp.rf.rf[5][1] ;
 wire \dp.rf.rf[5][20] ;
 wire \dp.rf.rf[5][21] ;
 wire \dp.rf.rf[5][22] ;
 wire \dp.rf.rf[5][23] ;
 wire \dp.rf.rf[5][24] ;
 wire \dp.rf.rf[5][25] ;
 wire \dp.rf.rf[5][26] ;
 wire \dp.rf.rf[5][27] ;
 wire \dp.rf.rf[5][28] ;
 wire \dp.rf.rf[5][29] ;
 wire \dp.rf.rf[5][2] ;
 wire \dp.rf.rf[5][30] ;
 wire \dp.rf.rf[5][31] ;
 wire \dp.rf.rf[5][3] ;
 wire \dp.rf.rf[5][4] ;
 wire \dp.rf.rf[5][5] ;
 wire \dp.rf.rf[5][6] ;
 wire \dp.rf.rf[5][7] ;
 wire \dp.rf.rf[5][8] ;
 wire \dp.rf.rf[5][9] ;
 wire \dp.rf.rf[6][0] ;
 wire \dp.rf.rf[6][10] ;
 wire \dp.rf.rf[6][11] ;
 wire \dp.rf.rf[6][12] ;
 wire \dp.rf.rf[6][13] ;
 wire \dp.rf.rf[6][14] ;
 wire \dp.rf.rf[6][15] ;
 wire \dp.rf.rf[6][16] ;
 wire \dp.rf.rf[6][17] ;
 wire \dp.rf.rf[6][18] ;
 wire \dp.rf.rf[6][19] ;
 wire \dp.rf.rf[6][1] ;
 wire \dp.rf.rf[6][20] ;
 wire \dp.rf.rf[6][21] ;
 wire \dp.rf.rf[6][22] ;
 wire \dp.rf.rf[6][23] ;
 wire \dp.rf.rf[6][24] ;
 wire \dp.rf.rf[6][25] ;
 wire \dp.rf.rf[6][26] ;
 wire \dp.rf.rf[6][27] ;
 wire \dp.rf.rf[6][28] ;
 wire \dp.rf.rf[6][29] ;
 wire \dp.rf.rf[6][2] ;
 wire \dp.rf.rf[6][30] ;
 wire \dp.rf.rf[6][31] ;
 wire \dp.rf.rf[6][3] ;
 wire \dp.rf.rf[6][4] ;
 wire \dp.rf.rf[6][5] ;
 wire \dp.rf.rf[6][6] ;
 wire \dp.rf.rf[6][7] ;
 wire \dp.rf.rf[6][8] ;
 wire \dp.rf.rf[6][9] ;
 wire \dp.rf.rf[7][0] ;
 wire \dp.rf.rf[7][10] ;
 wire \dp.rf.rf[7][11] ;
 wire \dp.rf.rf[7][12] ;
 wire \dp.rf.rf[7][13] ;
 wire \dp.rf.rf[7][14] ;
 wire \dp.rf.rf[7][15] ;
 wire \dp.rf.rf[7][16] ;
 wire \dp.rf.rf[7][17] ;
 wire \dp.rf.rf[7][18] ;
 wire \dp.rf.rf[7][19] ;
 wire \dp.rf.rf[7][1] ;
 wire \dp.rf.rf[7][20] ;
 wire \dp.rf.rf[7][21] ;
 wire \dp.rf.rf[7][22] ;
 wire \dp.rf.rf[7][23] ;
 wire \dp.rf.rf[7][24] ;
 wire \dp.rf.rf[7][25] ;
 wire \dp.rf.rf[7][26] ;
 wire \dp.rf.rf[7][27] ;
 wire \dp.rf.rf[7][28] ;
 wire \dp.rf.rf[7][29] ;
 wire \dp.rf.rf[7][2] ;
 wire \dp.rf.rf[7][30] ;
 wire \dp.rf.rf[7][31] ;
 wire \dp.rf.rf[7][3] ;
 wire \dp.rf.rf[7][4] ;
 wire \dp.rf.rf[7][5] ;
 wire \dp.rf.rf[7][6] ;
 wire \dp.rf.rf[7][7] ;
 wire \dp.rf.rf[7][8] ;
 wire \dp.rf.rf[7][9] ;
 wire \dp.rf.rf[8][0] ;
 wire \dp.rf.rf[8][10] ;
 wire \dp.rf.rf[8][11] ;
 wire \dp.rf.rf[8][12] ;
 wire \dp.rf.rf[8][13] ;
 wire \dp.rf.rf[8][14] ;
 wire \dp.rf.rf[8][15] ;
 wire \dp.rf.rf[8][16] ;
 wire \dp.rf.rf[8][17] ;
 wire \dp.rf.rf[8][18] ;
 wire \dp.rf.rf[8][19] ;
 wire \dp.rf.rf[8][1] ;
 wire \dp.rf.rf[8][20] ;
 wire \dp.rf.rf[8][21] ;
 wire \dp.rf.rf[8][22] ;
 wire \dp.rf.rf[8][23] ;
 wire \dp.rf.rf[8][24] ;
 wire \dp.rf.rf[8][25] ;
 wire \dp.rf.rf[8][26] ;
 wire \dp.rf.rf[8][27] ;
 wire \dp.rf.rf[8][28] ;
 wire \dp.rf.rf[8][29] ;
 wire \dp.rf.rf[8][2] ;
 wire \dp.rf.rf[8][30] ;
 wire \dp.rf.rf[8][31] ;
 wire \dp.rf.rf[8][3] ;
 wire \dp.rf.rf[8][4] ;
 wire \dp.rf.rf[8][5] ;
 wire \dp.rf.rf[8][6] ;
 wire \dp.rf.rf[8][7] ;
 wire \dp.rf.rf[8][8] ;
 wire \dp.rf.rf[8][9] ;
 wire \dp.rf.rf[9][0] ;
 wire \dp.rf.rf[9][10] ;
 wire \dp.rf.rf[9][11] ;
 wire \dp.rf.rf[9][12] ;
 wire \dp.rf.rf[9][13] ;
 wire \dp.rf.rf[9][14] ;
 wire \dp.rf.rf[9][15] ;
 wire \dp.rf.rf[9][16] ;
 wire \dp.rf.rf[9][17] ;
 wire \dp.rf.rf[9][18] ;
 wire \dp.rf.rf[9][19] ;
 wire \dp.rf.rf[9][1] ;
 wire \dp.rf.rf[9][20] ;
 wire \dp.rf.rf[9][21] ;
 wire \dp.rf.rf[9][22] ;
 wire \dp.rf.rf[9][23] ;
 wire \dp.rf.rf[9][24] ;
 wire \dp.rf.rf[9][25] ;
 wire \dp.rf.rf[9][26] ;
 wire \dp.rf.rf[9][27] ;
 wire \dp.rf.rf[9][28] ;
 wire \dp.rf.rf[9][29] ;
 wire \dp.rf.rf[9][2] ;
 wire \dp.rf.rf[9][30] ;
 wire \dp.rf.rf[9][31] ;
 wire \dp.rf.rf[9][3] ;
 wire \dp.rf.rf[9][4] ;
 wire \dp.rf.rf[9][5] ;
 wire \dp.rf.rf[9][6] ;
 wire \dp.rf.rf[9][7] ;
 wire \dp.rf.rf[9][8] ;
 wire \dp.rf.rf[9][9] ;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire [0:0] _05093_;
 wire [0:0] _05095_;
 wire [0:0] _05096_;
 wire [0:0] _05097_;
 wire [0:0] _05098_;
 wire [0:0] _05099_;
 wire [0:0] _05100_;
 wire [0:0] _05101_;
 wire [0:0] _05102_;
 wire [0:0] _05104_;
 wire [0:0] _05105_;
 wire [0:0] _05106_;
 wire [0:0] _05107_;
 wire [0:0] _05108_;
 wire [0:0] _05109_;
 wire [0:0] _05110_;
 wire [0:0] _05111_;
 wire [0:0] _05113_;
 wire [0:0] _05114_;
 wire [0:0] _05115_;
 wire [0:0] _05117_;
 wire [0:0] _05118_;
 wire [0:0] _05120_;
 wire [0:0] _05121_;
 wire [0:0] _05122_;
 wire [0:0] _05123_;
 wire [0:0] _05124_;
 wire [0:0] _05125_;
 wire [0:0] _05126_;
 wire [0:0] _05127_;
 wire [0:0] _05128_;
 wire [0:0] _05129_;
 wire [0:0] _05130_;
 wire [0:0] _05131_;
 wire [0:0] _05132_;
 wire [0:0] _05133_;
 wire [0:0] _05134_;
 wire [0:0] _05135_;
 wire [0:0] _05136_;
 wire [0:0] _05137_;
 wire [0:0] _05138_;
 wire [0:0] _05139_;
 wire [0:0] _05140_;
 wire [0:0] _05141_;
 wire [0:0] _05142_;
 wire [0:0] _05144_;
 wire [0:0] _05145_;
 wire [0:0] _05146_;
 wire [0:0] _05147_;
 wire [0:0] _05148_;
 wire [0:0] _05149_;
 wire [0:0] _05150_;
 wire [0:0] _05152_;
 wire [0:0] _05153_;
 wire [0:0] _05154_;
 wire [0:0] _05155_;
 wire [0:0] _05156_;
 wire [0:0] _05157_;
 wire [0:0] _05158_;
 wire [0:0] _05159_;
 wire [0:0] _05160_;
 wire [0:0] _05161_;
 wire [0:0] _05162_;
 wire [0:0] _05163_;
 wire [0:0] _05164_;
 wire [0:0] _05165_;
 wire [0:0] _05166_;
 wire [0:0] _05168_;
 wire [0:0] _05169_;
 wire [0:0] _05170_;
 wire [0:0] _05171_;
 wire [0:0] _05172_;
 wire [0:0] _05173_;
 wire [0:0] _05174_;
 wire [0:0] _05176_;
 wire [0:0] _05177_;
 wire [0:0] _05178_;
 wire [0:0] _05179_;
 wire [0:0] _05180_;
 wire [0:0] _05181_;
 wire [0:0] _05182_;
 wire [0:0] _05184_;
 wire [0:0] _05185_;
 wire [0:0] _05186_;
 wire [0:0] _05187_;
 wire [0:0] _05188_;
 wire [0:0] _05189_;
 wire [0:0] _05190_;
 wire [0:0] _05192_;
 wire [0:0] _05193_;
 wire [0:0] _05194_;
 wire [0:0] _05195_;
 wire [0:0] _05196_;
 wire [0:0] _05197_;
 wire [0:0] _05198_;
 wire [0:0] _05200_;
 wire [0:0] _05201_;
 wire [0:0] _05202_;
 wire [0:0] _05203_;
 wire [0:0] _05204_;
 wire [0:0] _05205_;
 wire [0:0] _05206_;
 wire [0:0] _05208_;
 wire [0:0] _05209_;
 wire [0:0] _05210_;
 wire [0:0] _05211_;
 wire [0:0] _05212_;
 wire [0:0] _05213_;
 wire [0:0] _05214_;
 wire [0:0] _05216_;
 wire [0:0] _05217_;
 wire [0:0] _05218_;
 wire [0:0] _05219_;
 wire [0:0] _05220_;
 wire [0:0] _05221_;
 wire [0:0] _05222_;
 wire [0:0] _05224_;
 wire [0:0] _05225_;
 wire [0:0] _05226_;
 wire [0:0] _05227_;
 wire [0:0] _05228_;
 wire [0:0] _05229_;
 wire [0:0] _05230_;
 wire [0:0] _05232_;
 wire [0:0] _05233_;
 wire [0:0] _05234_;
 wire [0:0] _05235_;
 wire [0:0] _05236_;
 wire [0:0] _05237_;
 wire [0:0] _05238_;
 wire [0:0] _05240_;
 wire [0:0] _05241_;
 wire [0:0] _05242_;
 wire [0:0] _05243_;
 wire [0:0] _05244_;
 wire [0:0] _05245_;
 wire [0:0] _05246_;
 wire [0:0] _05248_;
 wire [0:0] _05249_;
 wire [0:0] _05250_;
 wire [0:0] _05251_;
 wire [0:0] _05252_;
 wire [0:0] _05253_;
 wire [0:0] _05254_;
 wire [0:0] _05256_;
 wire [0:0] _05257_;
 wire [0:0] _05258_;
 wire [0:0] _05259_;
 wire [0:0] _05260_;
 wire [0:0] _05261_;
 wire [0:0] _05262_;
 wire [0:0] _05264_;
 wire [0:0] _05265_;
 wire [0:0] _05266_;
 wire [0:0] _05267_;
 wire [0:0] _05268_;
 wire [0:0] _05269_;
 wire [0:0] _05270_;
 wire [0:0] _05272_;
 wire [0:0] _05273_;
 wire [0:0] _05274_;
 wire [0:0] _05275_;
 wire [0:0] _05276_;
 wire [0:0] _05277_;
 wire [0:0] _05278_;
 wire [0:0] _05280_;
 wire [0:0] _05281_;
 wire [0:0] _05282_;
 wire [0:0] _05283_;
 wire [0:0] _05284_;
 wire [0:0] _05285_;
 wire [0:0] _05286_;
 wire [0:0] _05288_;
 wire [0:0] _05289_;
 wire [0:0] _05290_;
 wire [0:0] _05291_;
 wire [0:0] _05292_;
 wire [0:0] _05293_;
 wire [0:0] _05294_;
 wire [0:0] _05296_;
 wire [0:0] _05297_;
 wire [0:0] _05298_;
 wire [0:0] _05299_;
 wire [0:0] _05300_;
 wire [0:0] _05301_;
 wire [0:0] _05302_;
 wire [0:0] _05303_;
 wire [0:0] _05304_;
 wire [0:0] _05305_;
 wire [0:0] _05306_;
 wire [0:0] _05307_;
 wire [0:0] _05308_;
 wire [0:0] _05309_;
 wire [0:0] _05310_;
 wire [0:0] _05312_;
 wire [0:0] _05313_;
 wire [0:0] _05314_;
 wire [0:0] _05315_;
 wire [0:0] _05316_;
 wire [0:0] _05317_;
 wire [0:0] _05318_;
 wire [0:0] _05320_;
 wire [0:0] _05321_;
 wire [0:0] _05322_;
 wire [0:0] _05323_;
 wire [0:0] _05324_;
 wire [0:0] _05325_;
 wire [0:0] _05326_;
 wire [0:0] _05328_;
 wire [0:0] _05329_;
 wire [0:0] _05330_;
 wire [0:0] _05331_;
 wire [0:0] _05332_;
 wire [0:0] _05333_;
 wire [0:0] _05334_;
 wire [0:0] _05336_;
 wire [0:0] _05337_;
 wire [0:0] _05338_;
 wire [0:0] _05339_;
 wire [0:0] _05340_;
 wire [0:0] _05341_;
 wire [0:0] _05342_;
 wire [0:0] _05344_;
 wire [0:0] _05345_;
 wire [0:0] _05346_;
 wire [0:0] _05347_;
 wire [0:0] _05348_;
 wire [0:0] _05349_;
 wire [0:0] _05350_;
 wire [0:0] _05351_;
 wire [0:0] _05352_;
 wire [0:0] _05353_;
 wire [0:0] _05354_;
 wire [0:0] _05355_;
 wire [0:0] _05356_;
 wire [0:0] _05357_;
 wire [0:0] _05358_;
 wire [0:0] _05359_;
 wire [0:0] _05360_;
 wire [0:0] _05361_;
 wire [0:0] _05362_;
 wire [0:0] _05363_;
 wire [0:0] _05364_;
 wire [0:0] _05365_;
 wire [0:0] _05366_;
 wire [0:0] _05367_;
 wire [0:0] _05368_;
 wire [0:0] _05369_;
 wire [0:0] _05370_;
 wire [0:0] _05371_;
 wire [0:0] _05372_;
 wire [0:0] _05373_;
 wire [0:0] _05374_;
 wire [0:0] _05375_;
 wire [0:0] _05376_;
 wire [0:0] _05377_;
 wire [0:0] _05378_;
 wire [0:0] _05379_;
 wire [0:0] _05380_;
 wire [0:0] _05381_;
 wire [0:0] _05382_;
 wire [0:0] _05383_;
 wire [0:0] _05384_;
 wire [0:0] _05385_;
 wire [0:0] _05386_;
 wire [0:0] _05387_;
 wire [0:0] _05388_;
 wire [0:0] _05389_;
 wire [0:0] _05390_;
 wire [0:0] _05391_;
 wire [0:0] _05392_;
 wire [0:0] _05393_;
 wire [0:0] _05394_;
 wire [0:0] _05395_;
 wire [0:0] _05396_;
 wire [0:0] _05397_;
 wire [0:0] _05398_;
 wire [0:0] _05399_;
 wire [0:0] _05400_;
 wire [0:0] _05401_;
 wire [0:0] _05402_;
 wire [0:0] _05403_;
 wire [0:0] _05404_;
 wire [0:0] _05405_;
 wire [0:0] _05406_;
 wire [0:0] _05407_;
 wire [0:0] _05408_;
 wire [0:0] _05409_;
 wire [0:0] _05410_;
 wire [0:0] _05411_;
 wire [0:0] _05412_;
 wire [0:0] _05413_;
 wire [0:0] _05414_;
 wire [0:0] _05415_;
 wire [0:0] _05416_;
 wire [0:0] _05417_;
 wire [0:0] _05418_;
 wire [0:0] _05419_;
 wire [0:0] _05420_;
 wire [0:0] _05421_;
 wire [0:0] _05422_;
 wire [0:0] _05423_;
 wire [0:0] _05424_;
 wire [0:0] _05425_;
 wire [0:0] _05426_;
 wire [0:0] _05427_;
 wire [0:0] _05428_;
 wire [0:0] _05429_;
 wire [0:0] _05430_;
 wire [0:0] _05431_;
 wire [0:0] _05432_;
 wire [0:0] _05433_;
 wire [0:0] _05434_;
 wire [0:0] _05435_;
 wire [0:0] _05436_;
 wire [0:0] _05437_;
 wire [0:0] _05438_;
 wire [0:0] _05439_;
 wire [0:0] _05440_;
 wire [0:0] _05441_;
 wire [0:0] _05442_;
 wire [0:0] _05443_;
 wire [0:0] _05444_;
 wire [0:0] _05445_;
 wire [0:0] _05446_;
 wire [0:0] _05447_;
 wire [0:0] _05448_;
 wire [0:0] _05449_;
 wire [0:0] _05450_;
 wire [0:0] _05451_;
 wire [0:0] _05452_;
 wire [0:0] _05453_;
 wire [0:0] _05454_;
 wire [0:0] _05455_;
 wire [0:0] _05456_;
 wire [0:0] _05457_;
 wire [0:0] _05458_;
 wire [0:0] _05459_;
 wire [0:0] _05460_;
 wire [0:0] _05461_;
 wire [0:0] _05462_;
 wire [0:0] _05463_;
 wire [0:0] _05464_;
 wire [0:0] _05465_;
 wire [0:0] _05466_;
 wire [0:0] _05467_;
 wire [0:0] _05468_;
 wire [0:0] _05469_;
 wire [0:0] _05470_;
 wire [0:0] _05471_;
 wire [0:0] _05472_;
 wire [0:0] _05473_;
 wire [0:0] _05474_;
 wire [0:0] _05475_;
 wire [0:0] _05476_;
 wire [0:0] _05477_;
 wire [0:0] _05478_;
 wire [0:0] _05479_;

 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_48__f_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_6_48__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_47__f_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_6_47__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _05482_ (.I(net28),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05483_ (.A1(net1),
    .A2(net12),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_46__f_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_6_46__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05485_ (.A1(net26),
    .A2(net23),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _05486_ (.A1(net27),
    .A2(_01029_),
    .A3(net533),
    .A4(_01032_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05487_ (.A1(net29),
    .A2(_01033_),
    .ZN(net99));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_45__f_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_6_45__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_44__f_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_6_44__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _05490_ (.I(net14),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_43__f_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_6_43__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_42__f_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_6_42__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05493_ (.I0(\dp.rf.rf[17][0] ),
    .I1(\dp.rf.rf[21][0] ),
    .S(net15),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05494_ (.I0(\dp.rf.rf[16][0] ),
    .I1(\dp.rf.rf[20][0] ),
    .S(net15),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05495_ (.I0(\dp.rf.rf[25][0] ),
    .I1(\dp.rf.rf[29][0] ),
    .S(net15),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05496_ (.I0(\dp.rf.rf[24][0] ),
    .I1(\dp.rf.rf[28][0] ),
    .S(net15),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_41__f_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_6_41__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_40__f_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_6_40__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _05499_ (.I(net547),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_39__f_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_6_39__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05501_ (.I0(_01039_),
    .I1(_01040_),
    .I2(_01041_),
    .I3(_01042_),
    .S0(_01045_),
    .S1(net16),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _05502_ (.A1(net17),
    .A2(_01036_),
    .A3(_01047_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_38__f_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_6_38__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_37__f_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_6_37__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_36__f_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_6_36__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05506_ (.I0(\dp.rf.rf[0][0] ),
    .I1(\dp.rf.rf[1][0] ),
    .I2(\dp.rf.rf[2][0] ),
    .I3(\dp.rf.rf[3][0] ),
    .S0(net13),
    .S1(net546),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05507_ (.A1(net15),
    .A2(_01052_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_35__f_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_6_35__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _05509_ (.I(net15),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05510_ (.I0(\dp.rf.rf[4][0] ),
    .I1(\dp.rf.rf[5][0] ),
    .S(net13),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _05511_ (.A1(net14),
    .A2(net13),
    .A3(net15),
    .A4(net16),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _05512_ (.A1(net546),
    .A2(_01055_),
    .A3(_01056_),
    .B1(_01057_),
    .B2(net17),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_34__f_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_6_34__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05514_ (.A1(net546),
    .A2(net15),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_33__f_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_6_33__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05516_ (.I0(\dp.rf.rf[6][0] ),
    .I1(\dp.rf.rf[7][0] ),
    .S(net13),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05517_ (.A1(_01060_),
    .A2(_01062_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _05518_ (.I(net17),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_32__f_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_6_32__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _05520_ (.I(net16),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05521_ (.A1(_01064_),
    .A2(_01066_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _05522_ (.A1(_01053_),
    .A2(_01058_),
    .A3(_01063_),
    .A4(_01067_),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_31__f_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_6_31__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_30__f_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_6_30__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_29__f_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_6_29__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_28__f_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_6_28__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05527_ (.I0(\dp.rf.rf[26][0] ),
    .I1(\dp.rf.rf[27][0] ),
    .I2(\dp.rf.rf[30][0] ),
    .I3(\dp.rf.rf[31][0] ),
    .S0(net13),
    .S1(net15),
    .Z(_01073_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05528_ (.I0(\dp.rf.rf[18][0] ),
    .I1(\dp.rf.rf[19][0] ),
    .I2(\dp.rf.rf[22][0] ),
    .I3(\dp.rf.rf[23][0] ),
    .S0(net13),
    .S1(net15),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_27__f_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_6_27__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05530_ (.I0(_01073_),
    .I1(_01074_),
    .S(_01066_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _05531_ (.A1(net17),
    .A2(net546),
    .A3(_01076_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05532_ (.I0(\dp.rf.rf[10][0] ),
    .I1(\dp.rf.rf[11][0] ),
    .S(net13),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _05533_ (.A1(_01036_),
    .A2(net15),
    .A3(_01078_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_26__f_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_6_26__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05535_ (.I0(\dp.rf.rf[8][0] ),
    .I1(\dp.rf.rf[9][0] ),
    .I2(\dp.rf.rf[12][0] ),
    .I3(\dp.rf.rf[13][0] ),
    .S0(net13),
    .S1(net15),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05536_ (.A1(net546),
    .A2(_01081_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_25__f_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_6_25__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05538_ (.A1(_01064_),
    .A2(net16),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05539_ (.I0(\dp.rf.rf[14][0] ),
    .I1(\dp.rf.rf[15][0] ),
    .S(net13),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05540_ (.A1(_01060_),
    .A2(_01085_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _05541_ (.A1(_01079_),
    .A2(_01082_),
    .A3(_01084_),
    .A4(_01086_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _05542_ (.A1(_01048_),
    .A2(_01068_),
    .A3(_01077_),
    .A4(_01087_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05543_ (.I(_01088_),
    .ZN(net133));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05544_ (.I(net5),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_24__f_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_6_24__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_23__f_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_6_23__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _05547_ (.A1(net29),
    .A2(net533),
    .A3(_01032_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_22__f_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_6_22__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05549_ (.A1(net28),
    .A2(net24),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05550_ (.I(net4),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _05551_ (.A1(net28),
    .A2(_01095_),
    .A3(_01089_),
    .A4(net24),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05552_ (.A1(net5),
    .A2(_01094_),
    .B1(_01092_),
    .B2(_01096_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05553_ (.I(net27),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05554_ (.A1(_01089_),
    .A2(_01092_),
    .B1(_01097_),
    .B2(_01098_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05555_ (.I(net6),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05556_ (.A1(net23),
    .A2(net27),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_21__f_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_6_21__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05558_ (.A1(net29),
    .A2(_01101_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05559_ (.A1(net28),
    .A2(net29),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _05560_ (.A1(net23),
    .A2(net27),
    .A3(_01104_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05561_ (.I(net26),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05562_ (.A1(net1),
    .A2(net12),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _05563_ (.A1(_01103_),
    .A2(_01105_),
    .B(_01106_),
    .C(_01107_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05564_ (.A1(_01100_),
    .A2(_01108_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05565_ (.A1(_01099_),
    .A2(_01109_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_20__f_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_6_20__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05567_ (.A1(net26),
    .A2(net23),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05568_ (.I0(net29),
    .I1(net27),
    .S(net28),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05569_ (.I(_01113_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05570_ (.A1(net28),
    .A2(net29),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05571_ (.A1(net26),
    .A2(net29),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05572_ (.I0(_01115_),
    .I1(_01116_),
    .S(net27),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05573_ (.A1(_01112_),
    .A2(_01114_),
    .B1(_01117_),
    .B2(net23),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05574_ (.A1(net533),
    .A2(_01118_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_19__f_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_6_19__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_18__f_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_6_18__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05577_ (.A1(net26),
    .A2(net23),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _05578_ (.A1(_01098_),
    .A2(_01107_),
    .A3(_01115_),
    .A4(_01122_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_17__f_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_6_17__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05580_ (.A1(net26),
    .A2(net29),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _05581_ (.A1(_01125_),
    .A2(_01101_),
    .A3(_01030_),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_16__f_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_6_16__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _05583_ (.A1(net13),
    .A2(_01033_),
    .A3(_01123_),
    .A4(net528),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05584_ (.A1(net29),
    .A2(net31),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05585_ (.A1(_01036_),
    .A2(_01123_),
    .B1(_01129_),
    .B2(_01033_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05586_ (.I(net30),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _05587_ (.A1(net29),
    .A2(_01131_),
    .A3(_01033_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _05588_ (.A1(_01128_),
    .A2(_01130_),
    .A3(_01132_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _05589_ (.A1(net26),
    .A2(net23),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _05590_ (.A1(_01098_),
    .A2(_01107_),
    .A3(_01115_),
    .A4(_01134_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _05591_ (.A1(net533),
    .A2(_01118_),
    .A3(_01135_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _05592_ (.A1(_01088_),
    .A2(_01119_),
    .B1(_01133_),
    .B2(_01136_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_15__f_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_6_15__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_14__f_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_6_14__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _05595_ (.A1(_01110_),
    .A2(net509),
    .ZN(_05104_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05596_ (.I(_05104_[0]),
    .ZN(_05108_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _05597_ (.I(net8),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_13__f_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_6_13__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_12__f_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_6_12__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_11__f_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_6_11__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _05601_ (.I(net10),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_10__f_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_6_10__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_9__f_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_6_9__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05604_ (.A1(_01140_),
    .A2(_01144_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _05605_ (.I(net7),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_8__f_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_6_8__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_7__f_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_6_7__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_6__f_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_6_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_5__f_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_6_5__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_4__f_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_6_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05611_ (.A1(\dp.rf.rf[4][0] ),
    .A2(net531),
    .A3(net9),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_3__f_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_6_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_2__f_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_6_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_1__f_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_6_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_0__f_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_6_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05617_ (.I0(\dp.rf.rf[1][0] ),
    .I1(\dp.rf.rf[5][0] ),
    .S(net9),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05618_ (.A1(net7),
    .A2(_01160_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05621_ (.A1(_01147_),
    .A2(_01154_),
    .A3(_01161_),
    .B(net526),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _05622_ (.A1(net23),
    .A2(net27),
    .A3(_01107_),
    .A4(_01116_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _05624_ (.I(net9),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05625_ (.A1(net531),
    .A2(_01167_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05626_ (.A1(_01165_),
    .A2(_01168_),
    .B(\dp.rf.rf[0][0] ),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05627_ (.A1(_01164_),
    .A2(_01169_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05633_ (.I0(\dp.rf.rf[2][0] ),
    .I1(\dp.rf.rf[3][0] ),
    .I2(\dp.rf.rf[6][0] ),
    .I3(\dp.rf.rf[7][0] ),
    .S0(net542),
    .S1(net9),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05634_ (.A1(net533),
    .A2(net532),
    .A3(_01125_),
    .B(_01144_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05635_ (.A1(_01176_),
    .A2(_01177_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05636_ (.A1(net8),
    .A2(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05637_ (.A1(net533),
    .A2(net532),
    .A3(_01125_),
    .B(net8),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05641_ (.I0(\dp.rf.rf[14][0] ),
    .I1(\dp.rf.rf[15][0] ),
    .S(net542),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05642_ (.A1(_01167_),
    .A2(_01184_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _05643_ (.A1(net11),
    .A2(net523),
    .A3(_01185_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05644_ (.A1(net533),
    .A2(net532),
    .A3(_01125_),
    .B(net9),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05646_ (.I(\dp.rf.rf[10][0] ),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _05648_ (.A1(_01189_),
    .A2(_01030_),
    .A3(_01101_),
    .A4(_01125_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05651_ (.I0(\dp.rf.rf[10][0] ),
    .I1(\dp.rf.rf[11][0] ),
    .S(net542),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05652_ (.I(_01194_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _05653_ (.A1(net522),
    .A2(_01191_),
    .A3(_01195_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _05654_ (.A1(net7),
    .A2(net8),
    .A3(net9),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05655_ (.A1(_01144_),
    .A2(_01197_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_712_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_712_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_711_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_711_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_705_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_705_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_704_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_704_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_702_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_702_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05662_ (.I0(\dp.rf.rf[9][0] ),
    .I1(\dp.rf.rf[13][0] ),
    .S(net9),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _05663_ (.A1(net542),
    .A2(_01140_),
    .A3(net10),
    .A4(_01205_),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_700_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_700_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05665_ (.A1(net7),
    .A2(net8),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05666_ (.I0(\dp.rf.rf[8][0] ),
    .I1(\dp.rf.rf[12][0] ),
    .S(net9),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05667_ (.A1(net10),
    .A2(_01208_),
    .A3(_01209_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _05668_ (.A1(_01198_),
    .A2(_01206_),
    .A3(_01210_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _05669_ (.I(net11),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_698_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_698_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05671_ (.A1(_01212_),
    .A2(net526),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05672_ (.A1(_01186_),
    .A2(_01196_),
    .B1(_01211_),
    .B2(_01214_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05673_ (.A1(net11),
    .A2(net166),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_697_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_697_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_694_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_694_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05676_ (.I0(\dp.rf.rf[24][0] ),
    .I1(\dp.rf.rf[25][0] ),
    .I2(\dp.rf.rf[26][0] ),
    .I3(\dp.rf.rf[27][0] ),
    .S0(net542),
    .S1(net8),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05677_ (.I0(\dp.rf.rf[16][0] ),
    .I1(\dp.rf.rf[17][0] ),
    .I2(\dp.rf.rf[18][0] ),
    .I3(\dp.rf.rf[19][0] ),
    .S0(net542),
    .S1(net8),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05678_ (.I0(_01219_),
    .I1(_01220_),
    .S(_01144_),
    .Z(_01221_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05679_ (.I0(\dp.rf.rf[21][0] ),
    .I1(\dp.rf.rf[23][0] ),
    .I2(\dp.rf.rf[29][0] ),
    .I3(\dp.rf.rf[31][0] ),
    .S0(net8),
    .S1(net10),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05680_ (.I0(\dp.rf.rf[20][0] ),
    .I1(\dp.rf.rf[22][0] ),
    .I2(\dp.rf.rf[28][0] ),
    .I3(\dp.rf.rf[30][0] ),
    .S0(net8),
    .S1(net10),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05681_ (.I0(_01222_),
    .I1(_01223_),
    .S(net531),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_693_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_693_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_692_clk (.I(clknet_6_3__leaf_clk),
    .Z(clknet_leaf_692_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_689_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_689_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05685_ (.I0(_01221_),
    .I1(_01224_),
    .S(net9),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05686_ (.A1(_01216_),
    .A2(_01228_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05687_ (.A1(_01170_),
    .A2(_01179_),
    .A3(_01215_),
    .B(_01229_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_688_clk (.I(clknet_6_3__leaf_clk),
    .Z(clknet_leaf_688_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _05689_ (.I(_01230_),
    .ZN(_05107_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05690_ (.A1(net10),
    .A2(net11),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05691_ (.A1(net8),
    .A2(_01231_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _05692_ (.A1(_01165_),
    .A2(_01168_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05693_ (.I(\dp.rf.rf[3][31] ),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_687_clk (.I(clknet_6_3__leaf_clk),
    .Z(clknet_leaf_687_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05695_ (.I(\dp.rf.rf[7][31] ),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05696_ (.A1(_01234_),
    .A2(net537),
    .B1(net521),
    .B2(_01236_),
    .C(net540),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05697_ (.I(\dp.rf.rf[6][31] ),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05698_ (.A1(_01238_),
    .A2(net521),
    .B(_01148_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05699_ (.A1(\dp.rf.rf[2][31] ),
    .A2(_01233_),
    .B1(_01237_),
    .B2(_01239_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _05700_ (.A1(_01165_),
    .A2(_01232_),
    .A3(_01240_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _05701_ (.A1(_01212_),
    .A2(net168),
    .A3(_01198_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05702_ (.A1(_01140_),
    .A2(net165),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05703_ (.I(\dp.rf.rf[4][31] ),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05704_ (.A1(_01148_),
    .A2(net9),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05705_ (.I(\dp.rf.rf[1][31] ),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05706_ (.I(\dp.rf.rf[5][31] ),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05707_ (.I0(_01246_),
    .I1(_01247_),
    .S(net537),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05708_ (.A1(_01244_),
    .A2(net520),
    .B1(_01248_),
    .B2(_01148_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05709_ (.A1(net165),
    .A2(_01197_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05710_ (.A1(_01243_),
    .A2(_01249_),
    .B1(_01250_),
    .B2(\dp.rf.rf[0][31] ),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_685_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_685_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05712_ (.I0(\dp.rf.rf[17][31] ),
    .I1(\dp.rf.rf[19][31] ),
    .S(net8),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05713_ (.A1(net531),
    .A2(_01253_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05714_ (.I(\dp.rf.rf[18][31] ),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _05715_ (.A1(_01255_),
    .A2(net531),
    .A3(net8),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05716_ (.A1(net9),
    .A2(_01254_),
    .A3(_01256_),
    .B(net526),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05717_ (.I(\dp.rf.rf[16][31] ),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05718_ (.A1(_01258_),
    .A2(net530),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05719_ (.I(\dp.rf.rf[20][31] ),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05720_ (.I(\dp.rf.rf[21][31] ),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05721_ (.I(\dp.rf.rf[22][31] ),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05722_ (.I(\dp.rf.rf[23][31] ),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05723_ (.I0(_01260_),
    .I1(_01261_),
    .I2(_01262_),
    .I3(_01263_),
    .S0(net7),
    .S1(net8),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05724_ (.A1(net522),
    .A2(_01264_),
    .B(_01144_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05725_ (.A1(_01257_),
    .A2(_01259_),
    .B(_01265_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05726_ (.I(\dp.rf.rf[25][31] ),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _05727_ (.A1(_01267_),
    .A2(net540),
    .A3(_01140_),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05728_ (.A1(net540),
    .A2(net8),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05729_ (.I0(\dp.rf.rf[24][31] ),
    .I1(\dp.rf.rf[26][31] ),
    .S(net8),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05730_ (.A1(\dp.rf.rf[27][31] ),
    .A2(_01269_),
    .B1(_01270_),
    .B2(net540),
    .C(_01167_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05731_ (.A1(net165),
    .A2(_01268_),
    .B(_01271_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05732_ (.A1(_01030_),
    .A2(_01101_),
    .A3(_01125_),
    .B(net10),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_684_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_684_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05734_ (.I0(\dp.rf.rf[28][31] ),
    .I1(\dp.rf.rf[29][31] ),
    .I2(\dp.rf.rf[30][31] ),
    .I3(\dp.rf.rf[31][31] ),
    .S0(net540),
    .S1(net8),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05735_ (.A1(net9),
    .A2(_01275_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05736_ (.A1(_01272_),
    .A2(net519),
    .A3(_01276_),
    .B(_01216_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05737_ (.A1(net10),
    .A2(_01212_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _05738_ (.A1(_01140_),
    .A2(net167),
    .A3(_01278_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_682_clk (.I(clknet_6_3__leaf_clk),
    .Z(clknet_leaf_682_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _05740_ (.I0(\dp.rf.rf[8][31] ),
    .I1(\dp.rf.rf[9][31] ),
    .I2(\dp.rf.rf[12][31] ),
    .I3(\dp.rf.rf[13][31] ),
    .S0(net541),
    .S1(net9),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05741_ (.I0(\dp.rf.rf[10][31] ),
    .I1(\dp.rf.rf[11][31] ),
    .I2(\dp.rf.rf[14][31] ),
    .I3(\dp.rf.rf[15][31] ),
    .S0(net541),
    .S1(net9),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05742_ (.A1(_01278_),
    .A2(_01282_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05743_ (.A1(net8),
    .A2(net166),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05744_ (.A1(_01279_),
    .A2(_01281_),
    .B1(_01283_),
    .B2(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _05745_ (.A1(net516),
    .A2(_01251_),
    .B1(_01266_),
    .B2(_01277_),
    .C(_01285_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05746_ (.A1(_01241_),
    .A2(_01286_),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _05747_ (.I(_01287_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_681_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_681_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_680_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_680_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05750_ (.I(net25),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_679_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_679_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_678_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_678_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05753_ (.I0(\dp.rf.rf[24][31] ),
    .I1(\dp.rf.rf[25][31] ),
    .I2(\dp.rf.rf[26][31] ),
    .I3(\dp.rf.rf[27][31] ),
    .S0(net13),
    .S1(net14),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05754_ (.I0(\dp.rf.rf[16][31] ),
    .I1(\dp.rf.rf[17][31] ),
    .I2(\dp.rf.rf[18][31] ),
    .I3(\dp.rf.rf[19][31] ),
    .S0(net13),
    .S1(net546),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_675_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_675_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05756_ (.I0(\dp.rf.rf[28][31] ),
    .I1(\dp.rf.rf[29][31] ),
    .I2(\dp.rf.rf[30][31] ),
    .I3(\dp.rf.rf[31][31] ),
    .S0(net13),
    .S1(net14),
    .Z(_01296_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05757_ (.I0(\dp.rf.rf[20][31] ),
    .I1(\dp.rf.rf[21][31] ),
    .I2(\dp.rf.rf[22][31] ),
    .I3(\dp.rf.rf[23][31] ),
    .S0(net13),
    .S1(net546),
    .Z(_01297_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_673_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_673_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_670_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_670_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _05760_ (.I0(_01293_),
    .I1(_01294_),
    .I2(_01296_),
    .I3(_01297_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_668_clk (.I(clknet_6_3__leaf_clk),
    .Z(clknet_leaf_668_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05762_ (.I0(\dp.rf.rf[8][31] ),
    .I1(\dp.rf.rf[9][31] ),
    .I2(\dp.rf.rf[10][31] ),
    .I3(\dp.rf.rf[11][31] ),
    .S0(net549),
    .S1(net14),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05763_ (.I0(\dp.rf.rf[0][31] ),
    .I1(\dp.rf.rf[1][31] ),
    .I2(\dp.rf.rf[2][31] ),
    .I3(\dp.rf.rf[3][31] ),
    .S0(net549),
    .S1(net14),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05764_ (.I0(\dp.rf.rf[12][31] ),
    .I1(\dp.rf.rf[13][31] ),
    .I2(\dp.rf.rf[14][31] ),
    .I3(\dp.rf.rf[15][31] ),
    .S0(net549),
    .S1(net14),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05765_ (.I0(\dp.rf.rf[4][31] ),
    .I1(\dp.rf.rf[5][31] ),
    .I2(\dp.rf.rf[6][31] ),
    .I3(\dp.rf.rf[7][31] ),
    .S0(net549),
    .S1(net14),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_665_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_665_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_664_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_664_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _05768_ (.I0(_01302_),
    .I1(_01303_),
    .I2(_01304_),
    .I3(_01305_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05769_ (.A1(_01064_),
    .A2(_01057_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _05770_ (.A1(net17),
    .A2(_01300_),
    .B1(_01308_),
    .B2(_01309_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05771_ (.A1(net533),
    .A2(_01118_),
    .Z(_01311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05772_ (.I0(_01290_),
    .I1(_01310_),
    .S(_01311_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05773_ (.A1(net511),
    .A2(_01312_),
    .Z(_05111_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05774_ (.I(_05111_[0]),
    .ZN(_05115_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_662_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_662_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_658_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_658_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05777_ (.A1(_01123_),
    .A2(net527),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05778_ (.A1(_01033_),
    .A2(_01315_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _05779_ (.A1(_01098_),
    .A2(net28),
    .A3(_01107_),
    .A4(_01112_),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _05780_ (.A1(_01098_),
    .A2(_01107_),
    .A3(_01115_),
    .A4(_01122_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05781_ (.A1(_01317_),
    .A2(_01318_),
    .B(net25),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05782_ (.A1(_01316_),
    .A2(_01319_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_657_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_657_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_656_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_656_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05785_ (.A1(net24),
    .A2(_01165_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _05786_ (.A1(_01033_),
    .A2(_01123_),
    .A3(net527),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05787_ (.A1(_01290_),
    .A2(_01324_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_655_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_655_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05789_ (.A1(_01320_),
    .A2(_01323_),
    .B(_01325_),
    .ZN(_05477_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_654_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_654_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_652_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_652_clk));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05792_ (.A1(net17),
    .A2(_01057_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_651_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_651_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_649_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_649_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_647_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_647_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05796_ (.I0(\dp.rf.rf[24][30] ),
    .I1(\dp.rf.rf[25][30] ),
    .I2(\dp.rf.rf[26][30] ),
    .I3(\dp.rf.rf[27][30] ),
    .S0(net13),
    .S1(net14),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05797_ (.I0(\dp.rf.rf[16][30] ),
    .I1(\dp.rf.rf[17][30] ),
    .I2(\dp.rf.rf[18][30] ),
    .I3(\dp.rf.rf[19][30] ),
    .S0(net13),
    .S1(net14),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_645_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_645_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_642_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_642_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_641_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_641_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05801_ (.I0(\dp.rf.rf[28][30] ),
    .I1(\dp.rf.rf[29][30] ),
    .I2(\dp.rf.rf[30][30] ),
    .I3(\dp.rf.rf[31][30] ),
    .S0(net13),
    .S1(net14),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05802_ (.I0(\dp.rf.rf[20][30] ),
    .I1(\dp.rf.rf[21][30] ),
    .I2(\dp.rf.rf[22][30] ),
    .I3(\dp.rf.rf[23][30] ),
    .S0(net13),
    .S1(net14),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_640_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_640_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_639_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_639_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05805_ (.I0(_01333_),
    .I1(_01334_),
    .I2(_01338_),
    .I3(_01339_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05806_ (.I0(\dp.rf.rf[8][30] ),
    .I1(\dp.rf.rf[9][30] ),
    .I2(\dp.rf.rf[10][30] ),
    .I3(\dp.rf.rf[11][30] ),
    .S0(net13),
    .S1(net14),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05807_ (.I0(\dp.rf.rf[0][30] ),
    .I1(\dp.rf.rf[1][30] ),
    .I2(\dp.rf.rf[2][30] ),
    .I3(\dp.rf.rf[3][30] ),
    .S0(net13),
    .S1(net14),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05808_ (.I0(\dp.rf.rf[12][30] ),
    .I1(\dp.rf.rf[13][30] ),
    .I2(\dp.rf.rf[14][30] ),
    .I3(\dp.rf.rf[15][30] ),
    .S0(net13),
    .S1(net14),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05809_ (.I0(\dp.rf.rf[4][30] ),
    .I1(\dp.rf.rf[5][30] ),
    .I2(\dp.rf.rf[6][30] ),
    .I3(\dp.rf.rf[7][30] ),
    .S0(net13),
    .S1(net14),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05810_ (.I0(_01343_),
    .I1(_01344_),
    .I2(_01345_),
    .I3(_01346_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_638_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_638_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05812_ (.I0(_01342_),
    .I1(_01347_),
    .S(_01064_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05813_ (.A1(_01329_),
    .A2(_01349_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05814_ (.A1(_01311_),
    .A2(_01350_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05815_ (.A1(_01119_),
    .A2(_05477_[0]),
    .B(_01351_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05816_ (.A1(net511),
    .A2(_01352_),
    .Z(_05120_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05817_ (.I(_05120_[0]),
    .ZN(_05124_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_637_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_637_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_633_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_633_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_632_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_632_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05821_ (.I0(\dp.rf.rf[8][30] ),
    .I1(\dp.rf.rf[9][30] ),
    .I2(\dp.rf.rf[12][30] ),
    .I3(\dp.rf.rf[13][30] ),
    .S0(net7),
    .S1(net537),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_631_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_631_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_630_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_630_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05824_ (.I0(\dp.rf.rf[10][30] ),
    .I1(\dp.rf.rf[11][30] ),
    .S(net7),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05825_ (.I(_01359_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05826_ (.I0(\dp.rf.rf[14][30] ),
    .I1(\dp.rf.rf[15][30] ),
    .S(net543),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05827_ (.I(_01361_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_629_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_629_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_628_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_628_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05830_ (.A1(net521),
    .A2(_01360_),
    .B1(_01362_),
    .B2(net537),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05831_ (.I0(_01356_),
    .I1(_01365_),
    .S(net8),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_626_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_626_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05833_ (.A1(net533),
    .A2(net532),
    .A3(_01125_),
    .B(net7),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_624_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_624_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05835_ (.A1(\dp.rf.rf[2][30] ),
    .A2(_01368_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_623_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_623_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_622_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_622_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05838_ (.A1(\dp.rf.rf[3][30] ),
    .A2(net543),
    .B1(net537),
    .B2(net165),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05839_ (.I0(\dp.rf.rf[6][30] ),
    .I1(\dp.rf.rf[7][30] ),
    .S(net543),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05840_ (.A1(_01167_),
    .A2(_01374_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05841_ (.A1(_01370_),
    .A2(_01373_),
    .B(net523),
    .C(_01375_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05842_ (.A1(_01144_),
    .A2(net526),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_618_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_618_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_616_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_616_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05845_ (.I0(\dp.rf.rf[1][30] ),
    .I1(\dp.rf.rf[5][30] ),
    .S(net537),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_614_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_614_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_611_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_611_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05848_ (.A1(\dp.rf.rf[4][30] ),
    .A2(net520),
    .B1(_01380_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _05849_ (.A1(net7),
    .A2(net9),
    .A3(net10),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _05850_ (.A1(_01030_),
    .A2(_01101_),
    .A3(_01125_),
    .B(_01384_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_609_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_609_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05852_ (.I(\dp.rf.rf[0][30] ),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05853_ (.A1(_01377_),
    .A2(_01383_),
    .B1(_01385_),
    .B2(_01387_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_608_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_608_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_598_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_598_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05856_ (.A1(_01167_),
    .A2(net530),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05857_ (.A1(_01144_),
    .A2(_01391_),
    .B(_01165_),
    .C(net11),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05858_ (.A1(net519),
    .A2(_01366_),
    .B1(_01376_),
    .B2(_01388_),
    .C(_01392_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05859_ (.I0(\dp.rf.rf[24][30] ),
    .I1(\dp.rf.rf[25][30] ),
    .I2(\dp.rf.rf[28][30] ),
    .I3(\dp.rf.rf[29][30] ),
    .S0(net543),
    .S1(net537),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05860_ (.I0(\dp.rf.rf[26][30] ),
    .I1(\dp.rf.rf[27][30] ),
    .S(net543),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05861_ (.I(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05862_ (.I0(\dp.rf.rf[30][30] ),
    .I1(\dp.rf.rf[31][30] ),
    .S(net543),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05863_ (.I(_01397_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05864_ (.A1(net521),
    .A2(_01396_),
    .B1(_01398_),
    .B2(net537),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_597_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_597_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05866_ (.I0(_01394_),
    .I1(_01399_),
    .S(net8),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05867_ (.A1(\dp.rf.rf[18][30] ),
    .A2(_01368_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05868_ (.A1(\dp.rf.rf[19][30] ),
    .A2(net543),
    .B1(net537),
    .B2(net165),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05869_ (.I0(\dp.rf.rf[22][30] ),
    .I1(\dp.rf.rf[23][30] ),
    .S(net543),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05870_ (.A1(_01167_),
    .A2(_01404_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _05871_ (.A1(_01402_),
    .A2(_01403_),
    .B(net523),
    .C(_01405_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05872_ (.I(\dp.rf.rf[16][30] ),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_596_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_596_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05874_ (.I0(\dp.rf.rf[17][30] ),
    .I1(\dp.rf.rf[21][30] ),
    .S(net537),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_595_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_595_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05876_ (.A1(\dp.rf.rf[20][30] ),
    .A2(_01245_),
    .B1(_01409_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05877_ (.A1(_01407_),
    .A2(_01385_),
    .B1(_01411_),
    .B2(_01377_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05878_ (.A1(net519),
    .A2(_01401_),
    .B1(_01406_),
    .B2(_01412_),
    .C(net517),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05879_ (.A1(_01393_),
    .A2(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _05880_ (.I(_01414_),
    .ZN(_05123_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05881_ (.A1(net22),
    .A2(_01165_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05882_ (.A1(_01320_),
    .A2(_01415_),
    .B(_01325_),
    .ZN(_05473_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_592_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_592_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_591_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_591_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_590_clk (.I(clknet_6_15__leaf_clk),
    .Z(clknet_leaf_590_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_588_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_588_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05887_ (.I0(\dp.rf.rf[24][29] ),
    .I1(\dp.rf.rf[25][29] ),
    .I2(\dp.rf.rf[26][29] ),
    .I3(\dp.rf.rf[27][29] ),
    .S0(net549),
    .S1(net14),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05888_ (.I0(\dp.rf.rf[16][29] ),
    .I1(\dp.rf.rf[17][29] ),
    .I2(\dp.rf.rf[18][29] ),
    .I3(\dp.rf.rf[19][29] ),
    .S0(net13),
    .S1(net14),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_587_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_587_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_584_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_584_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05891_ (.I0(\dp.rf.rf[28][29] ),
    .I1(\dp.rf.rf[29][29] ),
    .I2(\dp.rf.rf[30][29] ),
    .I3(\dp.rf.rf[31][29] ),
    .S0(net549),
    .S1(net14),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05892_ (.I0(\dp.rf.rf[20][29] ),
    .I1(\dp.rf.rf[21][29] ),
    .I2(\dp.rf.rf[22][29] ),
    .I3(\dp.rf.rf[23][29] ),
    .S0(net13),
    .S1(net14),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_581_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_581_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_578_clk (.I(clknet_6_15__leaf_clk),
    .Z(clknet_leaf_578_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_572_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_572_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05896_ (.I0(_01420_),
    .I1(_01421_),
    .I2(_01424_),
    .I3(_01425_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05897_ (.I0(\dp.rf.rf[8][29] ),
    .I1(\dp.rf.rf[9][29] ),
    .I2(\dp.rf.rf[10][29] ),
    .I3(\dp.rf.rf[11][29] ),
    .S0(net551),
    .S1(net14),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05898_ (.I0(\dp.rf.rf[0][29] ),
    .I1(\dp.rf.rf[1][29] ),
    .I2(\dp.rf.rf[2][29] ),
    .I3(\dp.rf.rf[3][29] ),
    .S0(net551),
    .S1(net14),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05899_ (.I0(\dp.rf.rf[12][29] ),
    .I1(\dp.rf.rf[13][29] ),
    .I2(\dp.rf.rf[14][29] ),
    .I3(\dp.rf.rf[15][29] ),
    .S0(net551),
    .S1(net14),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05900_ (.I0(\dp.rf.rf[4][29] ),
    .I1(\dp.rf.rf[5][29] ),
    .I2(\dp.rf.rf[6][29] ),
    .I3(\dp.rf.rf[7][29] ),
    .S0(net551),
    .S1(net14),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_570_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_570_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05902_ (.I0(_01430_),
    .I1(_01431_),
    .I2(_01432_),
    .I3(_01433_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05903_ (.I0(_01429_),
    .I1(_01435_),
    .S(_01064_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05904_ (.A1(_01329_),
    .A2(_01436_),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05905_ (.A1(_01311_),
    .A2(_01437_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05906_ (.A1(_01119_),
    .A2(_05473_[0]),
    .B(_01438_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05907_ (.A1(net511),
    .A2(_01439_),
    .Z(_05128_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05908_ (.I(_05128_[0]),
    .ZN(_05132_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05909_ (.A1(net166),
    .A2(_01278_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05910_ (.I0(\dp.rf.rf[10][29] ),
    .I1(\dp.rf.rf[11][29] ),
    .I2(\dp.rf.rf[14][29] ),
    .I3(\dp.rf.rf[15][29] ),
    .S0(net7),
    .S1(net9),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_569_clk (.I(clknet_6_24__leaf_clk),
    .Z(clknet_leaf_569_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05912_ (.I0(\dp.rf.rf[8][29] ),
    .I1(\dp.rf.rf[9][29] ),
    .I2(\dp.rf.rf[12][29] ),
    .I3(\dp.rf.rf[13][29] ),
    .S0(net7),
    .S1(net9),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05913_ (.I0(_01441_),
    .I1(_01443_),
    .S(_01140_),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05914_ (.A1(_01440_),
    .A2(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_562_clk (.I(clknet_6_19__leaf_clk),
    .Z(clknet_leaf_562_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_561_clk (.I(clknet_6_24__leaf_clk),
    .Z(clknet_leaf_561_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05917_ (.I0(\dp.rf.rf[2][29] ),
    .I1(\dp.rf.rf[3][29] ),
    .I2(\dp.rf.rf[6][29] ),
    .I3(\dp.rf.rf[7][29] ),
    .S0(net7),
    .S1(net537),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05918_ (.A1(net8),
    .A2(_01448_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05919_ (.I(\dp.rf.rf[4][29] ),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05920_ (.A1(_01148_),
    .A2(net9),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05921_ (.I(\dp.rf.rf[1][29] ),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05922_ (.I(\dp.rf.rf[5][29] ),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05923_ (.I0(_01452_),
    .I1(_01453_),
    .S(net537),
    .Z(_01454_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_557_clk (.I(clknet_6_24__leaf_clk),
    .Z(clknet_leaf_557_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_546_clk (.I(clknet_6_19__leaf_clk),
    .Z(clknet_leaf_546_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _05926_ (.A1(_01450_),
    .A2(_01451_),
    .B1(_01454_),
    .B2(net7),
    .C(net8),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _05927_ (.A1(_01212_),
    .A2(net167),
    .A3(_01198_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_545_clk (.I(clknet_6_19__leaf_clk),
    .Z(clknet_leaf_545_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05929_ (.A1(_01449_),
    .A2(_01457_),
    .B(_01458_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05930_ (.A1(_01445_),
    .A2(_01460_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05931_ (.I0(\dp.rf.rf[22][29] ),
    .I1(\dp.rf.rf[23][29] ),
    .S(net543),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05932_ (.A1(\dp.rf.rf[18][29] ),
    .A2(_01368_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05933_ (.I(\dp.rf.rf[19][29] ),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _05934_ (.A1(_01464_),
    .A2(_01148_),
    .B(net521),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05935_ (.A1(_01167_),
    .A2(_01462_),
    .B1(_01463_),
    .B2(_01465_),
    .C(_01284_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _05936_ (.A1(net167),
    .A2(_01384_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_536_clk (.I(clknet_6_19__leaf_clk),
    .Z(clknet_leaf_536_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05938_ (.I(\dp.rf.rf[20][29] ),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05939_ (.I(\dp.rf.rf[17][29] ),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05940_ (.I(\dp.rf.rf[21][29] ),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05941_ (.I0(_01470_),
    .I1(_01471_),
    .S(net537),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _05942_ (.A1(_01469_),
    .A2(_01451_),
    .B1(_01472_),
    .B2(net543),
    .C(net8),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _05943_ (.A1(\dp.rf.rf[16][29] ),
    .A2(_01467_),
    .B1(_01473_),
    .B2(_01177_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _05944_ (.A1(net11),
    .A2(_01126_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05945_ (.I0(\dp.rf.rf[26][29] ),
    .I1(\dp.rf.rf[27][29] ),
    .I2(\dp.rf.rf[30][29] ),
    .I3(\dp.rf.rf[31][29] ),
    .S0(net7),
    .S1(net9),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05946_ (.I0(\dp.rf.rf[24][29] ),
    .I1(\dp.rf.rf[25][29] ),
    .I2(\dp.rf.rf[28][29] ),
    .I3(\dp.rf.rf[29][29] ),
    .S0(net7),
    .S1(net9),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05947_ (.I0(_01476_),
    .I1(_01477_),
    .S(_01140_),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05948_ (.A1(_01144_),
    .A2(_01478_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _05949_ (.A1(_01466_),
    .A2(_01474_),
    .B(net515),
    .C(_01479_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _05950_ (.A1(_01461_),
    .A2(_01480_),
    .Z(_05127_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _05951_ (.I(_05127_[0]),
    .ZN(_05131_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_534_clk (.I(clknet_6_18__leaf_clk),
    .Z(clknet_leaf_534_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_533_clk (.I(clknet_6_18__leaf_clk),
    .Z(clknet_leaf_533_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_530_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_530_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05955_ (.I0(\dp.rf.rf[28][28] ),
    .I1(\dp.rf.rf[29][28] ),
    .I2(\dp.rf.rf[30][28] ),
    .I3(\dp.rf.rf[31][28] ),
    .S0(net548),
    .S1(net14),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05956_ (.I0(\dp.rf.rf[20][28] ),
    .I1(\dp.rf.rf[21][28] ),
    .I2(\dp.rf.rf[22][28] ),
    .I3(\dp.rf.rf[23][28] ),
    .S0(net548),
    .S1(net14),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_528_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_528_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05958_ (.I0(\dp.rf.rf[24][28] ),
    .I1(\dp.rf.rf[25][28] ),
    .I2(\dp.rf.rf[26][28] ),
    .I3(\dp.rf.rf[27][28] ),
    .S0(net548),
    .S1(net14),
    .Z(_01487_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05959_ (.I0(\dp.rf.rf[16][28] ),
    .I1(\dp.rf.rf[17][28] ),
    .I2(\dp.rf.rf[18][28] ),
    .I3(\dp.rf.rf[19][28] ),
    .S0(net13),
    .S1(net14),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_526_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_526_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05961_ (.I0(_01484_),
    .I1(_01485_),
    .I2(_01487_),
    .I3(_01488_),
    .S0(_01066_),
    .S1(_01055_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05962_ (.A1(_01064_),
    .A2(_01490_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_516_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_516_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05964_ (.I0(\dp.rf.rf[12][28] ),
    .I1(\dp.rf.rf[13][28] ),
    .I2(\dp.rf.rf[14][28] ),
    .I3(\dp.rf.rf[15][28] ),
    .S0(net13),
    .S1(net14),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05965_ (.I0(\dp.rf.rf[8][28] ),
    .I1(\dp.rf.rf[9][28] ),
    .I2(\dp.rf.rf[10][28] ),
    .I3(\dp.rf.rf[11][28] ),
    .S0(net13),
    .S1(net14),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05966_ (.I0(_01493_),
    .I1(_01494_),
    .S(_01055_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05967_ (.I0(\dp.rf.rf[4][28] ),
    .I1(\dp.rf.rf[5][28] ),
    .I2(\dp.rf.rf[6][28] ),
    .I3(\dp.rf.rf[7][28] ),
    .S0(net548),
    .S1(net14),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05968_ (.I0(\dp.rf.rf[0][28] ),
    .I1(\dp.rf.rf[1][28] ),
    .I2(\dp.rf.rf[2][28] ),
    .I3(\dp.rf.rf[3][28] ),
    .S0(net548),
    .S1(net14),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05969_ (.I0(_01496_),
    .I1(_01497_),
    .S(_01055_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _05970_ (.A1(_01084_),
    .A2(_01495_),
    .B1(_01498_),
    .B2(_01067_),
    .C(_01329_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _05971_ (.A1(_01491_),
    .A2(_01499_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05972_ (.A1(net21),
    .A2(_01165_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05973_ (.A1(_01320_),
    .A2(_01501_),
    .B(_01325_),
    .ZN(_05469_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05974_ (.A1(_01119_),
    .A2(_05469_[0]),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05975_ (.A1(_01311_),
    .A2(_01500_),
    .B(_01502_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _05976_ (.A1(net511),
    .A2(_01503_),
    .Z(_05136_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05977_ (.I(_05136_[0]),
    .ZN(_05140_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_515_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_515_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05979_ (.I0(\dp.rf.rf[22][28] ),
    .I1(\dp.rf.rf[23][28] ),
    .S(net544),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05980_ (.I(_01505_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _05981_ (.A1(net536),
    .A2(_01506_),
    .B(net523),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05982_ (.I(\dp.rf.rf[18][28] ),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _05983_ (.A1(_01508_),
    .A2(net533),
    .A3(net532),
    .A4(_01125_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05984_ (.I0(\dp.rf.rf[18][28] ),
    .I1(\dp.rf.rf[19][28] ),
    .S(net543),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05985_ (.I(_01510_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _05986_ (.A1(net521),
    .A2(_01509_),
    .A3(_01511_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_513_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_513_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _05988_ (.I0(\dp.rf.rf[17][28] ),
    .I1(\dp.rf.rf[21][28] ),
    .S(net536),
    .Z(_01514_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _05989_ (.A1(_01148_),
    .A2(_01514_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_509_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_509_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_507_clk (.I(clknet_6_16__leaf_clk),
    .Z(clknet_leaf_507_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _05992_ (.A1(\dp.rf.rf[20][28] ),
    .A2(net544),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_505_clk (.I(clknet_6_16__leaf_clk),
    .Z(clknet_leaf_505_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _05994_ (.A1(_01515_),
    .A2(_01518_),
    .B(_01144_),
    .C(net165),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _05995_ (.I(\dp.rf.rf[16][28] ),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _05996_ (.A1(_01521_),
    .A2(_01385_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _05997_ (.A1(_01507_),
    .A2(_01512_),
    .B1(_01520_),
    .B2(_01522_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _05998_ (.I0(\dp.rf.rf[26][28] ),
    .I1(\dp.rf.rf[27][28] ),
    .I2(\dp.rf.rf[30][28] ),
    .I3(\dp.rf.rf[31][28] ),
    .S0(net544),
    .S1(net535),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _05999_ (.A1(net8),
    .A2(_01524_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06000_ (.I0(\dp.rf.rf[24][28] ),
    .I1(\dp.rf.rf[28][28] ),
    .S(net535),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06001_ (.A1(net530),
    .A2(_01526_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_502_clk (.I(clknet_6_16__leaf_clk),
    .Z(clknet_leaf_502_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_497_clk (.I(clknet_6_17__leaf_clk),
    .Z(clknet_leaf_497_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06004_ (.I0(\dp.rf.rf[25][28] ),
    .I1(\dp.rf.rf[29][28] ),
    .S(net535),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06005_ (.A1(net544),
    .A2(_01140_),
    .A3(_01530_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06006_ (.A1(net519),
    .A2(_01527_),
    .A3(_01531_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06007_ (.A1(_01525_),
    .A2(_01532_),
    .B(net517),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06008_ (.A1(net8),
    .A2(_01231_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06009_ (.A1(net526),
    .A2(_01534_),
    .Z(_01535_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_496_clk (.I(clknet_6_17__leaf_clk),
    .Z(clknet_leaf_496_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_494_clk (.I(clknet_6_17__leaf_clk),
    .Z(clknet_leaf_494_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_493_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_493_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06013_ (.I0(\dp.rf.rf[2][28] ),
    .I1(\dp.rf.rf[3][28] ),
    .I2(\dp.rf.rf[6][28] ),
    .I3(\dp.rf.rf[7][28] ),
    .S0(net544),
    .S1(net535),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06014_ (.I(\dp.rf.rf[4][28] ),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_492_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_492_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06016_ (.I0(\dp.rf.rf[1][28] ),
    .I1(\dp.rf.rf[5][28] ),
    .S(net535),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06017_ (.A1(_01148_),
    .A2(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06018_ (.A1(_01540_),
    .A2(_01451_),
    .B(_01543_),
    .C(net8),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06019_ (.I0(\dp.rf.rf[10][28] ),
    .I1(\dp.rf.rf[11][28] ),
    .I2(\dp.rf.rf[14][28] ),
    .I3(\dp.rf.rf[15][28] ),
    .S0(net544),
    .S1(net535),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06020_ (.I0(\dp.rf.rf[8][28] ),
    .I1(\dp.rf.rf[9][28] ),
    .I2(\dp.rf.rf[12][28] ),
    .I3(\dp.rf.rf[13][28] ),
    .S0(net544),
    .S1(net535),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06021_ (.I0(_01545_),
    .I1(_01546_),
    .S(_01140_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06022_ (.A1(net527),
    .A2(_01278_),
    .A3(_01547_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06023_ (.A1(_01535_),
    .A2(_01539_),
    .B1(_01544_),
    .B2(_01458_),
    .C(_01548_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06024_ (.A1(_01523_),
    .A2(_01533_),
    .B(_01549_),
    .ZN(_05135_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06025_ (.I(_05135_[0]),
    .ZN(_05139_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06026_ (.A1(net20),
    .A2(_01165_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06027_ (.A1(_01320_),
    .A2(_01550_),
    .B(_01325_),
    .ZN(_05465_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_491_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_491_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06029_ (.I0(\dp.rf.rf[24][27] ),
    .I1(\dp.rf.rf[25][27] ),
    .I2(\dp.rf.rf[26][27] ),
    .I3(\dp.rf.rf[27][27] ),
    .S0(net550),
    .S1(net14),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06030_ (.I0(\dp.rf.rf[16][27] ),
    .I1(\dp.rf.rf[17][27] ),
    .I2(\dp.rf.rf[18][27] ),
    .I3(\dp.rf.rf[19][27] ),
    .S0(net551),
    .S1(net14),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06031_ (.I0(_01552_),
    .I1(_01553_),
    .S(_01066_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06032_ (.I0(\dp.rf.rf[28][27] ),
    .I1(\dp.rf.rf[29][27] ),
    .I2(\dp.rf.rf[30][27] ),
    .I3(\dp.rf.rf[31][27] ),
    .S0(net550),
    .S1(net14),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06033_ (.I0(\dp.rf.rf[20][27] ),
    .I1(\dp.rf.rf[21][27] ),
    .I2(\dp.rf.rf[22][27] ),
    .I3(\dp.rf.rf[23][27] ),
    .S0(net551),
    .S1(net14),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06034_ (.I0(_01555_),
    .I1(_01556_),
    .S(_01066_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06035_ (.I0(_01554_),
    .I1(_01557_),
    .S(net15),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06036_ (.I0(\dp.rf.rf[8][27] ),
    .I1(\dp.rf.rf[9][27] ),
    .I2(\dp.rf.rf[10][27] ),
    .I3(\dp.rf.rf[11][27] ),
    .S0(net550),
    .S1(net14),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06037_ (.I0(\dp.rf.rf[0][27] ),
    .I1(\dp.rf.rf[1][27] ),
    .I2(\dp.rf.rf[2][27] ),
    .I3(\dp.rf.rf[3][27] ),
    .S0(net550),
    .S1(net14),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06038_ (.I0(_01559_),
    .I1(_01560_),
    .S(_01066_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06039_ (.I0(\dp.rf.rf[12][27] ),
    .I1(\dp.rf.rf[13][27] ),
    .I2(\dp.rf.rf[14][27] ),
    .I3(\dp.rf.rf[15][27] ),
    .S0(net550),
    .S1(net14),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06040_ (.I0(\dp.rf.rf[4][27] ),
    .I1(\dp.rf.rf[5][27] ),
    .I2(\dp.rf.rf[6][27] ),
    .I3(\dp.rf.rf[7][27] ),
    .S0(net550),
    .S1(net14),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06041_ (.I0(_01562_),
    .I1(_01563_),
    .S(_01066_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06042_ (.I0(_01561_),
    .I1(_01564_),
    .S(net15),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06043_ (.A1(net17),
    .A2(_01558_),
    .B1(_01565_),
    .B2(_01309_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06044_ (.A1(_01311_),
    .A2(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06045_ (.A1(_01311_),
    .A2(_05465_[0]),
    .B(_01567_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06046_ (.A1(net511),
    .A2(_01568_),
    .Z(_05144_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06047_ (.I(_05144_[0]),
    .ZN(_05148_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_488_clk (.I(clknet_6_17__leaf_clk),
    .Z(clknet_leaf_488_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_486_clk (.I(clknet_6_17__leaf_clk),
    .Z(clknet_leaf_486_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06050_ (.I0(\dp.rf.rf[18][27] ),
    .I1(\dp.rf.rf[19][27] ),
    .I2(\dp.rf.rf[22][27] ),
    .I3(\dp.rf.rf[23][27] ),
    .S0(net7),
    .S1(net536),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06051_ (.I0(\dp.rf.rf[17][27] ),
    .I1(\dp.rf.rf[21][27] ),
    .S(net536),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06052_ (.A1(_01148_),
    .A2(_01572_),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_484_clk (.I(clknet_6_22__leaf_clk),
    .Z(clknet_leaf_484_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06054_ (.A1(\dp.rf.rf[20][27] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06055_ (.A1(_01573_),
    .A2(_01575_),
    .B(_01144_),
    .C(net529),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06056_ (.I(\dp.rf.rf[16][27] ),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06057_ (.A1(_01577_),
    .A2(_01385_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06058_ (.A1(_01284_),
    .A2(_01571_),
    .B1(_01576_),
    .B2(_01578_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06059_ (.A1(net10),
    .A2(net166),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_481_clk (.I(clknet_6_22__leaf_clk),
    .Z(clknet_leaf_481_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06061_ (.I0(\dp.rf.rf[26][27] ),
    .I1(\dp.rf.rf[27][27] ),
    .I2(\dp.rf.rf[30][27] ),
    .I3(\dp.rf.rf[31][27] ),
    .S0(net7),
    .S1(net536),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06062_ (.A1(net8),
    .A2(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_473_clk (.I(clknet_6_23__leaf_clk),
    .Z(clknet_leaf_473_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06064_ (.A1(net7),
    .A2(_01140_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06065_ (.I0(\dp.rf.rf[25][27] ),
    .I1(\dp.rf.rf[29][27] ),
    .S(net536),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06066_ (.I0(\dp.rf.rf[24][27] ),
    .I1(\dp.rf.rf[28][27] ),
    .S(net536),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06067_ (.A1(_01585_),
    .A2(_01586_),
    .B1(_01587_),
    .B2(net530),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06068_ (.A1(_01580_),
    .A2(_01583_),
    .A3(_01588_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_469_clk (.I(clknet_6_21__leaf_clk),
    .Z(clknet_leaf_469_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06070_ (.A1(\dp.rf.rf[4][27] ),
    .A2(net7),
    .A3(_01167_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06071_ (.I0(\dp.rf.rf[1][27] ),
    .I1(\dp.rf.rf[5][27] ),
    .S(net9),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06072_ (.A1(_01148_),
    .A2(_01592_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06073_ (.I0(\dp.rf.rf[2][27] ),
    .I1(\dp.rf.rf[3][27] ),
    .I2(\dp.rf.rf[6][27] ),
    .I3(\dp.rf.rf[7][27] ),
    .S0(net7),
    .S1(net9),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06074_ (.A1(net8),
    .A2(_01594_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06075_ (.A1(net8),
    .A2(_01591_),
    .A3(_01593_),
    .B(_01595_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06076_ (.I0(\dp.rf.rf[10][27] ),
    .I1(\dp.rf.rf[11][27] ),
    .I2(\dp.rf.rf[14][27] ),
    .I3(\dp.rf.rf[15][27] ),
    .S0(net7),
    .S1(net9),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06077_ (.I0(\dp.rf.rf[8][27] ),
    .I1(\dp.rf.rf[9][27] ),
    .I2(\dp.rf.rf[12][27] ),
    .I3(\dp.rf.rf[13][27] ),
    .S0(net7),
    .S1(net9),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_468_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_468_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06079_ (.I0(_01597_),
    .I1(_01598_),
    .S(_01140_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06080_ (.A1(_01458_),
    .A2(_01596_),
    .B1(_01600_),
    .B2(_01440_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _06081_ (.A1(net515),
    .A2(_01579_),
    .A3(_01589_),
    .B(_01601_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_465_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_465_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06083_ (.I(_01602_),
    .ZN(_05147_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06084_ (.A1(net19),
    .A2(_01165_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06085_ (.A1(_01320_),
    .A2(_01603_),
    .B(_01325_),
    .ZN(_05461_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_459_clk (.I(clknet_6_23__leaf_clk),
    .Z(clknet_leaf_459_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_458_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_458_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_457_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_457_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_456_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_456_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_454_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_454_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06091_ (.I0(\dp.rf.rf[24][26] ),
    .I1(\dp.rf.rf[25][26] ),
    .I2(\dp.rf.rf[26][26] ),
    .I3(\dp.rf.rf[27][26] ),
    .S0(net13),
    .S1(net14),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06092_ (.I0(\dp.rf.rf[16][26] ),
    .I1(\dp.rf.rf[17][26] ),
    .I2(\dp.rf.rf[18][26] ),
    .I3(\dp.rf.rf[19][26] ),
    .S0(net13),
    .S1(net14),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_452_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_452_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_449_clk (.I(clknet_6_21__leaf_clk),
    .Z(clknet_leaf_449_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06095_ (.I0(\dp.rf.rf[28][26] ),
    .I1(\dp.rf.rf[29][26] ),
    .I2(\dp.rf.rf[30][26] ),
    .I3(\dp.rf.rf[31][26] ),
    .S0(net13),
    .S1(net14),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06096_ (.I0(\dp.rf.rf[20][26] ),
    .I1(\dp.rf.rf[21][26] ),
    .I2(\dp.rf.rf[22][26] ),
    .I3(\dp.rf.rf[23][26] ),
    .S0(net13),
    .S1(net14),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_448_clk (.I(clknet_6_23__leaf_clk),
    .Z(clknet_leaf_448_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06098_ (.I0(_01609_),
    .I1(_01610_),
    .I2(_01613_),
    .I3(_01614_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06099_ (.I0(\dp.rf.rf[8][26] ),
    .I1(\dp.rf.rf[9][26] ),
    .I2(\dp.rf.rf[10][26] ),
    .I3(\dp.rf.rf[11][26] ),
    .S0(net13),
    .S1(net14),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06100_ (.I0(\dp.rf.rf[0][26] ),
    .I1(\dp.rf.rf[1][26] ),
    .I2(\dp.rf.rf[2][26] ),
    .I3(\dp.rf.rf[3][26] ),
    .S0(net548),
    .S1(net14),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_446_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_446_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_442_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_442_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06103_ (.I0(\dp.rf.rf[12][26] ),
    .I1(\dp.rf.rf[13][26] ),
    .I2(\dp.rf.rf[14][26] ),
    .I3(\dp.rf.rf[15][26] ),
    .S0(net13),
    .S1(net14),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06104_ (.I0(\dp.rf.rf[4][26] ),
    .I1(\dp.rf.rf[5][26] ),
    .I2(\dp.rf.rf[6][26] ),
    .I3(\dp.rf.rf[7][26] ),
    .S0(net548),
    .S1(net14),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06105_ (.I0(_01617_),
    .I1(_01618_),
    .I2(_01621_),
    .I3(_01622_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_441_clk (.I(clknet_6_25__leaf_clk),
    .Z(clknet_leaf_441_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06107_ (.A1(net17),
    .A2(_01616_),
    .B1(_01623_),
    .B2(_01309_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06108_ (.I(_01625_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06109_ (.A1(_01311_),
    .A2(_01626_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06110_ (.A1(_01119_),
    .A2(_05461_[0]),
    .B(_01627_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06111_ (.A1(net511),
    .A2(_01628_),
    .Z(_05152_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06112_ (.I(_05152_[0]),
    .ZN(_05156_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06113_ (.I0(\dp.rf.rf[2][26] ),
    .I1(\dp.rf.rf[3][26] ),
    .I2(\dp.rf.rf[6][26] ),
    .I3(\dp.rf.rf[7][26] ),
    .S0(net544),
    .S1(net535),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06114_ (.I(_01629_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06115_ (.I0(\dp.rf.rf[1][26] ),
    .I1(\dp.rf.rf[5][26] ),
    .S(net535),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_438_clk (.I(clknet_6_25__leaf_clk),
    .Z(clknet_leaf_438_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06117_ (.A1(\dp.rf.rf[4][26] ),
    .A2(_01245_),
    .B1(_01631_),
    .B2(_01148_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06118_ (.I0(_01630_),
    .I1(_01633_),
    .S(_01140_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06119_ (.I0(\dp.rf.rf[10][26] ),
    .I1(\dp.rf.rf[11][26] ),
    .I2(\dp.rf.rf[14][26] ),
    .I3(\dp.rf.rf[15][26] ),
    .S0(net544),
    .S1(net535),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06120_ (.I0(\dp.rf.rf[8][26] ),
    .I1(\dp.rf.rf[9][26] ),
    .I2(\dp.rf.rf[12][26] ),
    .I3(\dp.rf.rf[13][26] ),
    .S0(net544),
    .S1(net535),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06121_ (.I0(_01635_),
    .I1(_01636_),
    .S(_01140_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06122_ (.A1(_01440_),
    .A2(_01637_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06123_ (.A1(net516),
    .A2(_01634_),
    .B(_01638_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_436_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_436_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06125_ (.I0(\dp.rf.rf[22][26] ),
    .I1(\dp.rf.rf[23][26] ),
    .S(net544),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06126_ (.A1(\dp.rf.rf[18][26] ),
    .A2(_01368_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06127_ (.A1(\dp.rf.rf[19][26] ),
    .A2(net543),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06128_ (.A1(net521),
    .A2(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06129_ (.A1(_01167_),
    .A2(_01641_),
    .B1(_01642_),
    .B2(_01644_),
    .C(_01284_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06130_ (.I(\dp.rf.rf[20][26] ),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06131_ (.I0(\dp.rf.rf[17][26] ),
    .I1(\dp.rf.rf[21][26] ),
    .S(net536),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06132_ (.A1(_01148_),
    .A2(_01647_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06133_ (.A1(_01646_),
    .A2(_01451_),
    .B(_01648_),
    .C(net8),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06134_ (.A1(\dp.rf.rf[16][26] ),
    .A2(_01467_),
    .B1(_01649_),
    .B2(_01177_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_432_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_432_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06136_ (.I0(\dp.rf.rf[26][26] ),
    .I1(\dp.rf.rf[27][26] ),
    .I2(\dp.rf.rf[30][26] ),
    .I3(\dp.rf.rf[31][26] ),
    .S0(net7),
    .S1(net535),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06137_ (.I0(\dp.rf.rf[24][26] ),
    .I1(\dp.rf.rf[25][26] ),
    .I2(\dp.rf.rf[28][26] ),
    .I3(\dp.rf.rf[29][26] ),
    .S0(net7),
    .S1(net535),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06138_ (.I0(_01652_),
    .I1(_01653_),
    .S(_01140_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06139_ (.A1(_01144_),
    .A2(_01654_),
    .B(net517),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06140_ (.A1(_01645_),
    .A2(_01650_),
    .B(_01655_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06141_ (.A1(_01639_),
    .A2(_01656_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_430_clk (.I(clknet_6_30__leaf_clk),
    .Z(clknet_leaf_430_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06143_ (.I(_01657_),
    .ZN(_05155_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06144_ (.A1(net18),
    .A2(_01165_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06145_ (.A1(_01320_),
    .A2(_01658_),
    .B(_01325_),
    .ZN(_05457_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06146_ (.I(\dp.rf.rf[28][25] ),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06147_ (.I(\dp.rf.rf[29][25] ),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06148_ (.I(\dp.rf.rf[30][25] ),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06149_ (.I(\dp.rf.rf[31][25] ),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06150_ (.I0(_01659_),
    .I1(_01660_),
    .I2(_01661_),
    .I3(_01662_),
    .S0(net549),
    .S1(net14),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06151_ (.I(\dp.rf.rf[20][25] ),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06152_ (.I(\dp.rf.rf[21][25] ),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06153_ (.I(\dp.rf.rf[22][25] ),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06154_ (.I(\dp.rf.rf[23][25] ),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06155_ (.I0(_01664_),
    .I1(_01665_),
    .I2(_01666_),
    .I3(_01667_),
    .S0(net13),
    .S1(net14),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06156_ (.I(\dp.rf.rf[24][25] ),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06157_ (.I(\dp.rf.rf[25][25] ),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06158_ (.I(\dp.rf.rf[26][25] ),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06159_ (.I(\dp.rf.rf[27][25] ),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06160_ (.I0(_01669_),
    .I1(_01670_),
    .I2(_01671_),
    .I3(_01672_),
    .S0(net549),
    .S1(net14),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06161_ (.I(\dp.rf.rf[16][25] ),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06162_ (.I(\dp.rf.rf[17][25] ),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06163_ (.I(\dp.rf.rf[18][25] ),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06164_ (.I(\dp.rf.rf[19][25] ),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06165_ (.I0(_01674_),
    .I1(_01675_),
    .I2(_01676_),
    .I3(_01677_),
    .S0(net13),
    .S1(net14),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_427_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_427_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06167_ (.I0(_01663_),
    .I1(_01668_),
    .I2(_01673_),
    .I3(_01678_),
    .S0(_01066_),
    .S1(_01055_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06168_ (.A1(net17),
    .A2(_01680_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06169_ (.I0(\dp.rf.rf[4][25] ),
    .I1(\dp.rf.rf[5][25] ),
    .I2(\dp.rf.rf[6][25] ),
    .I3(\dp.rf.rf[7][25] ),
    .S0(net551),
    .S1(net14),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06170_ (.I0(\dp.rf.rf[0][25] ),
    .I1(\dp.rf.rf[1][25] ),
    .I2(\dp.rf.rf[2][25] ),
    .I3(\dp.rf.rf[3][25] ),
    .S0(net551),
    .S1(net14),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_425_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_425_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06172_ (.I0(_01682_),
    .I1(_01683_),
    .S(_01055_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06173_ (.A1(_01067_),
    .A2(_01685_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_424_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_424_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_423_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_423_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06176_ (.I0(\dp.rf.rf[12][25] ),
    .I1(\dp.rf.rf[13][25] ),
    .I2(\dp.rf.rf[14][25] ),
    .I3(\dp.rf.rf[15][25] ),
    .S0(net550),
    .S1(net14),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06177_ (.I0(\dp.rf.rf[8][25] ),
    .I1(\dp.rf.rf[9][25] ),
    .I2(\dp.rf.rf[10][25] ),
    .I3(\dp.rf.rf[11][25] ),
    .S0(net550),
    .S1(net14),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06178_ (.I0(_01689_),
    .I1(_01690_),
    .S(_01055_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06179_ (.A1(_01084_),
    .A2(_01691_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _06180_ (.A1(_01329_),
    .A2(_01681_),
    .A3(_01686_),
    .A4(_01692_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06181_ (.A1(_01311_),
    .A2(_01693_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06182_ (.A1(_01119_),
    .A2(_05457_[0]),
    .B(_01694_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06183_ (.A1(net511),
    .A2(_01695_),
    .Z(_05160_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06184_ (.I(_05160_[0]),
    .ZN(_05164_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06185_ (.I(_01440_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06186_ (.A1(net7),
    .A2(net8),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_421_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_421_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06188_ (.I0(\dp.rf.rf[11][25] ),
    .I1(\dp.rf.rf[15][25] ),
    .S(net536),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_419_clk (.I(clknet_6_31__leaf_clk),
    .Z(clknet_leaf_419_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06190_ (.I0(\dp.rf.rf[10][25] ),
    .I1(\dp.rf.rf[14][25] ),
    .S(net536),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06191_ (.A1(_01148_),
    .A2(net8),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06192_ (.I0(\dp.rf.rf[8][25] ),
    .I1(\dp.rf.rf[9][25] ),
    .I2(\dp.rf.rf[12][25] ),
    .I3(\dp.rf.rf[13][25] ),
    .S0(net7),
    .S1(net536),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06193_ (.A1(_01140_),
    .A2(_01703_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06194_ (.A1(_01697_),
    .A2(_01699_),
    .B1(_01701_),
    .B2(_01702_),
    .C(_01704_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06195_ (.I0(\dp.rf.rf[2][25] ),
    .I1(\dp.rf.rf[3][25] ),
    .I2(\dp.rf.rf[6][25] ),
    .I3(\dp.rf.rf[7][25] ),
    .S0(net7),
    .S1(net537),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06196_ (.I(\dp.rf.rf[4][25] ),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06197_ (.I(\dp.rf.rf[1][25] ),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06198_ (.I(\dp.rf.rf[5][25] ),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06199_ (.I0(_01708_),
    .I1(_01709_),
    .S(net537),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06200_ (.A1(_01707_),
    .A2(_01451_),
    .B1(_01710_),
    .B2(net7),
    .C(net8),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06201_ (.A1(net8),
    .A2(_01706_),
    .B(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _06202_ (.A1(_01696_),
    .A2(_01705_),
    .B1(_01712_),
    .B2(net516),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06203_ (.I0(\dp.rf.rf[22][25] ),
    .I1(\dp.rf.rf[23][25] ),
    .S(net543),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06204_ (.A1(\dp.rf.rf[18][25] ),
    .A2(_01368_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06205_ (.A1(_01677_),
    .A2(_01148_),
    .B(net521),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06206_ (.A1(_01167_),
    .A2(_01714_),
    .B1(_01715_),
    .B2(_01716_),
    .C(_01284_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06207_ (.I0(_01675_),
    .I1(_01665_),
    .S(net537),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06208_ (.A1(_01664_),
    .A2(_01451_),
    .B1(_01718_),
    .B2(net543),
    .C(net8),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06209_ (.A1(\dp.rf.rf[16][25] ),
    .A2(_01467_),
    .B1(_01719_),
    .B2(_01177_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06210_ (.I0(\dp.rf.rf[26][25] ),
    .I1(\dp.rf.rf[27][25] ),
    .I2(\dp.rf.rf[30][25] ),
    .I3(\dp.rf.rf[31][25] ),
    .S0(net541),
    .S1(net9),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06211_ (.I0(\dp.rf.rf[24][25] ),
    .I1(\dp.rf.rf[25][25] ),
    .I2(\dp.rf.rf[28][25] ),
    .I3(\dp.rf.rf[29][25] ),
    .S0(net541),
    .S1(net9),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06212_ (.I0(_01721_),
    .I1(_01722_),
    .S(_01140_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06213_ (.A1(_01144_),
    .A2(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _06214_ (.A1(_01717_),
    .A2(_01720_),
    .B(net515),
    .C(_01724_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06215_ (.A1(_01713_),
    .A2(_01725_),
    .Z(_05159_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06216_ (.I(_05159_[0]),
    .ZN(_05163_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_418_clk (.I(clknet_6_31__leaf_clk),
    .Z(clknet_leaf_418_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_413_clk (.I(clknet_6_30__leaf_clk),
    .Z(clknet_leaf_413_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06219_ (.I0(\dp.rf.rf[24][24] ),
    .I1(\dp.rf.rf[25][24] ),
    .I2(\dp.rf.rf[26][24] ),
    .I3(\dp.rf.rf[27][24] ),
    .S0(net13),
    .S1(net14),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06220_ (.I0(\dp.rf.rf[16][24] ),
    .I1(\dp.rf.rf[17][24] ),
    .I2(\dp.rf.rf[18][24] ),
    .I3(\dp.rf.rf[19][24] ),
    .S0(net13),
    .S1(net14),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06221_ (.I0(_01728_),
    .I1(_01729_),
    .S(_01066_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06222_ (.I0(\dp.rf.rf[28][24] ),
    .I1(\dp.rf.rf[29][24] ),
    .I2(\dp.rf.rf[30][24] ),
    .I3(\dp.rf.rf[31][24] ),
    .S0(net13),
    .S1(net14),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06223_ (.I0(\dp.rf.rf[20][24] ),
    .I1(\dp.rf.rf[21][24] ),
    .I2(\dp.rf.rf[22][24] ),
    .I3(\dp.rf.rf[23][24] ),
    .S0(net548),
    .S1(net14),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06224_ (.I0(_01731_),
    .I1(_01732_),
    .S(_01066_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06225_ (.A1(net15),
    .A2(_01733_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06226_ (.A1(_01055_),
    .A2(_01730_),
    .B(_01734_),
    .C(_01064_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06227_ (.I0(\dp.rf.rf[12][24] ),
    .I1(\dp.rf.rf[13][24] ),
    .I2(\dp.rf.rf[14][24] ),
    .I3(\dp.rf.rf[15][24] ),
    .S0(net548),
    .S1(net14),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06228_ (.I0(\dp.rf.rf[8][24] ),
    .I1(\dp.rf.rf[9][24] ),
    .I2(\dp.rf.rf[10][24] ),
    .I3(\dp.rf.rf[11][24] ),
    .S0(net548),
    .S1(net14),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06229_ (.I0(_01736_),
    .I1(_01737_),
    .S(_01055_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06230_ (.I0(\dp.rf.rf[4][24] ),
    .I1(\dp.rf.rf[5][24] ),
    .I2(\dp.rf.rf[6][24] ),
    .I3(\dp.rf.rf[7][24] ),
    .S0(net548),
    .S1(net14),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06231_ (.I0(\dp.rf.rf[0][24] ),
    .I1(\dp.rf.rf[1][24] ),
    .I2(\dp.rf.rf[2][24] ),
    .I3(\dp.rf.rf[3][24] ),
    .S0(net548),
    .S1(net14),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06232_ (.I0(_01739_),
    .I1(_01740_),
    .S(_01055_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06233_ (.A1(_01084_),
    .A2(_01738_),
    .B1(_01741_),
    .B2(_01067_),
    .C(_01329_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06234_ (.A1(_01735_),
    .A2(_01742_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06235_ (.A1(net17),
    .A2(_01165_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06236_ (.A1(_01320_),
    .A2(_01744_),
    .B(_01325_),
    .ZN(_05453_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06237_ (.A1(_01119_),
    .A2(_05453_[0]),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06238_ (.A1(_01311_),
    .A2(_01743_),
    .B(_01745_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06239_ (.A1(net511),
    .A2(_01746_),
    .Z(_05168_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06240_ (.I(_05168_[0]),
    .ZN(_05172_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_411_clk (.I(clknet_6_31__leaf_clk),
    .Z(clknet_leaf_411_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06242_ (.I0(\dp.rf.rf[22][24] ),
    .I1(\dp.rf.rf[23][24] ),
    .S(net545),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06243_ (.I(_01748_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06244_ (.A1(net536),
    .A2(_01749_),
    .B(net523),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06245_ (.I(\dp.rf.rf[18][24] ),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _06246_ (.A1(_01751_),
    .A2(net533),
    .A3(net532),
    .A4(_01125_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06247_ (.I0(\dp.rf.rf[18][24] ),
    .I1(\dp.rf.rf[19][24] ),
    .S(net545),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06248_ (.I(_01753_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06249_ (.A1(net521),
    .A2(_01752_),
    .A3(_01754_),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_408_clk (.I(clknet_6_31__leaf_clk),
    .Z(clknet_leaf_408_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06251_ (.I0(\dp.rf.rf[17][24] ),
    .I1(\dp.rf.rf[21][24] ),
    .S(net535),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06252_ (.A1(_01148_),
    .A2(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_404_clk (.I(clknet_6_53__leaf_clk),
    .Z(clknet_leaf_404_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_403_clk (.I(clknet_6_30__leaf_clk),
    .Z(clknet_leaf_403_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_396_clk (.I(clknet_6_30__leaf_clk),
    .Z(clknet_leaf_396_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06256_ (.A1(\dp.rf.rf[20][24] ),
    .A2(net545),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_394_clk (.I(clknet_6_53__leaf_clk),
    .Z(clknet_leaf_394_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06258_ (.A1(_01758_),
    .A2(_01762_),
    .B(_01144_),
    .C(net529),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06259_ (.I(\dp.rf.rf[16][24] ),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_393_clk (.I(clknet_6_52__leaf_clk),
    .Z(clknet_leaf_393_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06261_ (.A1(_01765_),
    .A2(_01385_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06262_ (.A1(_01750_),
    .A2(_01755_),
    .B1(_01764_),
    .B2(_01767_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_390_clk (.I(clknet_6_52__leaf_clk),
    .Z(clknet_leaf_390_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06264_ (.I0(\dp.rf.rf[26][24] ),
    .I1(\dp.rf.rf[27][24] ),
    .I2(\dp.rf.rf[30][24] ),
    .I3(\dp.rf.rf[31][24] ),
    .S0(net545),
    .S1(net535),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06265_ (.A1(net8),
    .A2(_01770_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06266_ (.I0(\dp.rf.rf[24][24] ),
    .I1(\dp.rf.rf[28][24] ),
    .S(net535),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06267_ (.I0(\dp.rf.rf[25][24] ),
    .I1(\dp.rf.rf[29][24] ),
    .S(net535),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06268_ (.A1(net530),
    .A2(_01772_),
    .B1(_01773_),
    .B2(_01585_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06269_ (.A1(_01580_),
    .A2(_01771_),
    .A3(_01774_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06270_ (.I0(\dp.rf.rf[8][24] ),
    .I1(\dp.rf.rf[9][24] ),
    .I2(\dp.rf.rf[12][24] ),
    .I3(\dp.rf.rf[13][24] ),
    .S0(net544),
    .S1(net535),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06271_ (.I0(\dp.rf.rf[1][24] ),
    .I1(\dp.rf.rf[5][24] ),
    .S(net535),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06272_ (.A1(_01148_),
    .A2(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06273_ (.A1(\dp.rf.rf[4][24] ),
    .A2(net545),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01779_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06274_ (.A1(_01778_),
    .A2(_01779_),
    .B(net529),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _06275_ (.A1(net11),
    .A2(_01180_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06276_ (.I0(\dp.rf.rf[10][24] ),
    .I1(\dp.rf.rf[11][24] ),
    .I2(\dp.rf.rf[14][24] ),
    .I3(\dp.rf.rf[15][24] ),
    .S0(net544),
    .S1(net535),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06277_ (.I0(\dp.rf.rf[2][24] ),
    .I1(\dp.rf.rf[3][24] ),
    .I2(\dp.rf.rf[6][24] ),
    .I3(\dp.rf.rf[7][24] ),
    .S0(net545),
    .S1(net535),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06278_ (.I0(_01782_),
    .I1(_01783_),
    .S(_01144_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _06279_ (.A1(_01279_),
    .A2(_01776_),
    .B1(_01780_),
    .B2(_01458_),
    .C1(_01781_),
    .C2(_01784_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _06280_ (.A1(_01475_),
    .A2(_01768_),
    .A3(_01775_),
    .B(_01785_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_385_clk (.I(clknet_6_27__leaf_clk),
    .Z(clknet_leaf_385_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06282_ (.I(_01786_),
    .ZN(_05171_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06283_ (.A1(net16),
    .A2(_01165_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06284_ (.A1(_01320_),
    .A2(_01787_),
    .B(_01325_),
    .ZN(_05449_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06285_ (.I(\dp.rf.rf[24][23] ),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06286_ (.I(\dp.rf.rf[25][23] ),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06287_ (.I(\dp.rf.rf[26][23] ),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06288_ (.I(\dp.rf.rf[27][23] ),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_383_clk (.I(clknet_6_30__leaf_clk),
    .Z(clknet_leaf_383_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_380_clk (.I(clknet_6_27__leaf_clk),
    .Z(clknet_leaf_380_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06291_ (.I0(_01788_),
    .I1(_01789_),
    .I2(_01790_),
    .I3(_01791_),
    .S0(net549),
    .S1(net14),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06292_ (.I(\dp.rf.rf[16][23] ),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06293_ (.I(\dp.rf.rf[17][23] ),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06294_ (.I(\dp.rf.rf[18][23] ),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06295_ (.I(\dp.rf.rf[19][23] ),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06296_ (.I0(_01795_),
    .I1(_01796_),
    .I2(_01797_),
    .I3(_01798_),
    .S0(net549),
    .S1(net14),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06297_ (.I(\dp.rf.rf[28][23] ),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06298_ (.I(\dp.rf.rf[29][23] ),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06299_ (.I(\dp.rf.rf[30][23] ),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06300_ (.I(\dp.rf.rf[31][23] ),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06301_ (.I0(_01800_),
    .I1(_01801_),
    .I2(_01802_),
    .I3(_01803_),
    .S0(net549),
    .S1(net14),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06302_ (.I(\dp.rf.rf[20][23] ),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06303_ (.I(\dp.rf.rf[21][23] ),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06304_ (.I(\dp.rf.rf[22][23] ),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06305_ (.I(\dp.rf.rf[23][23] ),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06306_ (.I0(_01805_),
    .I1(_01806_),
    .I2(_01807_),
    .I3(_01808_),
    .S0(net549),
    .S1(net14),
    .Z(_01809_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_375_clk (.I(clknet_6_25__leaf_clk),
    .Z(clknet_leaf_375_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06308_ (.I0(_01794_),
    .I1(_01799_),
    .I2(_01804_),
    .I3(_01809_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_374_clk (.I(clknet_6_25__leaf_clk),
    .Z(clknet_leaf_374_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_372_clk (.I(clknet_6_25__leaf_clk),
    .Z(clknet_leaf_372_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06311_ (.I0(\dp.rf.rf[8][23] ),
    .I1(\dp.rf.rf[9][23] ),
    .I2(\dp.rf.rf[10][23] ),
    .I3(\dp.rf.rf[11][23] ),
    .S0(net550),
    .S1(net14),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06312_ (.I0(\dp.rf.rf[0][23] ),
    .I1(\dp.rf.rf[1][23] ),
    .I2(\dp.rf.rf[2][23] ),
    .I3(\dp.rf.rf[3][23] ),
    .S0(net550),
    .S1(net14),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06313_ (.I0(\dp.rf.rf[12][23] ),
    .I1(\dp.rf.rf[13][23] ),
    .I2(\dp.rf.rf[14][23] ),
    .I3(\dp.rf.rf[15][23] ),
    .S0(net550),
    .S1(net14),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06314_ (.I0(\dp.rf.rf[4][23] ),
    .I1(\dp.rf.rf[5][23] ),
    .I2(\dp.rf.rf[6][23] ),
    .I3(\dp.rf.rf[7][23] ),
    .S0(net550),
    .S1(net14),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06315_ (.I0(_01814_),
    .I1(_01815_),
    .I2(_01816_),
    .I3(_01817_),
    .S0(_01066_),
    .S1(net15),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06316_ (.A1(_01309_),
    .A2(_01818_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06317_ (.A1(_01064_),
    .A2(_01811_),
    .B(_01819_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _06318_ (.I(_01820_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06319_ (.A1(_01311_),
    .A2(_01821_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06320_ (.A1(_01311_),
    .A2(_05449_[0]),
    .B(_01822_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06321_ (.A1(net511),
    .A2(_01823_),
    .Z(_05176_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06322_ (.I(_05176_[0]),
    .ZN(_05180_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06323_ (.I0(\dp.rf.rf[18][23] ),
    .I1(\dp.rf.rf[19][23] ),
    .I2(\dp.rf.rf[22][23] ),
    .I3(\dp.rf.rf[23][23] ),
    .S0(net540),
    .S1(net9),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_370_clk (.I(clknet_6_24__leaf_clk),
    .Z(clknet_leaf_370_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06325_ (.I0(\dp.rf.rf[17][23] ),
    .I1(\dp.rf.rf[21][23] ),
    .S(net9),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06326_ (.I(_01826_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06327_ (.A1(_01805_),
    .A2(_01451_),
    .B1(_01827_),
    .B2(net540),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_369_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_369_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06329_ (.I0(_01824_),
    .I1(_01828_),
    .S(_01140_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06330_ (.A1(\dp.rf.rf[18][23] ),
    .A2(net8),
    .B(\dp.rf.rf[16][23] ),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06331_ (.A1(_01168_),
    .A2(_01831_),
    .B(_01212_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06332_ (.A1(_01377_),
    .A2(_01830_),
    .A3(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06333_ (.I(\dp.rf.rf[2][23] ),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06334_ (.I(\dp.rf.rf[3][23] ),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06335_ (.I(\dp.rf.rf[6][23] ),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06336_ (.I(\dp.rf.rf[7][23] ),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06337_ (.I0(_01834_),
    .I1(_01835_),
    .I2(_01836_),
    .I3(_01837_),
    .S0(net7),
    .S1(net537),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06338_ (.I0(\dp.rf.rf[1][23] ),
    .I1(\dp.rf.rf[5][23] ),
    .S(net537),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_366_clk (.I(clknet_6_27__leaf_clk),
    .Z(clknet_leaf_366_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06340_ (.A1(\dp.rf.rf[4][23] ),
    .A2(net520),
    .B1(_01839_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06341_ (.A1(_01140_),
    .A2(_01838_),
    .B(_01841_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06342_ (.I0(\dp.rf.rf[10][23] ),
    .I1(\dp.rf.rf[11][23] ),
    .I2(\dp.rf.rf[14][23] ),
    .I3(\dp.rf.rf[15][23] ),
    .S0(net541),
    .S1(net9),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06343_ (.I0(\dp.rf.rf[8][23] ),
    .I1(\dp.rf.rf[9][23] ),
    .I2(\dp.rf.rf[12][23] ),
    .I3(\dp.rf.rf[13][23] ),
    .S0(net541),
    .S1(net9),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06344_ (.I0(_01843_),
    .I1(_01844_),
    .S(_01140_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_365_clk (.I(clknet_6_27__leaf_clk),
    .Z(clknet_leaf_365_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06346_ (.I0(\dp.rf.rf[26][23] ),
    .I1(\dp.rf.rf[27][23] ),
    .I2(\dp.rf.rf[30][23] ),
    .I3(\dp.rf.rf[31][23] ),
    .S0(net541),
    .S1(net9),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06347_ (.I0(\dp.rf.rf[24][23] ),
    .I1(\dp.rf.rf[25][23] ),
    .I2(\dp.rf.rf[28][23] ),
    .I3(\dp.rf.rf[29][23] ),
    .S0(net541),
    .S1(net9),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06348_ (.I0(_01847_),
    .I1(_01848_),
    .S(_01140_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06349_ (.A1(net10),
    .A2(net517),
    .A3(_01849_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06350_ (.A1(_01458_),
    .A2(_01842_),
    .B1(_01845_),
    .B2(_01440_),
    .C(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06351_ (.A1(_01833_),
    .A2(_01851_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06352_ (.I(_01852_),
    .ZN(_05179_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06353_ (.A1(net15),
    .A2(_01165_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06354_ (.A1(_01320_),
    .A2(_01853_),
    .B(_01325_),
    .ZN(_05445_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06355_ (.I0(\dp.rf.rf[24][22] ),
    .I1(\dp.rf.rf[25][22] ),
    .I2(\dp.rf.rf[26][22] ),
    .I3(\dp.rf.rf[27][22] ),
    .S0(net13),
    .S1(net14),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06356_ (.I0(\dp.rf.rf[16][22] ),
    .I1(\dp.rf.rf[17][22] ),
    .I2(\dp.rf.rf[18][22] ),
    .I3(\dp.rf.rf[19][22] ),
    .S0(net13),
    .S1(net14),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06357_ (.I0(_01854_),
    .I1(_01855_),
    .S(_01066_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06358_ (.I0(\dp.rf.rf[28][22] ),
    .I1(\dp.rf.rf[29][22] ),
    .I2(\dp.rf.rf[30][22] ),
    .I3(\dp.rf.rf[31][22] ),
    .S0(net548),
    .S1(net14),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06359_ (.I0(\dp.rf.rf[20][22] ),
    .I1(\dp.rf.rf[21][22] ),
    .I2(\dp.rf.rf[22][22] ),
    .I3(\dp.rf.rf[23][22] ),
    .S0(net13),
    .S1(net14),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06360_ (.I0(_01857_),
    .I1(_01858_),
    .S(_01066_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06361_ (.I0(_01856_),
    .I1(_01859_),
    .S(net15),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06362_ (.I0(\dp.rf.rf[8][22] ),
    .I1(\dp.rf.rf[9][22] ),
    .I2(\dp.rf.rf[10][22] ),
    .I3(\dp.rf.rf[11][22] ),
    .S0(net548),
    .S1(net14),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06363_ (.I0(\dp.rf.rf[0][22] ),
    .I1(\dp.rf.rf[1][22] ),
    .I2(\dp.rf.rf[2][22] ),
    .I3(\dp.rf.rf[3][22] ),
    .S0(net548),
    .S1(net14),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06364_ (.I0(_01861_),
    .I1(_01862_),
    .S(_01066_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06365_ (.I0(\dp.rf.rf[12][22] ),
    .I1(\dp.rf.rf[13][22] ),
    .I2(\dp.rf.rf[14][22] ),
    .I3(\dp.rf.rf[15][22] ),
    .S0(net548),
    .S1(net14),
    .Z(_01864_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06366_ (.I0(\dp.rf.rf[4][22] ),
    .I1(\dp.rf.rf[5][22] ),
    .I2(\dp.rf.rf[6][22] ),
    .I3(\dp.rf.rf[7][22] ),
    .S0(net548),
    .S1(net14),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06367_ (.I0(_01864_),
    .I1(_01865_),
    .S(_01066_),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06368_ (.I0(_01863_),
    .I1(_01866_),
    .S(net15),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06369_ (.A1(net17),
    .A2(_01860_),
    .B1(_01867_),
    .B2(_01309_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06370_ (.A1(_01311_),
    .A2(_01868_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06371_ (.A1(_01311_),
    .A2(_05445_[0]),
    .B(_01869_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06372_ (.A1(net511),
    .A2(_01870_),
    .Z(_05184_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06373_ (.I(_05184_[0]),
    .ZN(_05188_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06374_ (.I0(\dp.rf.rf[26][22] ),
    .I1(\dp.rf.rf[27][22] ),
    .I2(\dp.rf.rf[30][22] ),
    .I3(\dp.rf.rf[31][22] ),
    .S0(net545),
    .S1(net535),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06375_ (.I0(\dp.rf.rf[24][22] ),
    .I1(\dp.rf.rf[25][22] ),
    .I2(\dp.rf.rf[28][22] ),
    .I3(\dp.rf.rf[29][22] ),
    .S0(net545),
    .S1(net535),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06376_ (.I0(_01871_),
    .I1(_01872_),
    .S(_01140_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06377_ (.A1(net519),
    .A2(_01873_),
    .B(net517),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06378_ (.I0(\dp.rf.rf[22][22] ),
    .I1(\dp.rf.rf[23][22] ),
    .S(net545),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06379_ (.I(_01875_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06380_ (.A1(net536),
    .A2(_01876_),
    .B(net523),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06381_ (.I(\dp.rf.rf[18][22] ),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _06382_ (.A1(_01878_),
    .A2(net533),
    .A3(net532),
    .A4(_01125_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06383_ (.I0(\dp.rf.rf[18][22] ),
    .I1(\dp.rf.rf[19][22] ),
    .S(net545),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06384_ (.I(_01880_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06385_ (.A1(net521),
    .A2(_01879_),
    .A3(_01881_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06386_ (.I0(\dp.rf.rf[17][22] ),
    .I1(\dp.rf.rf[21][22] ),
    .S(net535),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06387_ (.A1(_01148_),
    .A2(_01883_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06388_ (.A1(\dp.rf.rf[20][22] ),
    .A2(net545),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06389_ (.A1(_01884_),
    .A2(_01885_),
    .B(_01144_),
    .C(net529),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06390_ (.I(\dp.rf.rf[16][22] ),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06391_ (.A1(_01887_),
    .A2(_01385_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06392_ (.A1(_01877_),
    .A2(_01882_),
    .B1(_01886_),
    .B2(_01888_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06393_ (.I0(\dp.rf.rf[8][22] ),
    .I1(\dp.rf.rf[9][22] ),
    .I2(\dp.rf.rf[12][22] ),
    .I3(\dp.rf.rf[13][22] ),
    .S0(net545),
    .S1(net535),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06394_ (.I0(\dp.rf.rf[1][22] ),
    .I1(\dp.rf.rf[5][22] ),
    .S(net535),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06395_ (.A1(_01148_),
    .A2(_01891_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06396_ (.A1(\dp.rf.rf[4][22] ),
    .A2(net545),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06397_ (.A1(_01892_),
    .A2(_01893_),
    .B(net529),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06398_ (.I0(\dp.rf.rf[10][22] ),
    .I1(\dp.rf.rf[11][22] ),
    .I2(\dp.rf.rf[14][22] ),
    .I3(\dp.rf.rf[15][22] ),
    .S0(net545),
    .S1(net535),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06399_ (.I0(\dp.rf.rf[2][22] ),
    .I1(\dp.rf.rf[3][22] ),
    .I2(\dp.rf.rf[6][22] ),
    .I3(\dp.rf.rf[7][22] ),
    .S0(net545),
    .S1(net535),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06400_ (.I0(_01895_),
    .I1(_01896_),
    .S(_01144_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _06401_ (.A1(_01279_),
    .A2(_01890_),
    .B1(_01894_),
    .B2(_01458_),
    .C1(_01781_),
    .C2(_01897_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06402_ (.A1(_01874_),
    .A2(_01889_),
    .B(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_360_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_360_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06404_ (.I(_01899_),
    .ZN(_05187_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_358_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_358_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06406_ (.A1(net14),
    .A2(_01165_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06407_ (.A1(_01320_),
    .A2(_01901_),
    .B(_01325_),
    .ZN(_05441_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06408_ (.I0(\dp.rf.rf[24][21] ),
    .I1(\dp.rf.rf[25][21] ),
    .I2(\dp.rf.rf[26][21] ),
    .I3(\dp.rf.rf[27][21] ),
    .S0(net13),
    .S1(net14),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06409_ (.I0(\dp.rf.rf[16][21] ),
    .I1(\dp.rf.rf[17][21] ),
    .I2(\dp.rf.rf[18][21] ),
    .I3(\dp.rf.rf[19][21] ),
    .S0(net548),
    .S1(net14),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06410_ (.I0(_01902_),
    .I1(_01903_),
    .S(_01066_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06411_ (.I0(\dp.rf.rf[28][21] ),
    .I1(\dp.rf.rf[29][21] ),
    .I2(\dp.rf.rf[30][21] ),
    .I3(\dp.rf.rf[31][21] ),
    .S0(net13),
    .S1(net14),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06412_ (.I0(\dp.rf.rf[20][21] ),
    .I1(\dp.rf.rf[21][21] ),
    .I2(\dp.rf.rf[22][21] ),
    .I3(\dp.rf.rf[23][21] ),
    .S0(net548),
    .S1(net14),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06413_ (.I0(_01905_),
    .I1(_01906_),
    .S(_01066_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06414_ (.I0(_01904_),
    .I1(_01907_),
    .S(net15),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06415_ (.I0(\dp.rf.rf[8][21] ),
    .I1(\dp.rf.rf[9][21] ),
    .I2(\dp.rf.rf[10][21] ),
    .I3(\dp.rf.rf[11][21] ),
    .S0(net548),
    .S1(net14),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06416_ (.I0(\dp.rf.rf[0][21] ),
    .I1(\dp.rf.rf[1][21] ),
    .I2(\dp.rf.rf[2][21] ),
    .I3(\dp.rf.rf[3][21] ),
    .S0(net548),
    .S1(net14),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06417_ (.I0(_01909_),
    .I1(_01910_),
    .S(_01066_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06418_ (.I0(\dp.rf.rf[12][21] ),
    .I1(\dp.rf.rf[13][21] ),
    .I2(\dp.rf.rf[14][21] ),
    .I3(\dp.rf.rf[15][21] ),
    .S0(net548),
    .S1(net14),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06419_ (.I0(\dp.rf.rf[4][21] ),
    .I1(\dp.rf.rf[5][21] ),
    .I2(\dp.rf.rf[6][21] ),
    .I3(\dp.rf.rf[7][21] ),
    .S0(net548),
    .S1(net14),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06420_ (.I0(_01912_),
    .I1(_01913_),
    .S(_01066_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06421_ (.I0(_01911_),
    .I1(_01914_),
    .S(net15),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06422_ (.A1(net17),
    .A2(_01908_),
    .B1(_01915_),
    .B2(_01309_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06423_ (.A1(_01311_),
    .A2(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06424_ (.A1(_01311_),
    .A2(_05441_[0]),
    .B(_01917_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06425_ (.A1(net511),
    .A2(_01918_),
    .Z(_05192_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06426_ (.I(_05192_[0]),
    .ZN(_05196_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06427_ (.I0(\dp.rf.rf[26][21] ),
    .I1(\dp.rf.rf[27][21] ),
    .I2(\dp.rf.rf[30][21] ),
    .I3(\dp.rf.rf[31][21] ),
    .S0(net544),
    .S1(net535),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06428_ (.I0(\dp.rf.rf[24][21] ),
    .I1(\dp.rf.rf[25][21] ),
    .I2(\dp.rf.rf[28][21] ),
    .I3(\dp.rf.rf[29][21] ),
    .S0(net544),
    .S1(net535),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06429_ (.I0(_01919_),
    .I1(_01920_),
    .S(_01140_),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06430_ (.A1(net519),
    .A2(_01921_),
    .B(net517),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06431_ (.I0(\dp.rf.rf[22][21] ),
    .I1(\dp.rf.rf[23][21] ),
    .S(net545),
    .Z(_01923_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06432_ (.A1(_01167_),
    .A2(_01923_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06433_ (.A1(net523),
    .A2(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06434_ (.I(\dp.rf.rf[18][21] ),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _06435_ (.A1(_01926_),
    .A2(net533),
    .A3(net532),
    .A4(_01125_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06436_ (.I0(\dp.rf.rf[18][21] ),
    .I1(\dp.rf.rf[19][21] ),
    .S(net545),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06437_ (.I(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06438_ (.A1(net521),
    .A2(_01927_),
    .A3(_01929_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06439_ (.I0(\dp.rf.rf[17][21] ),
    .I1(\dp.rf.rf[21][21] ),
    .S(net535),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06440_ (.A1(_01148_),
    .A2(_01931_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06441_ (.A1(\dp.rf.rf[20][21] ),
    .A2(net545),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06442_ (.A1(_01932_),
    .A2(_01933_),
    .B(_01144_),
    .C(net529),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06443_ (.I(\dp.rf.rf[16][21] ),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06444_ (.A1(_01935_),
    .A2(_01385_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06445_ (.A1(_01925_),
    .A2(_01930_),
    .B1(_01934_),
    .B2(_01936_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06446_ (.I0(\dp.rf.rf[8][21] ),
    .I1(\dp.rf.rf[9][21] ),
    .I2(\dp.rf.rf[12][21] ),
    .I3(\dp.rf.rf[13][21] ),
    .S0(net544),
    .S1(net535),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06447_ (.I0(\dp.rf.rf[1][21] ),
    .I1(\dp.rf.rf[5][21] ),
    .S(net535),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06448_ (.A1(_01148_),
    .A2(_01939_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06449_ (.A1(\dp.rf.rf[4][21] ),
    .A2(net545),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06450_ (.A1(_01940_),
    .A2(_01941_),
    .B(net529),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06451_ (.I0(\dp.rf.rf[10][21] ),
    .I1(\dp.rf.rf[11][21] ),
    .I2(\dp.rf.rf[14][21] ),
    .I3(\dp.rf.rf[15][21] ),
    .S0(net544),
    .S1(net535),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06452_ (.I0(\dp.rf.rf[2][21] ),
    .I1(\dp.rf.rf[3][21] ),
    .I2(\dp.rf.rf[6][21] ),
    .I3(\dp.rf.rf[7][21] ),
    .S0(net544),
    .S1(net535),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06453_ (.I0(_01943_),
    .I1(_01944_),
    .S(_01144_),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _06454_ (.A1(_01279_),
    .A2(_01938_),
    .B1(_01942_),
    .B2(_01458_),
    .C1(_01781_),
    .C2(_01945_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06455_ (.A1(_01922_),
    .A2(_01937_),
    .B(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_351_clk (.I(clknet_6_48__leaf_clk),
    .Z(clknet_leaf_351_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06457_ (.I(_01947_),
    .ZN(_05195_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06458_ (.A1(net13),
    .A2(_01165_),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06459_ (.A1(_01320_),
    .A2(_01948_),
    .B(_01325_),
    .ZN(_05437_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06460_ (.I0(\dp.rf.rf[28][20] ),
    .I1(\dp.rf.rf[29][20] ),
    .I2(\dp.rf.rf[30][20] ),
    .I3(\dp.rf.rf[31][20] ),
    .S0(net549),
    .S1(net14),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06461_ (.I0(\dp.rf.rf[20][20] ),
    .I1(\dp.rf.rf[21][20] ),
    .I2(\dp.rf.rf[22][20] ),
    .I3(\dp.rf.rf[23][20] ),
    .S0(net13),
    .S1(net546),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06462_ (.I0(\dp.rf.rf[24][20] ),
    .I1(\dp.rf.rf[25][20] ),
    .I2(\dp.rf.rf[26][20] ),
    .I3(\dp.rf.rf[27][20] ),
    .S0(net549),
    .S1(net14),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06463_ (.I0(\dp.rf.rf[16][20] ),
    .I1(\dp.rf.rf[17][20] ),
    .I2(\dp.rf.rf[18][20] ),
    .I3(\dp.rf.rf[19][20] ),
    .S0(net13),
    .S1(net546),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06464_ (.I0(_01949_),
    .I1(_01950_),
    .I2(_01951_),
    .I3(_01952_),
    .S0(_01066_),
    .S1(_01055_),
    .Z(_01953_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06465_ (.A1(_01064_),
    .A2(_01953_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_349_clk (.I(clknet_6_48__leaf_clk),
    .Z(clknet_leaf_349_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06467_ (.I0(\dp.rf.rf[12][20] ),
    .I1(\dp.rf.rf[13][20] ),
    .I2(\dp.rf.rf[14][20] ),
    .I3(\dp.rf.rf[15][20] ),
    .S0(net13),
    .S1(net14),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06468_ (.I0(\dp.rf.rf[8][20] ),
    .I1(\dp.rf.rf[9][20] ),
    .I2(\dp.rf.rf[10][20] ),
    .I3(\dp.rf.rf[11][20] ),
    .S0(net13),
    .S1(net14),
    .Z(_01957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06469_ (.I0(_01956_),
    .I1(_01957_),
    .S(_01055_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06470_ (.A1(_01084_),
    .A2(_01958_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06471_ (.I0(\dp.rf.rf[4][20] ),
    .I1(\dp.rf.rf[5][20] ),
    .I2(\dp.rf.rf[6][20] ),
    .I3(\dp.rf.rf[7][20] ),
    .S0(net550),
    .S1(net14),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06472_ (.I0(\dp.rf.rf[0][20] ),
    .I1(\dp.rf.rf[1][20] ),
    .I2(\dp.rf.rf[2][20] ),
    .I3(\dp.rf.rf[3][20] ),
    .S0(net550),
    .S1(net14),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06473_ (.I0(_01960_),
    .I1(_01961_),
    .S(_01055_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _06474_ (.A1(_01067_),
    .A2(_01962_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06475_ (.A1(_01329_),
    .A2(_01963_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06476_ (.A1(_01954_),
    .A2(_01959_),
    .A3(_01964_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06477_ (.A1(_01311_),
    .A2(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06478_ (.A1(_01119_),
    .A2(_05437_[0]),
    .B(_01966_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06479_ (.A1(net511),
    .A2(_01967_),
    .Z(_05200_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06480_ (.I(_05200_[0]),
    .ZN(_05204_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06481_ (.I0(\dp.rf.rf[26][20] ),
    .I1(\dp.rf.rf[27][20] ),
    .I2(\dp.rf.rf[30][20] ),
    .I3(\dp.rf.rf[31][20] ),
    .S0(net7),
    .S1(net9),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06482_ (.I0(\dp.rf.rf[24][20] ),
    .I1(\dp.rf.rf[25][20] ),
    .I2(\dp.rf.rf[28][20] ),
    .I3(\dp.rf.rf[29][20] ),
    .S0(net7),
    .S1(net9),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_348_clk (.I(clknet_6_49__leaf_clk),
    .Z(clknet_leaf_348_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06484_ (.I0(_01968_),
    .I1(_01969_),
    .S(_01140_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06485_ (.A1(net519),
    .A2(_01971_),
    .B(net517),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06486_ (.I0(\dp.rf.rf[22][20] ),
    .I1(\dp.rf.rf[23][20] ),
    .S(net7),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06487_ (.I(_01973_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06488_ (.A1(net537),
    .A2(_01974_),
    .B(net523),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06489_ (.I(\dp.rf.rf[18][20] ),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06490_ (.A1(_01976_),
    .A2(_01030_),
    .A3(_01101_),
    .A4(_01125_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06491_ (.I0(\dp.rf.rf[18][20] ),
    .I1(\dp.rf.rf[19][20] ),
    .S(net7),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06492_ (.I(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06493_ (.A1(net522),
    .A2(_01977_),
    .A3(_01979_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06494_ (.I0(\dp.rf.rf[17][20] ),
    .I1(\dp.rf.rf[21][20] ),
    .S(net9),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06495_ (.A1(_01148_),
    .A2(_01981_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06496_ (.A1(\dp.rf.rf[20][20] ),
    .A2(net540),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06497_ (.A1(_01982_),
    .A2(_01983_),
    .B(_01144_),
    .C(net165),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06498_ (.I(\dp.rf.rf[16][20] ),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06499_ (.A1(_01985_),
    .A2(_01385_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06500_ (.A1(_01975_),
    .A2(_01980_),
    .B1(_01984_),
    .B2(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06501_ (.I0(\dp.rf.rf[8][20] ),
    .I1(\dp.rf.rf[9][20] ),
    .I2(\dp.rf.rf[12][20] ),
    .I3(\dp.rf.rf[13][20] ),
    .S0(net541),
    .S1(net9),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06502_ (.I0(\dp.rf.rf[1][20] ),
    .I1(\dp.rf.rf[5][20] ),
    .S(net9),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06503_ (.A1(_01148_),
    .A2(_01989_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06504_ (.A1(\dp.rf.rf[4][20] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06505_ (.A1(_01990_),
    .A2(_01991_),
    .B(net529),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06506_ (.I0(\dp.rf.rf[10][20] ),
    .I1(\dp.rf.rf[11][20] ),
    .I2(\dp.rf.rf[14][20] ),
    .I3(\dp.rf.rf[15][20] ),
    .S0(net541),
    .S1(net9),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06507_ (.I0(\dp.rf.rf[2][20] ),
    .I1(\dp.rf.rf[3][20] ),
    .I2(\dp.rf.rf[6][20] ),
    .I3(\dp.rf.rf[7][20] ),
    .S0(net541),
    .S1(net9),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06508_ (.I0(_01993_),
    .I1(_01994_),
    .S(_01144_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _06509_ (.A1(_01279_),
    .A2(_01988_),
    .B1(_01992_),
    .B2(_01458_),
    .C1(_01781_),
    .C2(_01995_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06510_ (.A1(_01972_),
    .A2(_01987_),
    .B(_01996_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_334_clk (.I(clknet_6_54__leaf_clk),
    .Z(clknet_leaf_334_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06512_ (.I(_01997_),
    .ZN(_05203_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_333_clk (.I(clknet_6_54__leaf_clk),
    .Z(clknet_leaf_333_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06514_ (.A1(net25),
    .A2(_01315_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06515_ (.A1(_01212_),
    .A2(_01123_),
    .B1(net528),
    .B2(_01144_),
    .C(_01999_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06516_ (.A1(net11),
    .A2(_01165_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06517_ (.A1(_01320_),
    .A2(_02001_),
    .B(_01325_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06518_ (.A1(_01098_),
    .A2(_01107_),
    .A3(_01115_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06519_ (.A1(_02003_),
    .A2(_01134_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06520_ (.I0(_02000_),
    .I1(_02002_),
    .S(_02004_),
    .Z(_05433_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06521_ (.I0(\dp.rf.rf[24][19] ),
    .I1(\dp.rf.rf[25][19] ),
    .I2(\dp.rf.rf[26][19] ),
    .I3(\dp.rf.rf[27][19] ),
    .S0(net547),
    .S1(net546),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06522_ (.I0(\dp.rf.rf[16][19] ),
    .I1(\dp.rf.rf[17][19] ),
    .I2(\dp.rf.rf[18][19] ),
    .I3(\dp.rf.rf[19][19] ),
    .S0(net547),
    .S1(net546),
    .Z(_02006_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06523_ (.I0(\dp.rf.rf[28][19] ),
    .I1(\dp.rf.rf[29][19] ),
    .I2(\dp.rf.rf[30][19] ),
    .I3(\dp.rf.rf[31][19] ),
    .S0(net547),
    .S1(net546),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06524_ (.I0(\dp.rf.rf[20][19] ),
    .I1(\dp.rf.rf[21][19] ),
    .I2(\dp.rf.rf[22][19] ),
    .I3(\dp.rf.rf[23][19] ),
    .S0(net547),
    .S1(net546),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06525_ (.I0(_02005_),
    .I1(_02006_),
    .I2(_02007_),
    .I3(_02008_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06526_ (.I0(\dp.rf.rf[8][19] ),
    .I1(\dp.rf.rf[9][19] ),
    .I2(\dp.rf.rf[10][19] ),
    .I3(\dp.rf.rf[11][19] ),
    .S0(net547),
    .S1(net546),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06527_ (.I0(\dp.rf.rf[0][19] ),
    .I1(\dp.rf.rf[1][19] ),
    .I2(\dp.rf.rf[2][19] ),
    .I3(\dp.rf.rf[3][19] ),
    .S0(net547),
    .S1(net546),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06528_ (.I0(\dp.rf.rf[12][19] ),
    .I1(\dp.rf.rf[13][19] ),
    .I2(\dp.rf.rf[14][19] ),
    .I3(\dp.rf.rf[15][19] ),
    .S0(net547),
    .S1(net546),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06529_ (.I0(\dp.rf.rf[4][19] ),
    .I1(\dp.rf.rf[5][19] ),
    .I2(\dp.rf.rf[6][19] ),
    .I3(\dp.rf.rf[7][19] ),
    .S0(net547),
    .S1(net546),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06530_ (.I0(_02010_),
    .I1(_02011_),
    .I2(_02012_),
    .I3(_02013_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06531_ (.A1(net17),
    .A2(_02009_),
    .B1(_02014_),
    .B2(_01309_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06532_ (.A1(_01311_),
    .A2(_02015_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06533_ (.A1(_01311_),
    .A2(_05433_[0]),
    .B(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06534_ (.A1(_01110_),
    .A2(_02017_),
    .Z(_05208_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06535_ (.I(_05208_[0]),
    .ZN(_05212_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06536_ (.I0(\dp.rf.rf[10][19] ),
    .I1(\dp.rf.rf[11][19] ),
    .I2(\dp.rf.rf[14][19] ),
    .I3(\dp.rf.rf[15][19] ),
    .S0(net539),
    .S1(net534),
    .Z(_02018_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06537_ (.I0(\dp.rf.rf[8][19] ),
    .I1(\dp.rf.rf[9][19] ),
    .I2(\dp.rf.rf[12][19] ),
    .I3(\dp.rf.rf[13][19] ),
    .S0(net539),
    .S1(net534),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06538_ (.I0(_02018_),
    .I1(_02019_),
    .S(_01140_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06539_ (.A1(_01440_),
    .A2(_02020_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06540_ (.I0(\dp.rf.rf[2][19] ),
    .I1(\dp.rf.rf[3][19] ),
    .I2(\dp.rf.rf[6][19] ),
    .I3(\dp.rf.rf[7][19] ),
    .S0(net539),
    .S1(net534),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06541_ (.A1(_01535_),
    .A2(_02022_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_330_clk (.I(clknet_6_54__leaf_clk),
    .Z(clknet_leaf_330_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06543_ (.I0(\dp.rf.rf[1][19] ),
    .I1(\dp.rf.rf[5][19] ),
    .S(net534),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06544_ (.A1(\dp.rf.rf[4][19] ),
    .A2(_01245_),
    .B1(_02025_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06545_ (.A1(net526),
    .A2(_02026_),
    .B(_01242_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _06546_ (.A1(_02021_),
    .A2(_02023_),
    .A3(_02027_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06547_ (.I0(\dp.rf.rf[22][19] ),
    .I1(\dp.rf.rf[23][19] ),
    .S(net538),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06548_ (.A1(\dp.rf.rf[18][19] ),
    .A2(_01368_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06549_ (.A1(\dp.rf.rf[19][19] ),
    .A2(net538),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06550_ (.A1(net522),
    .A2(_02031_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06551_ (.A1(_01167_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_02032_),
    .C(_01284_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06552_ (.I(\dp.rf.rf[20][19] ),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06553_ (.I0(\dp.rf.rf[17][19] ),
    .I1(\dp.rf.rf[21][19] ),
    .S(net534),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06554_ (.A1(_01148_),
    .A2(_02035_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06555_ (.A1(_02034_),
    .A2(_01451_),
    .B(_02036_),
    .C(net8),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06556_ (.A1(\dp.rf.rf[16][19] ),
    .A2(_01467_),
    .B1(_02037_),
    .B2(net524),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06557_ (.I0(\dp.rf.rf[26][19] ),
    .I1(\dp.rf.rf[27][19] ),
    .I2(\dp.rf.rf[30][19] ),
    .I3(\dp.rf.rf[31][19] ),
    .S0(net539),
    .S1(net534),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06558_ (.I0(\dp.rf.rf[24][19] ),
    .I1(\dp.rf.rf[25][19] ),
    .I2(\dp.rf.rf[28][19] ),
    .I3(\dp.rf.rf[29][19] ),
    .S0(net539),
    .S1(net534),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06559_ (.I0(_02039_),
    .I1(_02040_),
    .S(_01140_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06560_ (.A1(_01144_),
    .A2(_02041_),
    .B(_01216_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06561_ (.A1(_02033_),
    .A2(_02038_),
    .B(_02042_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06562_ (.A1(_02028_),
    .A2(_02043_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _06563_ (.I(_02044_),
    .ZN(_05211_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06564_ (.A1(_01144_),
    .A2(_01123_),
    .B1(net528),
    .B2(_01167_),
    .C(_01999_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_328_clk (.I(clknet_6_51__leaf_clk),
    .Z(clknet_leaf_328_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06566_ (.I0(_02000_),
    .I1(_02045_),
    .S(_01135_),
    .Z(_05429_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_326_clk (.I(clknet_6_51__leaf_clk),
    .Z(clknet_leaf_326_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_324_clk (.I(clknet_6_51__leaf_clk),
    .Z(clknet_leaf_324_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06569_ (.I0(\dp.rf.rf[24][18] ),
    .I1(\dp.rf.rf[25][18] ),
    .I2(\dp.rf.rf[26][18] ),
    .I3(\dp.rf.rf[27][18] ),
    .S0(net547),
    .S1(net546),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06570_ (.I0(\dp.rf.rf[16][18] ),
    .I1(\dp.rf.rf[17][18] ),
    .I2(\dp.rf.rf[18][18] ),
    .I3(\dp.rf.rf[19][18] ),
    .S0(net547),
    .S1(net546),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_319_clk (.I(clknet_6_56__leaf_clk),
    .Z(clknet_leaf_319_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06572_ (.I0(\dp.rf.rf[28][18] ),
    .I1(\dp.rf.rf[29][18] ),
    .I2(\dp.rf.rf[30][18] ),
    .I3(\dp.rf.rf[31][18] ),
    .S0(net547),
    .S1(net546),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06573_ (.I0(\dp.rf.rf[20][18] ),
    .I1(\dp.rf.rf[21][18] ),
    .I2(\dp.rf.rf[22][18] ),
    .I3(\dp.rf.rf[23][18] ),
    .S0(net547),
    .S1(net546),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06574_ (.I0(_02049_),
    .I1(_02050_),
    .I2(_02052_),
    .I3(_02053_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06575_ (.I0(\dp.rf.rf[8][18] ),
    .I1(\dp.rf.rf[9][18] ),
    .I2(\dp.rf.rf[10][18] ),
    .I3(\dp.rf.rf[11][18] ),
    .S0(net547),
    .S1(net546),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06576_ (.I0(\dp.rf.rf[0][18] ),
    .I1(\dp.rf.rf[1][18] ),
    .I2(\dp.rf.rf[2][18] ),
    .I3(\dp.rf.rf[3][18] ),
    .S0(net547),
    .S1(net546),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06577_ (.I0(\dp.rf.rf[12][18] ),
    .I1(\dp.rf.rf[13][18] ),
    .I2(\dp.rf.rf[14][18] ),
    .I3(\dp.rf.rf[15][18] ),
    .S0(net547),
    .S1(net546),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06578_ (.I0(\dp.rf.rf[4][18] ),
    .I1(\dp.rf.rf[5][18] ),
    .I2(\dp.rf.rf[6][18] ),
    .I3(\dp.rf.rf[7][18] ),
    .S0(net547),
    .S1(net546),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06579_ (.I0(_02055_),
    .I1(_02056_),
    .I2(_02057_),
    .I3(_02058_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06580_ (.A1(net17),
    .A2(_02054_),
    .B1(_02059_),
    .B2(_01309_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06581_ (.A1(_01311_),
    .A2(_02060_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06582_ (.A1(_01311_),
    .A2(_05429_[0]),
    .B(_02061_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06583_ (.A1(_01110_),
    .A2(_02062_),
    .Z(_05216_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06584_ (.I(_05216_[0]),
    .ZN(_05220_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06585_ (.I0(\dp.rf.rf[10][18] ),
    .I1(\dp.rf.rf[11][18] ),
    .I2(\dp.rf.rf[14][18] ),
    .I3(\dp.rf.rf[15][18] ),
    .S0(net539),
    .S1(net534),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06586_ (.I0(\dp.rf.rf[8][18] ),
    .I1(\dp.rf.rf[9][18] ),
    .I2(\dp.rf.rf[12][18] ),
    .I3(\dp.rf.rf[13][18] ),
    .S0(net539),
    .S1(net534),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06587_ (.I0(_02063_),
    .I1(_02064_),
    .S(_01140_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06588_ (.A1(_01440_),
    .A2(_02065_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06589_ (.I0(\dp.rf.rf[2][18] ),
    .I1(\dp.rf.rf[3][18] ),
    .I2(\dp.rf.rf[6][18] ),
    .I3(\dp.rf.rf[7][18] ),
    .S0(net539),
    .S1(net534),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06590_ (.A1(_01535_),
    .A2(_02067_),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06591_ (.I0(\dp.rf.rf[1][18] ),
    .I1(\dp.rf.rf[5][18] ),
    .S(net534),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06592_ (.A1(\dp.rf.rf[4][18] ),
    .A2(_01245_),
    .B1(_02069_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _06593_ (.A1(net526),
    .A2(_02070_),
    .B(_01242_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _06594_ (.A1(_02066_),
    .A2(_02068_),
    .A3(_02071_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06595_ (.I0(\dp.rf.rf[26][18] ),
    .I1(\dp.rf.rf[27][18] ),
    .I2(\dp.rf.rf[30][18] ),
    .I3(\dp.rf.rf[31][18] ),
    .S0(net539),
    .S1(net534),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06596_ (.I0(\dp.rf.rf[24][18] ),
    .I1(\dp.rf.rf[25][18] ),
    .I2(\dp.rf.rf[28][18] ),
    .I3(\dp.rf.rf[29][18] ),
    .S0(net539),
    .S1(net534),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06597_ (.I0(_02073_),
    .I1(_02074_),
    .S(_01140_),
    .Z(_02075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06598_ (.I0(\dp.rf.rf[22][18] ),
    .I1(\dp.rf.rf[23][18] ),
    .S(net538),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06599_ (.A1(_01167_),
    .A2(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06600_ (.A1(\dp.rf.rf[19][18] ),
    .A2(net538),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06601_ (.A1(net534),
    .A2(net526),
    .B1(_01368_),
    .B2(\dp.rf.rf[18][18] ),
    .C(_02078_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06602_ (.A1(net523),
    .A2(_02077_),
    .A3(_02079_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06603_ (.I(\dp.rf.rf[16][18] ),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06604_ (.I0(\dp.rf.rf[17][18] ),
    .I1(\dp.rf.rf[21][18] ),
    .S(net534),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06605_ (.A1(\dp.rf.rf[20][18] ),
    .A2(_01245_),
    .B1(_02082_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06606_ (.A1(_02081_),
    .A2(net518),
    .B1(_02083_),
    .B2(_01377_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06607_ (.A1(_01273_),
    .A2(_02075_),
    .B1(_02080_),
    .B2(_02084_),
    .C(_01216_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06608_ (.A1(_02072_),
    .A2(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _06609_ (.I(_02086_),
    .ZN(_05219_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06610_ (.A1(_01167_),
    .A2(_01123_),
    .B1(net528),
    .B2(_01140_),
    .C(_01999_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06611_ (.I0(_02045_),
    .I1(_02087_),
    .S(_01135_),
    .Z(_05425_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06612_ (.I0(\dp.rf.rf[6][17] ),
    .I1(\dp.rf.rf[7][17] ),
    .I2(\dp.rf.rf[14][17] ),
    .I3(\dp.rf.rf[15][17] ),
    .S0(net13),
    .S1(net16),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06613_ (.I0(\dp.rf.rf[2][17] ),
    .I1(\dp.rf.rf[3][17] ),
    .I2(\dp.rf.rf[10][17] ),
    .I3(\dp.rf.rf[11][17] ),
    .S0(net13),
    .S1(net16),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06614_ (.I0(_02088_),
    .I1(_02089_),
    .S(_01055_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06615_ (.A1(_01064_),
    .A2(net546),
    .A3(_02090_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06616_ (.A1(net17),
    .A2(net15),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06617_ (.I0(\dp.rf.rf[28][17] ),
    .I1(\dp.rf.rf[29][17] ),
    .I2(\dp.rf.rf[30][17] ),
    .I3(\dp.rf.rf[31][17] ),
    .S0(net13),
    .S1(net546),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06618_ (.I0(\dp.rf.rf[20][17] ),
    .I1(\dp.rf.rf[21][17] ),
    .I2(\dp.rf.rf[22][17] ),
    .I3(\dp.rf.rf[23][17] ),
    .S0(net13),
    .S1(net546),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06619_ (.I0(_02093_),
    .I1(_02094_),
    .S(_01066_),
    .Z(_02095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06620_ (.A1(_02092_),
    .A2(_02095_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06621_ (.I0(\dp.rf.rf[1][17] ),
    .I1(\dp.rf.rf[5][17] ),
    .I2(\dp.rf.rf[9][17] ),
    .I3(\dp.rf.rf[13][17] ),
    .S0(net15),
    .S1(net16),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06622_ (.I0(\dp.rf.rf[0][17] ),
    .I1(\dp.rf.rf[4][17] ),
    .I2(\dp.rf.rf[8][17] ),
    .I3(\dp.rf.rf[12][17] ),
    .S0(net15),
    .S1(net16),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06623_ (.I0(_02097_),
    .I1(_02098_),
    .S(_01045_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06624_ (.A1(_01036_),
    .A2(_01309_),
    .A3(_02099_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06625_ (.I0(\dp.rf.rf[24][17] ),
    .I1(\dp.rf.rf[25][17] ),
    .S(net547),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06626_ (.A1(net546),
    .A2(_01066_),
    .A3(_02101_),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06627_ (.I0(\dp.rf.rf[18][17] ),
    .I1(\dp.rf.rf[19][17] ),
    .S(net13),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06628_ (.A1(_01036_),
    .A2(net16),
    .A3(_02103_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06629_ (.A1(net17),
    .A2(_01055_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06630_ (.A1(net14),
    .A2(net16),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06631_ (.I0(\dp.rf.rf[26][17] ),
    .I1(\dp.rf.rf[27][17] ),
    .S(net547),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06632_ (.I0(\dp.rf.rf[16][17] ),
    .I1(\dp.rf.rf[17][17] ),
    .S(net13),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06633_ (.A1(net546),
    .A2(net16),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06634_ (.A1(_02106_),
    .A2(_02107_),
    .B1(_02108_),
    .B2(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06635_ (.A1(_02102_),
    .A2(_02104_),
    .A3(_02105_),
    .A4(_02110_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _06636_ (.A1(_02091_),
    .A2(_02096_),
    .A3(_02100_),
    .A4(_02111_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06637_ (.A1(_01311_),
    .A2(_02112_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06638_ (.A1(_01311_),
    .A2(_05425_[0]),
    .B(_02113_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06639_ (.A1(_01110_),
    .A2(_02114_),
    .Z(_05224_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06640_ (.I(_05224_[0]),
    .ZN(_05228_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06641_ (.A1(_01140_),
    .A2(net165),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06642_ (.I0(\dp.rf.rf[8][17] ),
    .I1(\dp.rf.rf[9][17] ),
    .I2(\dp.rf.rf[12][17] ),
    .I3(\dp.rf.rf[13][17] ),
    .S0(net540),
    .S1(net9),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06643_ (.I(\dp.rf.rf[4][17] ),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06644_ (.I0(\dp.rf.rf[1][17] ),
    .I1(\dp.rf.rf[5][17] ),
    .S(net9),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06645_ (.A1(net531),
    .A2(_02118_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06646_ (.A1(_02117_),
    .A2(_01451_),
    .B(_02119_),
    .C(net11),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06647_ (.A1(_01278_),
    .A2(_02116_),
    .B1(_02120_),
    .B2(_01198_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06648_ (.I0(\dp.rf.rf[18][17] ),
    .I1(\dp.rf.rf[19][17] ),
    .I2(\dp.rf.rf[22][17] ),
    .I3(\dp.rf.rf[23][17] ),
    .S0(net542),
    .S1(net9),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06649_ (.I0(\dp.rf.rf[17][17] ),
    .I1(\dp.rf.rf[21][17] ),
    .S(net9),
    .Z(_02123_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06650_ (.A1(net531),
    .A2(_02123_),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06651_ (.A1(\dp.rf.rf[20][17] ),
    .A2(net542),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06652_ (.A1(_02124_),
    .A2(_02125_),
    .B(_01144_),
    .C(net166),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06653_ (.I(\dp.rf.rf[16][17] ),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06654_ (.A1(_02127_),
    .A2(net518),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06655_ (.A1(_01284_),
    .A2(_02122_),
    .B1(_02126_),
    .B2(_02128_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06656_ (.I0(\dp.rf.rf[26][17] ),
    .I1(\dp.rf.rf[27][17] ),
    .I2(\dp.rf.rf[30][17] ),
    .I3(\dp.rf.rf[31][17] ),
    .S0(net540),
    .S1(net9),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06657_ (.A1(net8),
    .A2(_02130_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06658_ (.I0(\dp.rf.rf[24][17] ),
    .I1(\dp.rf.rf[28][17] ),
    .S(net9),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06659_ (.A1(_01208_),
    .A2(_02132_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06660_ (.I0(\dp.rf.rf[25][17] ),
    .I1(\dp.rf.rf[29][17] ),
    .S(net9),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06661_ (.A1(net540),
    .A2(_01140_),
    .A3(_02134_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _06662_ (.A1(net519),
    .A2(_02131_),
    .A3(_02133_),
    .A4(_02135_),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06663_ (.A1(_01216_),
    .A2(_02136_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06664_ (.I0(\dp.rf.rf[3][17] ),
    .I1(\dp.rf.rf[7][17] ),
    .I2(\dp.rf.rf[11][17] ),
    .I3(\dp.rf.rf[15][17] ),
    .S0(net9),
    .S1(net10),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06665_ (.I0(\dp.rf.rf[2][17] ),
    .I1(\dp.rf.rf[6][17] ),
    .I2(\dp.rf.rf[10][17] ),
    .I3(\dp.rf.rf[14][17] ),
    .S0(net9),
    .S1(net10),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06666_ (.I0(_02138_),
    .I1(_02139_),
    .S(net531),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06667_ (.A1(_01781_),
    .A2(_02140_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _06668_ (.A1(_02115_),
    .A2(_02121_),
    .B1(_02129_),
    .B2(_02137_),
    .C(_02141_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_317_clk (.I(clknet_6_56__leaf_clk),
    .Z(clknet_leaf_317_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06670_ (.I(_02142_),
    .ZN(_05227_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06671_ (.A1(_01140_),
    .A2(_01123_),
    .B1(net528),
    .B2(net531),
    .C(_01999_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06672_ (.I0(_02087_),
    .I1(_02143_),
    .S(_01135_),
    .Z(_05421_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06673_ (.I0(\dp.rf.rf[6][16] ),
    .I1(\dp.rf.rf[7][16] ),
    .I2(\dp.rf.rf[14][16] ),
    .I3(\dp.rf.rf[15][16] ),
    .S0(net549),
    .S1(net16),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06674_ (.I0(\dp.rf.rf[2][16] ),
    .I1(\dp.rf.rf[3][16] ),
    .I2(\dp.rf.rf[10][16] ),
    .I3(\dp.rf.rf[11][16] ),
    .S0(net549),
    .S1(net16),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06675_ (.I0(_02144_),
    .I1(_02145_),
    .S(_01055_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06676_ (.A1(_01064_),
    .A2(net14),
    .A3(_02146_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06677_ (.I0(\dp.rf.rf[28][16] ),
    .I1(\dp.rf.rf[29][16] ),
    .I2(\dp.rf.rf[30][16] ),
    .I3(\dp.rf.rf[31][16] ),
    .S0(net13),
    .S1(net14),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06678_ (.I0(\dp.rf.rf[20][16] ),
    .I1(\dp.rf.rf[21][16] ),
    .I2(\dp.rf.rf[22][16] ),
    .I3(\dp.rf.rf[23][16] ),
    .S0(net13),
    .S1(net546),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06679_ (.I0(_02148_),
    .I1(_02149_),
    .S(_01066_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06680_ (.A1(_02092_),
    .A2(_02150_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06681_ (.I0(\dp.rf.rf[1][16] ),
    .I1(\dp.rf.rf[5][16] ),
    .I2(\dp.rf.rf[9][16] ),
    .I3(\dp.rf.rf[13][16] ),
    .S0(net15),
    .S1(net16),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06682_ (.I0(\dp.rf.rf[0][16] ),
    .I1(\dp.rf.rf[4][16] ),
    .I2(\dp.rf.rf[8][16] ),
    .I3(\dp.rf.rf[12][16] ),
    .S0(net15),
    .S1(net16),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06683_ (.I0(_02152_),
    .I1(_02153_),
    .S(_01045_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06684_ (.A1(_01036_),
    .A2(_01309_),
    .A3(_02154_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06685_ (.I0(\dp.rf.rf[24][16] ),
    .I1(\dp.rf.rf[25][16] ),
    .S(net13),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06686_ (.A1(net14),
    .A2(_01066_),
    .A3(_02156_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06687_ (.I0(\dp.rf.rf[18][16] ),
    .I1(\dp.rf.rf[19][16] ),
    .S(net13),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06688_ (.A1(_01036_),
    .A2(net16),
    .A3(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06689_ (.I0(\dp.rf.rf[26][16] ),
    .I1(\dp.rf.rf[27][16] ),
    .S(net13),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06690_ (.I0(\dp.rf.rf[16][16] ),
    .I1(\dp.rf.rf[17][16] ),
    .S(net13),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06691_ (.A1(_02106_),
    .A2(_02160_),
    .B1(_02161_),
    .B2(_02109_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06692_ (.A1(_02105_),
    .A2(_02157_),
    .A3(_02159_),
    .A4(_02162_),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _06693_ (.A1(_02147_),
    .A2(_02151_),
    .A3(_02155_),
    .A4(_02163_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06694_ (.A1(_01311_),
    .A2(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06695_ (.A1(_01311_),
    .A2(_05421_[0]),
    .B(_02165_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06696_ (.A1(_01110_),
    .A2(_02166_),
    .Z(_05232_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06697_ (.I(_05232_[0]),
    .ZN(_05236_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06698_ (.I0(\dp.rf.rf[18][16] ),
    .I1(\dp.rf.rf[19][16] ),
    .I2(\dp.rf.rf[22][16] ),
    .I3(\dp.rf.rf[23][16] ),
    .S0(net7),
    .S1(net9),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06699_ (.I0(\dp.rf.rf[17][16] ),
    .I1(\dp.rf.rf[21][16] ),
    .S(net9),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06700_ (.A1(net531),
    .A2(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06701_ (.A1(\dp.rf.rf[20][16] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06702_ (.A1(_02169_),
    .A2(_02170_),
    .B(_01144_),
    .C(net165),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06703_ (.I(\dp.rf.rf[16][16] ),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06704_ (.A1(_02172_),
    .A2(net518),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06705_ (.A1(_01284_),
    .A2(_02167_),
    .B1(_02171_),
    .B2(_02173_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06706_ (.I0(\dp.rf.rf[26][16] ),
    .I1(\dp.rf.rf[27][16] ),
    .I2(\dp.rf.rf[30][16] ),
    .I3(\dp.rf.rf[31][16] ),
    .S0(net540),
    .S1(net9),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06707_ (.A1(net8),
    .A2(_02175_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06708_ (.I0(\dp.rf.rf[25][16] ),
    .I1(\dp.rf.rf[29][16] ),
    .S(net9),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06709_ (.I0(\dp.rf.rf[24][16] ),
    .I1(\dp.rf.rf[28][16] ),
    .S(net9),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06710_ (.A1(_01585_),
    .A2(_02177_),
    .B1(_02178_),
    .B2(_01208_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06711_ (.A1(_01580_),
    .A2(_02176_),
    .A3(_02179_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06712_ (.I0(\dp.rf.rf[10][16] ),
    .I1(\dp.rf.rf[11][16] ),
    .I2(\dp.rf.rf[14][16] ),
    .I3(\dp.rf.rf[15][16] ),
    .S0(net7),
    .S1(net9),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06713_ (.I0(\dp.rf.rf[8][16] ),
    .I1(\dp.rf.rf[9][16] ),
    .I2(\dp.rf.rf[12][16] ),
    .I3(\dp.rf.rf[13][16] ),
    .S0(net7),
    .S1(net9),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06714_ (.I0(_02181_),
    .I1(_02182_),
    .S(_01140_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _06715_ (.A1(_01140_),
    .A2(_01197_),
    .A3(_01231_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06716_ (.A1(\dp.rf.rf[4][16] ),
    .A2(net541),
    .A3(_01167_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06717_ (.I0(\dp.rf.rf[1][16] ),
    .I1(\dp.rf.rf[5][16] ),
    .S(net9),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06718_ (.A1(_01148_),
    .A2(_02186_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06719_ (.I0(\dp.rf.rf[2][16] ),
    .I1(\dp.rf.rf[3][16] ),
    .I2(\dp.rf.rf[6][16] ),
    .I3(\dp.rf.rf[7][16] ),
    .S0(net7),
    .S1(net9),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06720_ (.I(_02188_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06721_ (.A1(_02184_),
    .A2(_02185_),
    .A3(_02187_),
    .B1(_02189_),
    .B2(_01232_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06722_ (.A1(_01440_),
    .A2(_02183_),
    .B1(_02190_),
    .B2(net165),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _06723_ (.A1(net515),
    .A2(_02174_),
    .A3(_02180_),
    .B(_02191_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06724_ (.I(net508),
    .ZN(_05235_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_316_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_316_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06726_ (.A1(net531),
    .A2(_01123_),
    .B1(net528),
    .B2(_01100_),
    .C(_01999_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06727_ (.I0(_02143_),
    .I1(_02194_),
    .S(_01135_),
    .Z(_05417_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06728_ (.I0(\dp.rf.rf[24][15] ),
    .I1(\dp.rf.rf[25][15] ),
    .I2(\dp.rf.rf[26][15] ),
    .I3(\dp.rf.rf[27][15] ),
    .S0(net547),
    .S1(net546),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06729_ (.I0(\dp.rf.rf[16][15] ),
    .I1(\dp.rf.rf[17][15] ),
    .I2(\dp.rf.rf[18][15] ),
    .I3(\dp.rf.rf[19][15] ),
    .S0(net547),
    .S1(net546),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_315_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_315_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06731_ (.I0(\dp.rf.rf[28][15] ),
    .I1(\dp.rf.rf[29][15] ),
    .I2(\dp.rf.rf[30][15] ),
    .I3(\dp.rf.rf[31][15] ),
    .S0(net547),
    .S1(net546),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06732_ (.I0(\dp.rf.rf[20][15] ),
    .I1(\dp.rf.rf[21][15] ),
    .I2(\dp.rf.rf[22][15] ),
    .I3(\dp.rf.rf[23][15] ),
    .S0(net547),
    .S1(net546),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06733_ (.I0(_02195_),
    .I1(_02196_),
    .I2(_02198_),
    .I3(_02199_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_313_clk (.I(clknet_6_55__leaf_clk),
    .Z(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06735_ (.I0(\dp.rf.rf[8][15] ),
    .I1(\dp.rf.rf[9][15] ),
    .I2(\dp.rf.rf[10][15] ),
    .I3(\dp.rf.rf[11][15] ),
    .S0(net547),
    .S1(net546),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06736_ (.I0(\dp.rf.rf[0][15] ),
    .I1(\dp.rf.rf[1][15] ),
    .I2(\dp.rf.rf[2][15] ),
    .I3(\dp.rf.rf[3][15] ),
    .S0(net547),
    .S1(net546),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06737_ (.I0(\dp.rf.rf[12][15] ),
    .I1(\dp.rf.rf[13][15] ),
    .I2(\dp.rf.rf[14][15] ),
    .I3(\dp.rf.rf[15][15] ),
    .S0(net547),
    .S1(net546),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06738_ (.I0(\dp.rf.rf[4][15] ),
    .I1(\dp.rf.rf[5][15] ),
    .I2(\dp.rf.rf[6][15] ),
    .I3(\dp.rf.rf[7][15] ),
    .S0(net547),
    .S1(net546),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _06739_ (.I0(_02202_),
    .I1(_02203_),
    .I2(_02204_),
    .I3(_02205_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06740_ (.A1(net17),
    .A2(_02200_),
    .B1(_02206_),
    .B2(_01309_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06741_ (.A1(_01311_),
    .A2(_02207_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06742_ (.A1(_01311_),
    .A2(_05417_[0]),
    .B(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06743_ (.A1(_01110_),
    .A2(_02209_),
    .Z(_05240_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06744_ (.I(_05240_[0]),
    .ZN(_05244_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06745_ (.I0(\dp.rf.rf[1][15] ),
    .I1(\dp.rf.rf[5][15] ),
    .S(net9),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06746_ (.A1(\dp.rf.rf[4][15] ),
    .A2(_01245_),
    .B1(_02210_),
    .B2(_01148_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06747_ (.I0(\dp.rf.rf[10][15] ),
    .I1(\dp.rf.rf[11][15] ),
    .I2(\dp.rf.rf[14][15] ),
    .I3(\dp.rf.rf[15][15] ),
    .S0(net7),
    .S1(net9),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06748_ (.I0(\dp.rf.rf[8][15] ),
    .I1(\dp.rf.rf[9][15] ),
    .I2(\dp.rf.rf[12][15] ),
    .I3(\dp.rf.rf[13][15] ),
    .S0(net7),
    .S1(net9),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06749_ (.I0(_02212_),
    .I1(_02213_),
    .S(_01140_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06750_ (.A1(_01278_),
    .A2(_02214_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06751_ (.I0(\dp.rf.rf[2][15] ),
    .I1(\dp.rf.rf[3][15] ),
    .I2(\dp.rf.rf[6][15] ),
    .I3(\dp.rf.rf[7][15] ),
    .S0(net7),
    .S1(net9),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06752_ (.A1(_01534_),
    .A2(_02216_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06753_ (.A1(_02184_),
    .A2(_02211_),
    .B(_02215_),
    .C(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06754_ (.A1(net525),
    .A2(_02218_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06755_ (.I0(\dp.rf.rf[22][15] ),
    .I1(\dp.rf.rf[23][15] ),
    .S(net542),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06756_ (.A1(\dp.rf.rf[18][15] ),
    .A2(_01368_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06757_ (.A1(\dp.rf.rf[19][15] ),
    .A2(net542),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06758_ (.A1(net522),
    .A2(_02222_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06759_ (.A1(_01167_),
    .A2(_02220_),
    .B1(_02221_),
    .B2(_02223_),
    .C(_01284_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06760_ (.I(\dp.rf.rf[20][15] ),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06761_ (.I0(\dp.rf.rf[17][15] ),
    .I1(\dp.rf.rf[21][15] ),
    .S(net534),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06762_ (.A1(_01148_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06763_ (.A1(_02225_),
    .A2(_01451_),
    .B(_02227_),
    .C(net8),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06764_ (.A1(\dp.rf.rf[16][15] ),
    .A2(_01467_),
    .B1(_02228_),
    .B2(_01177_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06765_ (.I0(\dp.rf.rf[26][15] ),
    .I1(\dp.rf.rf[27][15] ),
    .I2(\dp.rf.rf[30][15] ),
    .I3(\dp.rf.rf[31][15] ),
    .S0(net7),
    .S1(net9),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06766_ (.A1(net8),
    .A2(_02230_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06767_ (.I0(\dp.rf.rf[24][15] ),
    .I1(\dp.rf.rf[28][15] ),
    .S(net9),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06768_ (.I0(\dp.rf.rf[25][15] ),
    .I1(\dp.rf.rf[29][15] ),
    .S(net9),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06769_ (.A1(_01208_),
    .A2(_02232_),
    .B1(_02233_),
    .B2(_01585_),
    .C(_01273_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06770_ (.A1(_02224_),
    .A2(_02229_),
    .B1(_02231_),
    .B2(_02234_),
    .C(net514),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06771_ (.A1(_02219_),
    .A2(_02235_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _06772_ (.I(_02236_),
    .ZN(_05243_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06773_ (.A1(_01100_),
    .A2(_01123_),
    .B1(net528),
    .B2(_01089_),
    .C(_01999_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06774_ (.I0(_02194_),
    .I1(_02237_),
    .S(_01135_),
    .Z(_05413_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06775_ (.I0(\dp.rf.rf[24][14] ),
    .I1(\dp.rf.rf[25][14] ),
    .I2(\dp.rf.rf[26][14] ),
    .I3(\dp.rf.rf[27][14] ),
    .S0(net547),
    .S1(net546),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06776_ (.I0(\dp.rf.rf[16][14] ),
    .I1(\dp.rf.rf[17][14] ),
    .I2(\dp.rf.rf[18][14] ),
    .I3(\dp.rf.rf[19][14] ),
    .S0(net547),
    .S1(net546),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06777_ (.I0(_02238_),
    .I1(_02239_),
    .S(_01066_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06778_ (.A1(net15),
    .A2(_02240_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06779_ (.I0(\dp.rf.rf[28][14] ),
    .I1(\dp.rf.rf[29][14] ),
    .I2(\dp.rf.rf[30][14] ),
    .I3(\dp.rf.rf[31][14] ),
    .S0(net547),
    .S1(net546),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06780_ (.I0(\dp.rf.rf[20][14] ),
    .I1(\dp.rf.rf[21][14] ),
    .I2(\dp.rf.rf[22][14] ),
    .I3(\dp.rf.rf[23][14] ),
    .S0(net547),
    .S1(net546),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06781_ (.I0(_02242_),
    .I1(_02243_),
    .S(_01066_),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06782_ (.A1(_01055_),
    .A2(_02244_),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06783_ (.I0(\dp.rf.rf[12][14] ),
    .I1(\dp.rf.rf[13][14] ),
    .I2(\dp.rf.rf[14][14] ),
    .I3(\dp.rf.rf[15][14] ),
    .S0(net547),
    .S1(net546),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06784_ (.I0(\dp.rf.rf[4][14] ),
    .I1(\dp.rf.rf[5][14] ),
    .I2(\dp.rf.rf[6][14] ),
    .I3(\dp.rf.rf[7][14] ),
    .S0(net547),
    .S1(net546),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06785_ (.I0(_02246_),
    .I1(_02247_),
    .S(_01066_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06786_ (.A1(_01055_),
    .A2(_02248_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06787_ (.I0(\dp.rf.rf[8][14] ),
    .I1(\dp.rf.rf[9][14] ),
    .I2(\dp.rf.rf[10][14] ),
    .I3(\dp.rf.rf[11][14] ),
    .S0(net547),
    .S1(net546),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06788_ (.I0(\dp.rf.rf[0][14] ),
    .I1(\dp.rf.rf[1][14] ),
    .I2(\dp.rf.rf[2][14] ),
    .I3(\dp.rf.rf[3][14] ),
    .S0(net547),
    .S1(net546),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06789_ (.I0(_02250_),
    .I1(_02251_),
    .S(_01066_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06790_ (.A1(net15),
    .A2(_02252_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _06791_ (.A1(_01064_),
    .A2(_01057_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_4 _06792_ (.A1(_01064_),
    .A2(_02241_),
    .A3(_02245_),
    .B1(_02249_),
    .B2(_02253_),
    .B3(_02254_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06793_ (.I0(_05413_[0]),
    .I1(_02255_),
    .S(_01311_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _06794_ (.A1(_01110_),
    .A2(_02256_),
    .ZN(_05248_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06795_ (.I(_05248_[0]),
    .ZN(_05252_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_310_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_310_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06797_ (.I0(\dp.rf.rf[18][14] ),
    .I1(\dp.rf.rf[19][14] ),
    .I2(\dp.rf.rf[22][14] ),
    .I3(\dp.rf.rf[23][14] ),
    .S0(net538),
    .S1(net9),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06798_ (.I0(\dp.rf.rf[17][14] ),
    .I1(\dp.rf.rf[21][14] ),
    .S(net9),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06799_ (.A1(_01148_),
    .A2(_02259_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06800_ (.A1(\dp.rf.rf[20][14] ),
    .A2(net538),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06801_ (.A1(_02260_),
    .A2(_02261_),
    .B(_01144_),
    .C(net525),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06802_ (.I(\dp.rf.rf[16][14] ),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06803_ (.A1(_02263_),
    .A2(net518),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06804_ (.A1(_01284_),
    .A2(_02258_),
    .B1(_02262_),
    .B2(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06805_ (.I0(\dp.rf.rf[26][14] ),
    .I1(\dp.rf.rf[27][14] ),
    .I2(\dp.rf.rf[30][14] ),
    .I3(\dp.rf.rf[31][14] ),
    .S0(net7),
    .S1(net9),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06806_ (.A1(net8),
    .A2(_02266_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06807_ (.I0(\dp.rf.rf[25][14] ),
    .I1(\dp.rf.rf[29][14] ),
    .S(net9),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06808_ (.A1(net7),
    .A2(_01140_),
    .A3(_02268_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06809_ (.I0(\dp.rf.rf[24][14] ),
    .I1(\dp.rf.rf[28][14] ),
    .S(net9),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06810_ (.A1(_01208_),
    .A2(_02270_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _06811_ (.A1(_01273_),
    .A2(_02267_),
    .A3(_02269_),
    .A4(_02271_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06812_ (.A1(_01216_),
    .A2(_02272_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06813_ (.A1(\dp.rf.rf[4][14] ),
    .A2(net7),
    .A3(_01167_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06814_ (.I0(\dp.rf.rf[1][14] ),
    .I1(\dp.rf.rf[5][14] ),
    .S(net9),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06815_ (.A1(_01148_),
    .A2(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06816_ (.I0(\dp.rf.rf[2][14] ),
    .I1(\dp.rf.rf[3][14] ),
    .I2(\dp.rf.rf[6][14] ),
    .I3(\dp.rf.rf[7][14] ),
    .S0(net7),
    .S1(net9),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06817_ (.I(_02277_),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06818_ (.A1(_02184_),
    .A2(_02274_),
    .A3(_02276_),
    .B1(_02278_),
    .B2(_01232_),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06819_ (.I0(\dp.rf.rf[10][14] ),
    .I1(\dp.rf.rf[11][14] ),
    .I2(\dp.rf.rf[14][14] ),
    .I3(\dp.rf.rf[15][14] ),
    .S0(net7),
    .S1(net9),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06820_ (.I0(\dp.rf.rf[8][14] ),
    .I1(\dp.rf.rf[9][14] ),
    .I2(\dp.rf.rf[12][14] ),
    .I3(\dp.rf.rf[13][14] ),
    .S0(net7),
    .S1(net9),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06821_ (.I0(_02280_),
    .I1(_02281_),
    .S(_01140_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06822_ (.A1(net525),
    .A2(_02279_),
    .B1(_02282_),
    .B2(_01440_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06823_ (.A1(_02265_),
    .A2(_02273_),
    .B(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _06824_ (.I(_02284_),
    .ZN(_05251_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06825_ (.A1(_01089_),
    .A2(_01123_),
    .B1(net528),
    .B2(_01095_),
    .C(_01999_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06826_ (.I0(_02237_),
    .I1(_02285_),
    .S(_01135_),
    .Z(_05409_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06827_ (.I0(\dp.rf.rf[24][13] ),
    .I1(\dp.rf.rf[25][13] ),
    .I2(\dp.rf.rf[26][13] ),
    .I3(\dp.rf.rf[27][13] ),
    .S0(net547),
    .S1(net546),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06828_ (.I0(\dp.rf.rf[16][13] ),
    .I1(\dp.rf.rf[17][13] ),
    .I2(\dp.rf.rf[18][13] ),
    .I3(\dp.rf.rf[19][13] ),
    .S0(net547),
    .S1(net546),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06829_ (.I0(\dp.rf.rf[28][13] ),
    .I1(\dp.rf.rf[29][13] ),
    .I2(\dp.rf.rf[30][13] ),
    .I3(\dp.rf.rf[31][13] ),
    .S0(net547),
    .S1(net546),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06830_ (.I0(\dp.rf.rf[20][13] ),
    .I1(\dp.rf.rf[21][13] ),
    .I2(\dp.rf.rf[22][13] ),
    .I3(\dp.rf.rf[23][13] ),
    .S0(net547),
    .S1(net546),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06831_ (.I0(_02286_),
    .I1(_02287_),
    .I2(_02288_),
    .I3(_02289_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06832_ (.I0(\dp.rf.rf[12][13] ),
    .I1(\dp.rf.rf[13][13] ),
    .I2(\dp.rf.rf[14][13] ),
    .I3(\dp.rf.rf[15][13] ),
    .S0(net547),
    .S1(net546),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06833_ (.I0(\dp.rf.rf[8][13] ),
    .I1(\dp.rf.rf[9][13] ),
    .I2(\dp.rf.rf[10][13] ),
    .I3(\dp.rf.rf[11][13] ),
    .S0(net547),
    .S1(net546),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06834_ (.I0(\dp.rf.rf[4][13] ),
    .I1(\dp.rf.rf[5][13] ),
    .I2(\dp.rf.rf[6][13] ),
    .I3(\dp.rf.rf[7][13] ),
    .S0(net547),
    .S1(net546),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06835_ (.I0(\dp.rf.rf[0][13] ),
    .I1(\dp.rf.rf[1][13] ),
    .I2(\dp.rf.rf[2][13] ),
    .I3(\dp.rf.rf[3][13] ),
    .S0(net547),
    .S1(net546),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06836_ (.I0(_02291_),
    .I1(_02292_),
    .I2(_02293_),
    .I3(_02294_),
    .S0(_01055_),
    .S1(_01066_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06837_ (.I0(_02290_),
    .I1(_02295_),
    .S(_01064_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06838_ (.A1(_01329_),
    .A2(_02296_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06839_ (.A1(_01311_),
    .A2(_02297_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06840_ (.A1(_01119_),
    .A2(_05409_[0]),
    .B(_02298_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06841_ (.A1(_01110_),
    .A2(_02299_),
    .Z(_05256_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06842_ (.I(_05256_[0]),
    .ZN(_05260_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06843_ (.I0(\dp.rf.rf[2][13] ),
    .I1(\dp.rf.rf[3][13] ),
    .I2(\dp.rf.rf[6][13] ),
    .I3(\dp.rf.rf[7][13] ),
    .S0(net7),
    .S1(net534),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06844_ (.I(\dp.rf.rf[4][13] ),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06845_ (.I0(\dp.rf.rf[1][13] ),
    .I1(\dp.rf.rf[5][13] ),
    .S(net534),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06846_ (.A1(_01148_),
    .A2(_02302_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06847_ (.A1(_02301_),
    .A2(_01451_),
    .B(_02184_),
    .C(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06848_ (.A1(_01534_),
    .A2(_02300_),
    .B(_02304_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06849_ (.I0(\dp.rf.rf[10][13] ),
    .I1(\dp.rf.rf[11][13] ),
    .I2(\dp.rf.rf[14][13] ),
    .I3(\dp.rf.rf[15][13] ),
    .S0(net7),
    .S1(net534),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06850_ (.I0(\dp.rf.rf[8][13] ),
    .I1(\dp.rf.rf[9][13] ),
    .I2(\dp.rf.rf[12][13] ),
    .I3(\dp.rf.rf[13][13] ),
    .S0(net7),
    .S1(net534),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06851_ (.I0(_02306_),
    .I1(_02307_),
    .S(_01140_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06852_ (.A1(_01440_),
    .A2(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06853_ (.A1(_01165_),
    .A2(_02305_),
    .B(_02309_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06854_ (.I0(\dp.rf.rf[22][13] ),
    .I1(\dp.rf.rf[23][13] ),
    .S(net538),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06855_ (.A1(\dp.rf.rf[18][13] ),
    .A2(_01368_),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06856_ (.A1(\dp.rf.rf[19][13] ),
    .A2(net538),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06857_ (.A1(net522),
    .A2(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06858_ (.A1(_01167_),
    .A2(_02311_),
    .B1(_02312_),
    .B2(_02314_),
    .C(_01284_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06859_ (.I(\dp.rf.rf[20][13] ),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06860_ (.I0(\dp.rf.rf[17][13] ),
    .I1(\dp.rf.rf[21][13] ),
    .S(net534),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06861_ (.A1(_01148_),
    .A2(_02317_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06862_ (.A1(_02316_),
    .A2(_01451_),
    .B(_02318_),
    .C(net8),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _06863_ (.A1(\dp.rf.rf[16][13] ),
    .A2(_01467_),
    .B1(_02319_),
    .B2(net524),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06864_ (.I0(\dp.rf.rf[26][13] ),
    .I1(\dp.rf.rf[27][13] ),
    .I2(\dp.rf.rf[30][13] ),
    .I3(\dp.rf.rf[31][13] ),
    .S0(net538),
    .S1(net534),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06865_ (.A1(net8),
    .A2(_02321_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06866_ (.I0(\dp.rf.rf[24][13] ),
    .I1(\dp.rf.rf[28][13] ),
    .S(net534),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06867_ (.I0(\dp.rf.rf[25][13] ),
    .I1(\dp.rf.rf[29][13] ),
    .S(net534),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06868_ (.A1(_01208_),
    .A2(_02323_),
    .B1(_02324_),
    .B2(_01585_),
    .C(_01273_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06869_ (.A1(_02315_),
    .A2(_02320_),
    .B1(_02322_),
    .B2(_02325_),
    .C(net514),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _06870_ (.A1(_02310_),
    .A2(_02326_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _06871_ (.I(_02327_),
    .ZN(_05259_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06872_ (.I0(\dp.rf.rf[24][12] ),
    .I1(\dp.rf.rf[25][12] ),
    .I2(\dp.rf.rf[26][12] ),
    .I3(\dp.rf.rf[27][12] ),
    .S0(net547),
    .S1(net546),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06873_ (.I0(\dp.rf.rf[16][12] ),
    .I1(\dp.rf.rf[17][12] ),
    .I2(\dp.rf.rf[18][12] ),
    .I3(\dp.rf.rf[19][12] ),
    .S0(net547),
    .S1(net546),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06874_ (.I0(_02328_),
    .I1(_02329_),
    .S(_01066_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06875_ (.A1(_01055_),
    .A2(_02330_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06876_ (.I0(\dp.rf.rf[28][12] ),
    .I1(\dp.rf.rf[29][12] ),
    .I2(\dp.rf.rf[30][12] ),
    .I3(\dp.rf.rf[31][12] ),
    .S0(net547),
    .S1(net546),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06877_ (.I0(\dp.rf.rf[20][12] ),
    .I1(\dp.rf.rf[21][12] ),
    .I2(\dp.rf.rf[22][12] ),
    .I3(\dp.rf.rf[23][12] ),
    .S0(net547),
    .S1(net546),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06878_ (.I0(_02332_),
    .I1(_02333_),
    .S(_01066_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06879_ (.A1(net15),
    .A2(_02334_),
    .B(_01064_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06880_ (.I0(\dp.rf.rf[12][12] ),
    .I1(\dp.rf.rf[13][12] ),
    .I2(\dp.rf.rf[14][12] ),
    .I3(\dp.rf.rf[15][12] ),
    .S0(net547),
    .S1(net546),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06881_ (.I0(\dp.rf.rf[8][12] ),
    .I1(\dp.rf.rf[9][12] ),
    .I2(\dp.rf.rf[10][12] ),
    .I3(\dp.rf.rf[11][12] ),
    .S0(net547),
    .S1(net546),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06882_ (.I0(_02336_),
    .I1(_02337_),
    .S(_01055_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06883_ (.I0(\dp.rf.rf[4][12] ),
    .I1(\dp.rf.rf[5][12] ),
    .I2(\dp.rf.rf[6][12] ),
    .I3(\dp.rf.rf[7][12] ),
    .S0(net547),
    .S1(net546),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06884_ (.I0(\dp.rf.rf[0][12] ),
    .I1(\dp.rf.rf[1][12] ),
    .I2(\dp.rf.rf[2][12] ),
    .I3(\dp.rf.rf[3][12] ),
    .S0(net547),
    .S1(net546),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06885_ (.I0(_02339_),
    .I1(_02340_),
    .S(_01055_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _06886_ (.A1(_01084_),
    .A2(_02338_),
    .B1(_02341_),
    .B2(_01067_),
    .C(_01329_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06887_ (.A1(_02331_),
    .A2(_02335_),
    .B(_02342_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06888_ (.A1(_01095_),
    .A2(_01315_),
    .B(_01999_),
    .ZN(_05405_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06889_ (.A1(_01119_),
    .A2(_05405_[0]),
    .Z(_02344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06890_ (.A1(_01311_),
    .A2(_02343_),
    .B(_02344_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06891_ (.A1(_01110_),
    .A2(_02345_),
    .Z(_05264_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06892_ (.I(_05264_[0]),
    .ZN(_05268_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06893_ (.I0(\dp.rf.rf[22][12] ),
    .I1(\dp.rf.rf[23][12] ),
    .S(net538),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06894_ (.I(_02346_),
    .ZN(_02347_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _06895_ (.A1(net534),
    .A2(_02347_),
    .B(net523),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06896_ (.I(\dp.rf.rf[18][12] ),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _06897_ (.A1(_02349_),
    .A2(net533),
    .A3(_01101_),
    .A4(_01125_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06898_ (.I0(\dp.rf.rf[18][12] ),
    .I1(\dp.rf.rf[19][12] ),
    .S(net538),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06899_ (.I(_02351_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _06900_ (.A1(net522),
    .A2(_02350_),
    .A3(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06901_ (.I0(\dp.rf.rf[17][12] ),
    .I1(\dp.rf.rf[21][12] ),
    .S(net534),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06902_ (.A1(_01148_),
    .A2(_02354_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06903_ (.A1(\dp.rf.rf[20][12] ),
    .A2(net538),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06904_ (.A1(_02355_),
    .A2(_02356_),
    .B(_01144_),
    .C(net526),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06905_ (.I(\dp.rf.rf[16][12] ),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06906_ (.A1(_02358_),
    .A2(net518),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06907_ (.A1(_02348_),
    .A2(_02353_),
    .B1(_02357_),
    .B2(_02359_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06908_ (.I0(\dp.rf.rf[26][12] ),
    .I1(\dp.rf.rf[27][12] ),
    .I2(\dp.rf.rf[30][12] ),
    .I3(\dp.rf.rf[31][12] ),
    .S0(net538),
    .S1(net534),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06909_ (.A1(net8),
    .A2(_02361_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06910_ (.I0(\dp.rf.rf[25][12] ),
    .I1(\dp.rf.rf[29][12] ),
    .S(net534),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06911_ (.A1(net538),
    .A2(_01140_),
    .A3(_02363_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06912_ (.I0(\dp.rf.rf[24][12] ),
    .I1(\dp.rf.rf[28][12] ),
    .S(net534),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06913_ (.A1(_01208_),
    .A2(_02365_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _06914_ (.A1(_01273_),
    .A2(_02364_),
    .A3(_02366_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06915_ (.A1(_02362_),
    .A2(_02367_),
    .B(_01216_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06916_ (.I0(\dp.rf.rf[8][12] ),
    .I1(\dp.rf.rf[9][12] ),
    .I2(\dp.rf.rf[12][12] ),
    .I3(\dp.rf.rf[13][12] ),
    .S0(net539),
    .S1(net534),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06917_ (.A1(_01140_),
    .A2(_02369_),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06918_ (.I0(\dp.rf.rf[11][12] ),
    .I1(\dp.rf.rf[15][12] ),
    .S(net534),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06919_ (.A1(_01697_),
    .A2(_02371_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06920_ (.I0(\dp.rf.rf[10][12] ),
    .I1(\dp.rf.rf[14][12] ),
    .S(net534),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06921_ (.A1(_01148_),
    .A2(net8),
    .A3(_02373_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _06922_ (.A1(_02370_),
    .A2(_02372_),
    .A3(_02374_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06923_ (.I0(\dp.rf.rf[0][12] ),
    .I1(\dp.rf.rf[1][12] ),
    .I2(\dp.rf.rf[4][12] ),
    .I3(\dp.rf.rf[5][12] ),
    .S0(net538),
    .S1(net534),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _06924_ (.A1(_01140_),
    .A2(_02376_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _06925_ (.A1(_01212_),
    .A2(net526),
    .A3(_01198_),
    .A4(_02377_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06926_ (.I0(\dp.rf.rf[2][12] ),
    .I1(\dp.rf.rf[3][12] ),
    .I2(\dp.rf.rf[6][12] ),
    .I3(\dp.rf.rf[7][12] ),
    .S0(net538),
    .S1(net534),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06927_ (.A1(net526),
    .A2(_01534_),
    .A3(_02379_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _06928_ (.A1(_01440_),
    .A2(_02375_),
    .B(_02378_),
    .C(_02380_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _06929_ (.A1(_02360_),
    .A2(_02368_),
    .B(_02381_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_309_clk (.I(clknet_6_55__leaf_clk),
    .Z(clknet_leaf_309_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _06931_ (.I(_02382_),
    .ZN(_05267_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06932_ (.A1(_01107_),
    .A2(_01112_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06933_ (.A1(_01098_),
    .A2(_01115_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06934_ (.A1(_02383_),
    .A2(_02384_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _06935_ (.A1(net25),
    .A2(net528),
    .A3(_02004_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _06936_ (.A1(net13),
    .A2(_01318_),
    .B1(_02385_),
    .B2(net30),
    .C(_02386_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06937_ (.I0(\dp.rf.rf[24][11] ),
    .I1(\dp.rf.rf[25][11] ),
    .I2(\dp.rf.rf[26][11] ),
    .I3(\dp.rf.rf[27][11] ),
    .S0(net547),
    .S1(net546),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06938_ (.I0(\dp.rf.rf[16][11] ),
    .I1(\dp.rf.rf[17][11] ),
    .I2(\dp.rf.rf[18][11] ),
    .I3(\dp.rf.rf[19][11] ),
    .S0(net547),
    .S1(net546),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06939_ (.I0(_02388_),
    .I1(_02389_),
    .S(_01066_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06940_ (.I0(\dp.rf.rf[28][11] ),
    .I1(\dp.rf.rf[29][11] ),
    .I2(\dp.rf.rf[30][11] ),
    .I3(\dp.rf.rf[31][11] ),
    .S0(net547),
    .S1(net546),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06941_ (.I0(\dp.rf.rf[20][11] ),
    .I1(\dp.rf.rf[21][11] ),
    .I2(\dp.rf.rf[22][11] ),
    .I3(\dp.rf.rf[23][11] ),
    .S0(net547),
    .S1(net546),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06942_ (.I0(_02391_),
    .I1(_02392_),
    .S(_01066_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06943_ (.I0(_02390_),
    .I1(_02393_),
    .S(net15),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06944_ (.I0(\dp.rf.rf[8][11] ),
    .I1(\dp.rf.rf[9][11] ),
    .I2(\dp.rf.rf[10][11] ),
    .I3(\dp.rf.rf[11][11] ),
    .S0(net547),
    .S1(net546),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06945_ (.I0(\dp.rf.rf[0][11] ),
    .I1(\dp.rf.rf[1][11] ),
    .I2(\dp.rf.rf[2][11] ),
    .I3(\dp.rf.rf[3][11] ),
    .S0(net547),
    .S1(net546),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06946_ (.I0(_02395_),
    .I1(_02396_),
    .S(_01066_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06947_ (.I0(\dp.rf.rf[12][11] ),
    .I1(\dp.rf.rf[13][11] ),
    .I2(\dp.rf.rf[14][11] ),
    .I3(\dp.rf.rf[15][11] ),
    .S0(net547),
    .S1(net546),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06948_ (.I0(\dp.rf.rf[4][11] ),
    .I1(\dp.rf.rf[5][11] ),
    .I2(\dp.rf.rf[6][11] ),
    .I3(\dp.rf.rf[7][11] ),
    .S0(net547),
    .S1(net546),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06949_ (.I0(_02398_),
    .I1(_02399_),
    .S(_01066_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06950_ (.I0(_02397_),
    .I1(_02400_),
    .S(net15),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06951_ (.A1(net17),
    .A2(_02394_),
    .B1(_02401_),
    .B2(_01309_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06952_ (.I0(_02387_),
    .I1(_02402_),
    .S(_01311_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06953_ (.A1(_01110_),
    .A2(_02403_),
    .Z(_05272_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06954_ (.I(_05272_[0]),
    .ZN(_05276_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06955_ (.I0(\dp.rf.rf[18][11] ),
    .I1(\dp.rf.rf[19][11] ),
    .I2(\dp.rf.rf[22][11] ),
    .I3(\dp.rf.rf[23][11] ),
    .S0(net542),
    .S1(net9),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06956_ (.I0(\dp.rf.rf[17][11] ),
    .I1(\dp.rf.rf[21][11] ),
    .S(net9),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06957_ (.A1(net531),
    .A2(_02405_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _06958_ (.A1(\dp.rf.rf[20][11] ),
    .A2(net542),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _06959_ (.A1(_02406_),
    .A2(_02407_),
    .B(_01144_),
    .C(net525),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06960_ (.I(\dp.rf.rf[16][11] ),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06961_ (.A1(_02409_),
    .A2(net518),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06962_ (.A1(_01284_),
    .A2(_02404_),
    .B1(_02408_),
    .B2(_02410_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06963_ (.I0(\dp.rf.rf[26][11] ),
    .I1(\dp.rf.rf[27][11] ),
    .I2(\dp.rf.rf[30][11] ),
    .I3(\dp.rf.rf[31][11] ),
    .S0(net7),
    .S1(net9),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06964_ (.A1(net8),
    .A2(_02412_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06965_ (.I0(\dp.rf.rf[24][11] ),
    .I1(\dp.rf.rf[28][11] ),
    .S(net9),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06966_ (.I0(\dp.rf.rf[25][11] ),
    .I1(\dp.rf.rf[29][11] ),
    .S(net9),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06967_ (.A1(_01208_),
    .A2(_02414_),
    .B1(_02415_),
    .B2(_01585_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _06968_ (.A1(_01580_),
    .A2(_02413_),
    .A3(_02416_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _06969_ (.A1(\dp.rf.rf[4][11] ),
    .A2(net7),
    .A3(_01167_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06970_ (.I0(\dp.rf.rf[1][11] ),
    .I1(\dp.rf.rf[5][11] ),
    .S(net9),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _06971_ (.A1(_01148_),
    .A2(_02419_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06972_ (.I0(\dp.rf.rf[2][11] ),
    .I1(\dp.rf.rf[3][11] ),
    .I2(\dp.rf.rf[6][11] ),
    .I3(\dp.rf.rf[7][11] ),
    .S0(net7),
    .S1(net9),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06973_ (.I(_02421_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _06974_ (.A1(_02184_),
    .A2(_02418_),
    .A3(_02420_),
    .B1(_02422_),
    .B2(_01232_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06975_ (.I0(\dp.rf.rf[10][11] ),
    .I1(\dp.rf.rf[11][11] ),
    .I2(\dp.rf.rf[14][11] ),
    .I3(\dp.rf.rf[15][11] ),
    .S0(net7),
    .S1(net9),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06976_ (.I0(\dp.rf.rf[8][11] ),
    .I1(\dp.rf.rf[9][11] ),
    .I2(\dp.rf.rf[12][11] ),
    .I3(\dp.rf.rf[13][11] ),
    .S0(net7),
    .S1(net9),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06977_ (.I0(_02424_),
    .I1(_02425_),
    .S(_01140_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _06978_ (.A1(net525),
    .A2(_02423_),
    .B1(_02426_),
    .B2(_01440_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _06979_ (.A1(net514),
    .A2(_02411_),
    .A3(_02417_),
    .B(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _06980_ (.I(_02428_),
    .ZN(_05275_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _06981_ (.A1(net24),
    .A2(net528),
    .Z(_05397_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06982_ (.I0(\dp.rf.rf[24][10] ),
    .I1(\dp.rf.rf[25][10] ),
    .I2(\dp.rf.rf[26][10] ),
    .I3(\dp.rf.rf[27][10] ),
    .S0(net547),
    .S1(net546),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06983_ (.I0(\dp.rf.rf[16][10] ),
    .I1(\dp.rf.rf[17][10] ),
    .I2(\dp.rf.rf[18][10] ),
    .I3(\dp.rf.rf[19][10] ),
    .S0(net547),
    .S1(net546),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06984_ (.I0(_02429_),
    .I1(_02430_),
    .S(_01066_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06985_ (.I0(\dp.rf.rf[28][10] ),
    .I1(\dp.rf.rf[29][10] ),
    .I2(\dp.rf.rf[30][10] ),
    .I3(\dp.rf.rf[31][10] ),
    .S0(net547),
    .S1(net546),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06986_ (.I0(\dp.rf.rf[20][10] ),
    .I1(\dp.rf.rf[21][10] ),
    .I2(\dp.rf.rf[22][10] ),
    .I3(\dp.rf.rf[23][10] ),
    .S0(net547),
    .S1(net546),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06987_ (.I0(_02432_),
    .I1(_02433_),
    .S(_01066_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06988_ (.I0(_02431_),
    .I1(_02434_),
    .S(net15),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06989_ (.I0(\dp.rf.rf[8][10] ),
    .I1(\dp.rf.rf[9][10] ),
    .I2(\dp.rf.rf[10][10] ),
    .I3(\dp.rf.rf[11][10] ),
    .S0(net547),
    .S1(net546),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06990_ (.I0(\dp.rf.rf[0][10] ),
    .I1(\dp.rf.rf[1][10] ),
    .I2(\dp.rf.rf[2][10] ),
    .I3(\dp.rf.rf[3][10] ),
    .S0(net547),
    .S1(net546),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06991_ (.I0(_02436_),
    .I1(_02437_),
    .S(_01066_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06992_ (.I0(\dp.rf.rf[12][10] ),
    .I1(\dp.rf.rf[13][10] ),
    .I2(\dp.rf.rf[14][10] ),
    .I3(\dp.rf.rf[15][10] ),
    .S0(net547),
    .S1(net546),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _06993_ (.I0(\dp.rf.rf[4][10] ),
    .I1(\dp.rf.rf[5][10] ),
    .I2(\dp.rf.rf[6][10] ),
    .I3(\dp.rf.rf[7][10] ),
    .S0(net547),
    .S1(net546),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06994_ (.I0(_02439_),
    .I1(_02440_),
    .S(_01066_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _06995_ (.I0(_02438_),
    .I1(_02441_),
    .S(net15),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _06996_ (.A1(net17),
    .A2(_02435_),
    .B1(_02442_),
    .B2(_01309_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _06997_ (.A1(_01311_),
    .A2(_02443_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _06998_ (.A1(_01311_),
    .A2(_05397_[0]),
    .B(_02444_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _06999_ (.A1(_01110_),
    .A2(_02445_),
    .Z(_05280_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07000_ (.I(_05280_[0]),
    .ZN(_05284_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07001_ (.I0(\dp.rf.rf[18][10] ),
    .I1(\dp.rf.rf[19][10] ),
    .I2(\dp.rf.rf[22][10] ),
    .I3(\dp.rf.rf[23][10] ),
    .S0(net542),
    .S1(net9),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07002_ (.I0(\dp.rf.rf[17][10] ),
    .I1(\dp.rf.rf[21][10] ),
    .S(net9),
    .Z(_02447_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07003_ (.A1(net531),
    .A2(_02447_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07004_ (.A1(\dp.rf.rf[20][10] ),
    .A2(net542),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07005_ (.A1(_02448_),
    .A2(_02449_),
    .B(_01144_),
    .C(net525),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07006_ (.I(\dp.rf.rf[16][10] ),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07007_ (.A1(_02451_),
    .A2(net518),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07008_ (.A1(_01284_),
    .A2(_02446_),
    .B1(_02450_),
    .B2(_02452_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07009_ (.I0(\dp.rf.rf[26][10] ),
    .I1(\dp.rf.rf[27][10] ),
    .I2(\dp.rf.rf[30][10] ),
    .I3(\dp.rf.rf[31][10] ),
    .S0(net7),
    .S1(net9),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07010_ (.A1(net8),
    .A2(_02454_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07011_ (.I0(\dp.rf.rf[24][10] ),
    .I1(\dp.rf.rf[28][10] ),
    .S(net9),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07012_ (.I0(\dp.rf.rf[25][10] ),
    .I1(\dp.rf.rf[29][10] ),
    .S(net9),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07013_ (.A1(_01208_),
    .A2(_02456_),
    .B1(_02457_),
    .B2(_01585_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07014_ (.A1(_01580_),
    .A2(_02455_),
    .A3(_02458_),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07015_ (.A1(\dp.rf.rf[4][10] ),
    .A2(net7),
    .A3(_01167_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07016_ (.I0(\dp.rf.rf[1][10] ),
    .I1(\dp.rf.rf[5][10] ),
    .S(net9),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07017_ (.A1(_01148_),
    .A2(_02461_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07018_ (.I0(\dp.rf.rf[2][10] ),
    .I1(\dp.rf.rf[3][10] ),
    .I2(\dp.rf.rf[6][10] ),
    .I3(\dp.rf.rf[7][10] ),
    .S0(net7),
    .S1(net9),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07019_ (.I(_02463_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _07020_ (.A1(_02184_),
    .A2(_02460_),
    .A3(_02462_),
    .B1(_02464_),
    .B2(_01232_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07021_ (.I0(\dp.rf.rf[10][10] ),
    .I1(\dp.rf.rf[11][10] ),
    .I2(\dp.rf.rf[14][10] ),
    .I3(\dp.rf.rf[15][10] ),
    .S0(net7),
    .S1(net9),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07022_ (.I0(\dp.rf.rf[8][10] ),
    .I1(\dp.rf.rf[9][10] ),
    .I2(\dp.rf.rf[12][10] ),
    .I3(\dp.rf.rf[13][10] ),
    .S0(net7),
    .S1(net9),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07023_ (.I0(_02466_),
    .I1(_02467_),
    .S(_01140_),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07024_ (.A1(net525),
    .A2(_02465_),
    .B1(_02468_),
    .B2(_01440_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07025_ (.A1(net514),
    .A2(_02453_),
    .A3(_02459_),
    .B(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07026_ (.I(_02470_),
    .ZN(_05283_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07027_ (.A1(net22),
    .A2(net527),
    .Z(_05393_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07028_ (.I0(\dp.rf.rf[24][9] ),
    .I1(\dp.rf.rf[25][9] ),
    .I2(\dp.rf.rf[26][9] ),
    .I3(\dp.rf.rf[27][9] ),
    .S0(net13),
    .S1(net14),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07029_ (.I0(\dp.rf.rf[16][9] ),
    .I1(\dp.rf.rf[17][9] ),
    .I2(\dp.rf.rf[18][9] ),
    .I3(\dp.rf.rf[19][9] ),
    .S0(net13),
    .S1(net14),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07030_ (.I0(_02471_),
    .I1(_02472_),
    .S(_01066_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07031_ (.I0(\dp.rf.rf[28][9] ),
    .I1(\dp.rf.rf[29][9] ),
    .I2(\dp.rf.rf[30][9] ),
    .I3(\dp.rf.rf[31][9] ),
    .S0(net13),
    .S1(net14),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07032_ (.I0(\dp.rf.rf[20][9] ),
    .I1(\dp.rf.rf[21][9] ),
    .I2(\dp.rf.rf[22][9] ),
    .I3(\dp.rf.rf[23][9] ),
    .S0(net13),
    .S1(net14),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07033_ (.I0(_02474_),
    .I1(_02475_),
    .S(_01066_),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07034_ (.A1(_01055_),
    .A2(_02476_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07035_ (.A1(net15),
    .A2(_02473_),
    .B(_02477_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07036_ (.I0(\dp.rf.rf[12][9] ),
    .I1(\dp.rf.rf[13][9] ),
    .I2(\dp.rf.rf[14][9] ),
    .I3(\dp.rf.rf[15][9] ),
    .S0(net13),
    .S1(net14),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07037_ (.I0(\dp.rf.rf[8][9] ),
    .I1(\dp.rf.rf[9][9] ),
    .I2(\dp.rf.rf[10][9] ),
    .I3(\dp.rf.rf[11][9] ),
    .S0(net13),
    .S1(net14),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07038_ (.I0(_02479_),
    .I1(_02480_),
    .S(_01055_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07039_ (.I0(\dp.rf.rf[4][9] ),
    .I1(\dp.rf.rf[5][9] ),
    .I2(\dp.rf.rf[6][9] ),
    .I3(\dp.rf.rf[7][9] ),
    .S0(net13),
    .S1(net14),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07040_ (.I0(\dp.rf.rf[0][9] ),
    .I1(\dp.rf.rf[1][9] ),
    .I2(\dp.rf.rf[2][9] ),
    .I3(\dp.rf.rf[3][9] ),
    .S0(net13),
    .S1(net14),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07041_ (.I0(_02482_),
    .I1(_02483_),
    .S(_01055_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07042_ (.A1(_01084_),
    .A2(_02481_),
    .B1(_02484_),
    .B2(_01067_),
    .C(_01329_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07043_ (.A1(net17),
    .A2(_02478_),
    .B(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07044_ (.I0(_05393_[0]),
    .I1(_02486_),
    .S(_01311_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07045_ (.A1(_01110_),
    .A2(_02487_),
    .ZN(_05288_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07046_ (.I(_05288_[0]),
    .ZN(_05292_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07047_ (.I0(\dp.rf.rf[22][9] ),
    .I1(\dp.rf.rf[23][9] ),
    .S(net7),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07048_ (.I(_02488_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07049_ (.A1(net536),
    .A2(_02489_),
    .B(net523),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07050_ (.I(\dp.rf.rf[18][9] ),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07051_ (.A1(_02491_),
    .A2(net533),
    .A3(net532),
    .A4(_01125_),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07052_ (.I0(\dp.rf.rf[18][9] ),
    .I1(\dp.rf.rf[19][9] ),
    .S(net7),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07053_ (.I(_02493_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07054_ (.A1(net521),
    .A2(_02492_),
    .A3(_02494_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07055_ (.I0(\dp.rf.rf[17][9] ),
    .I1(\dp.rf.rf[21][9] ),
    .S(net536),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07056_ (.A1(_01148_),
    .A2(_02496_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07057_ (.A1(\dp.rf.rf[20][9] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07058_ (.A1(_02497_),
    .A2(_02498_),
    .B(_01144_),
    .C(net529),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07059_ (.I(\dp.rf.rf[16][9] ),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07060_ (.A1(_02500_),
    .A2(_01385_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07061_ (.A1(_02490_),
    .A2(_02495_),
    .B1(_02499_),
    .B2(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07062_ (.I0(\dp.rf.rf[26][9] ),
    .I1(\dp.rf.rf[27][9] ),
    .I2(\dp.rf.rf[30][9] ),
    .I3(\dp.rf.rf[31][9] ),
    .S0(net7),
    .S1(net535),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07063_ (.A1(net8),
    .A2(_02503_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07064_ (.I0(\dp.rf.rf[24][9] ),
    .I1(\dp.rf.rf[28][9] ),
    .S(net535),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07065_ (.I0(\dp.rf.rf[25][9] ),
    .I1(\dp.rf.rf[29][9] ),
    .S(net535),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07066_ (.A1(_01208_),
    .A2(_02505_),
    .B1(_02506_),
    .B2(_01585_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07067_ (.A1(_01580_),
    .A2(_02504_),
    .A3(_02507_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07068_ (.I0(\dp.rf.rf[8][9] ),
    .I1(\dp.rf.rf[9][9] ),
    .I2(\dp.rf.rf[12][9] ),
    .I3(\dp.rf.rf[13][9] ),
    .S0(net7),
    .S1(net9),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07069_ (.I0(\dp.rf.rf[1][9] ),
    .I1(\dp.rf.rf[5][9] ),
    .S(net535),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07070_ (.A1(_01148_),
    .A2(_02510_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07071_ (.A1(\dp.rf.rf[4][9] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07072_ (.A1(_02511_),
    .A2(_02512_),
    .B(net529),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07073_ (.I0(\dp.rf.rf[10][9] ),
    .I1(\dp.rf.rf[11][9] ),
    .I2(\dp.rf.rf[14][9] ),
    .I3(\dp.rf.rf[15][9] ),
    .S0(net7),
    .S1(net9),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07074_ (.I0(\dp.rf.rf[2][9] ),
    .I1(\dp.rf.rf[3][9] ),
    .I2(\dp.rf.rf[6][9] ),
    .I3(\dp.rf.rf[7][9] ),
    .S0(net7),
    .S1(net9),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07075_ (.I0(_02514_),
    .I1(_02515_),
    .S(_01144_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07076_ (.A1(_01279_),
    .A2(_02509_),
    .B1(_02513_),
    .B2(_01458_),
    .C1(_01781_),
    .C2(_02516_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07077_ (.A1(_01475_),
    .A2(_02502_),
    .A3(_02508_),
    .B(_02517_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07078_ (.I(_02518_),
    .ZN(_05291_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07079_ (.A1(net21),
    .A2(net527),
    .Z(_05389_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07080_ (.I0(\dp.rf.rf[28][8] ),
    .I1(\dp.rf.rf[29][8] ),
    .I2(\dp.rf.rf[30][8] ),
    .I3(\dp.rf.rf[31][8] ),
    .S0(net13),
    .S1(net14),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07081_ (.I0(\dp.rf.rf[20][8] ),
    .I1(\dp.rf.rf[21][8] ),
    .I2(\dp.rf.rf[22][8] ),
    .I3(\dp.rf.rf[23][8] ),
    .S0(net13),
    .S1(net14),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07082_ (.I0(\dp.rf.rf[24][8] ),
    .I1(\dp.rf.rf[25][8] ),
    .I2(\dp.rf.rf[26][8] ),
    .I3(\dp.rf.rf[27][8] ),
    .S0(net13),
    .S1(net14),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07083_ (.I0(\dp.rf.rf[16][8] ),
    .I1(\dp.rf.rf[17][8] ),
    .I2(\dp.rf.rf[18][8] ),
    .I3(\dp.rf.rf[19][8] ),
    .S0(net13),
    .S1(net14),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07084_ (.I0(_02519_),
    .I1(_02520_),
    .I2(_02521_),
    .I3(_02522_),
    .S0(_01066_),
    .S1(_01055_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07085_ (.I0(\dp.rf.rf[4][8] ),
    .I1(\dp.rf.rf[5][8] ),
    .I2(\dp.rf.rf[6][8] ),
    .I3(\dp.rf.rf[7][8] ),
    .S0(net13),
    .S1(net14),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07086_ (.I0(\dp.rf.rf[0][8] ),
    .I1(\dp.rf.rf[1][8] ),
    .I2(\dp.rf.rf[2][8] ),
    .I3(\dp.rf.rf[3][8] ),
    .S0(net13),
    .S1(net14),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07087_ (.I0(_02524_),
    .I1(_02525_),
    .S(_01055_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07088_ (.I0(\dp.rf.rf[12][8] ),
    .I1(\dp.rf.rf[13][8] ),
    .I2(\dp.rf.rf[14][8] ),
    .I3(\dp.rf.rf[15][8] ),
    .S0(net13),
    .S1(net14),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07089_ (.I0(\dp.rf.rf[8][8] ),
    .I1(\dp.rf.rf[9][8] ),
    .I2(\dp.rf.rf[10][8] ),
    .I3(\dp.rf.rf[11][8] ),
    .S0(net13),
    .S1(net14),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07090_ (.I0(_02527_),
    .I1(_02528_),
    .S(_01055_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07091_ (.A1(_01084_),
    .A2(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07092_ (.A1(_01329_),
    .A2(_02530_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _07093_ (.A1(_01064_),
    .A2(_02523_),
    .B1(_02526_),
    .B2(_01067_),
    .C(_02531_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07094_ (.I(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07095_ (.I0(_05389_[0]),
    .I1(_02533_),
    .S(_01311_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07096_ (.A1(_01110_),
    .A2(_02534_),
    .ZN(_05296_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07097_ (.I(_05296_[0]),
    .ZN(_05300_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07098_ (.I0(\dp.rf.rf[2][8] ),
    .I1(\dp.rf.rf[3][8] ),
    .I2(\dp.rf.rf[6][8] ),
    .I3(\dp.rf.rf[7][8] ),
    .S0(net7),
    .S1(net9),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07099_ (.I(_02535_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07100_ (.I0(\dp.rf.rf[1][8] ),
    .I1(\dp.rf.rf[5][8] ),
    .S(net9),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07101_ (.A1(\dp.rf.rf[4][8] ),
    .A2(_01245_),
    .B1(_02537_),
    .B2(_01148_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07102_ (.I0(_02536_),
    .I1(_02538_),
    .S(_01140_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07103_ (.I0(\dp.rf.rf[26][8] ),
    .I1(\dp.rf.rf[27][8] ),
    .S(net7),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07104_ (.I(_02540_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07105_ (.I0(\dp.rf.rf[30][8] ),
    .I1(\dp.rf.rf[31][8] ),
    .S(net7),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07106_ (.A1(_01167_),
    .A2(_02542_),
    .B(net8),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07107_ (.A1(net522),
    .A2(_02541_),
    .B(_02543_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07108_ (.I0(\dp.rf.rf[24][8] ),
    .I1(\dp.rf.rf[25][8] ),
    .I2(\dp.rf.rf[28][8] ),
    .I3(\dp.rf.rf[29][8] ),
    .S0(net7),
    .S1(net9),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07109_ (.A1(_01140_),
    .A2(_02545_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07110_ (.A1(net519),
    .A2(_02544_),
    .A3(_02546_),
    .B(_01216_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07111_ (.I0(\dp.rf.rf[18][8] ),
    .I1(\dp.rf.rf[19][8] ),
    .I2(\dp.rf.rf[22][8] ),
    .I3(\dp.rf.rf[23][8] ),
    .S0(net540),
    .S1(net9),
    .Z(_02548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07112_ (.I0(\dp.rf.rf[17][8] ),
    .I1(\dp.rf.rf[21][8] ),
    .S(net9),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07113_ (.A1(_01148_),
    .A2(_02549_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07114_ (.A1(\dp.rf.rf[20][8] ),
    .A2(net540),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07115_ (.A1(_02550_),
    .A2(_02551_),
    .B(_01144_),
    .C(net165),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07116_ (.I(\dp.rf.rf[16][8] ),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07117_ (.A1(_02553_),
    .A2(net518),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07118_ (.A1(_01284_),
    .A2(_02548_),
    .B1(_02552_),
    .B2(_02554_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07119_ (.I0(\dp.rf.rf[10][8] ),
    .I1(\dp.rf.rf[11][8] ),
    .I2(\dp.rf.rf[14][8] ),
    .I3(\dp.rf.rf[15][8] ),
    .S0(net7),
    .S1(net9),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07120_ (.I0(\dp.rf.rf[8][8] ),
    .I1(\dp.rf.rf[9][8] ),
    .I2(\dp.rf.rf[12][8] ),
    .I3(\dp.rf.rf[13][8] ),
    .S0(net7),
    .S1(net9),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07121_ (.I0(_02556_),
    .I1(_02557_),
    .S(_01140_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07122_ (.A1(_01440_),
    .A2(_02558_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _07123_ (.A1(net516),
    .A2(_02539_),
    .B1(_02547_),
    .B2(_02555_),
    .C(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07124_ (.I(net507),
    .ZN(_05299_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07125_ (.I0(\dp.rf.rf[24][7] ),
    .I1(\dp.rf.rf[25][7] ),
    .I2(\dp.rf.rf[26][7] ),
    .I3(\dp.rf.rf[27][7] ),
    .S0(net547),
    .S1(net546),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07126_ (.I0(\dp.rf.rf[16][7] ),
    .I1(\dp.rf.rf[17][7] ),
    .I2(\dp.rf.rf[18][7] ),
    .I3(\dp.rf.rf[19][7] ),
    .S0(net547),
    .S1(net546),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07127_ (.I0(\dp.rf.rf[28][7] ),
    .I1(\dp.rf.rf[29][7] ),
    .I2(\dp.rf.rf[30][7] ),
    .I3(\dp.rf.rf[31][7] ),
    .S0(net547),
    .S1(net546),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07128_ (.I0(\dp.rf.rf[20][7] ),
    .I1(\dp.rf.rf[21][7] ),
    .I2(\dp.rf.rf[22][7] ),
    .I3(\dp.rf.rf[23][7] ),
    .S0(net547),
    .S1(net546),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07129_ (.I0(_02561_),
    .I1(_02562_),
    .I2(_02563_),
    .I3(_02564_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02565_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07130_ (.I0(\dp.rf.rf[8][7] ),
    .I1(\dp.rf.rf[9][7] ),
    .I2(\dp.rf.rf[10][7] ),
    .I3(\dp.rf.rf[11][7] ),
    .S0(net547),
    .S1(net546),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07131_ (.I0(\dp.rf.rf[0][7] ),
    .I1(\dp.rf.rf[1][7] ),
    .I2(\dp.rf.rf[2][7] ),
    .I3(\dp.rf.rf[3][7] ),
    .S0(net547),
    .S1(net546),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07132_ (.I0(\dp.rf.rf[12][7] ),
    .I1(\dp.rf.rf[13][7] ),
    .I2(\dp.rf.rf[14][7] ),
    .I3(\dp.rf.rf[15][7] ),
    .S0(net547),
    .S1(net546),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07133_ (.I0(\dp.rf.rf[4][7] ),
    .I1(\dp.rf.rf[5][7] ),
    .I2(\dp.rf.rf[6][7] ),
    .I3(\dp.rf.rf[7][7] ),
    .S0(net547),
    .S1(net546),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07134_ (.I0(_02566_),
    .I1(_02567_),
    .I2(_02568_),
    .I3(_02569_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07135_ (.I0(_02565_),
    .I1(_02570_),
    .S(_01064_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07136_ (.A1(_01329_),
    .A2(_02571_),
    .Z(net162));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07137_ (.A1(net20),
    .A2(net527),
    .Z(_05385_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07138_ (.I0(net162),
    .I1(_05385_[0]),
    .S(_01119_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07139_ (.A1(_01110_),
    .A2(_02572_),
    .ZN(_05304_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07140_ (.I(_05304_[0]),
    .ZN(_05308_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07141_ (.I0(\dp.rf.rf[2][7] ),
    .I1(\dp.rf.rf[3][7] ),
    .I2(\dp.rf.rf[6][7] ),
    .I3(\dp.rf.rf[7][7] ),
    .S0(net539),
    .S1(net534),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07142_ (.I(_02573_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07143_ (.I0(\dp.rf.rf[1][7] ),
    .I1(\dp.rf.rf[5][7] ),
    .S(net534),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07144_ (.A1(\dp.rf.rf[4][7] ),
    .A2(_01245_),
    .B1(_02575_),
    .B2(_01148_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07145_ (.I0(_02574_),
    .I1(_02576_),
    .S(_01140_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07146_ (.I0(\dp.rf.rf[10][7] ),
    .I1(\dp.rf.rf[11][7] ),
    .I2(\dp.rf.rf[14][7] ),
    .I3(\dp.rf.rf[15][7] ),
    .S0(net539),
    .S1(net534),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07147_ (.I0(\dp.rf.rf[8][7] ),
    .I1(\dp.rf.rf[9][7] ),
    .I2(\dp.rf.rf[12][7] ),
    .I3(\dp.rf.rf[13][7] ),
    .S0(net539),
    .S1(net534),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07148_ (.I0(_02578_),
    .I1(_02579_),
    .S(_01140_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07149_ (.A1(_01440_),
    .A2(_02580_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07150_ (.A1(_01242_),
    .A2(_02577_),
    .B(_02581_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07151_ (.I0(\dp.rf.rf[22][7] ),
    .I1(\dp.rf.rf[23][7] ),
    .S(net538),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07152_ (.A1(\dp.rf.rf[18][7] ),
    .A2(_01368_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07153_ (.A1(\dp.rf.rf[19][7] ),
    .A2(net538),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07154_ (.A1(net522),
    .A2(_02585_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07155_ (.A1(_01167_),
    .A2(_02583_),
    .B1(_02584_),
    .B2(_02586_),
    .C(_01284_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07156_ (.I(\dp.rf.rf[20][7] ),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07157_ (.I0(\dp.rf.rf[17][7] ),
    .I1(\dp.rf.rf[21][7] ),
    .S(net534),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07158_ (.A1(_01148_),
    .A2(_02589_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07159_ (.A1(_02588_),
    .A2(_01451_),
    .B(_02590_),
    .C(net8),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07160_ (.A1(\dp.rf.rf[16][7] ),
    .A2(_01467_),
    .B1(_02591_),
    .B2(_01177_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07161_ (.I0(\dp.rf.rf[26][7] ),
    .I1(\dp.rf.rf[27][7] ),
    .I2(\dp.rf.rf[30][7] ),
    .I3(\dp.rf.rf[31][7] ),
    .S0(net539),
    .S1(net534),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07162_ (.I0(\dp.rf.rf[24][7] ),
    .I1(\dp.rf.rf[25][7] ),
    .I2(\dp.rf.rf[28][7] ),
    .I3(\dp.rf.rf[29][7] ),
    .S0(net539),
    .S1(net534),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07163_ (.I0(_02593_),
    .I1(_02594_),
    .S(_01140_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07164_ (.A1(_01144_),
    .A2(_02595_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _07165_ (.A1(_02587_),
    .A2(_02592_),
    .B(net514),
    .C(_02596_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07166_ (.A1(_02582_),
    .A2(_02597_),
    .Z(_05303_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _07167_ (.I(_05303_[0]),
    .ZN(_05307_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07168_ (.I0(\dp.rf.rf[24][6] ),
    .I1(\dp.rf.rf[25][6] ),
    .I2(\dp.rf.rf[26][6] ),
    .I3(\dp.rf.rf[27][6] ),
    .S0(net549),
    .S1(net14),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07169_ (.I0(\dp.rf.rf[16][6] ),
    .I1(\dp.rf.rf[17][6] ),
    .I2(\dp.rf.rf[18][6] ),
    .I3(\dp.rf.rf[19][6] ),
    .S0(net13),
    .S1(net546),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07170_ (.I0(_02598_),
    .I1(_02599_),
    .S(_01066_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07171_ (.I0(\dp.rf.rf[28][6] ),
    .I1(\dp.rf.rf[29][6] ),
    .I2(\dp.rf.rf[30][6] ),
    .I3(\dp.rf.rf[31][6] ),
    .S0(net549),
    .S1(net14),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07172_ (.I0(\dp.rf.rf[20][6] ),
    .I1(\dp.rf.rf[21][6] ),
    .I2(\dp.rf.rf[22][6] ),
    .I3(\dp.rf.rf[23][6] ),
    .S0(net13),
    .S1(net546),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07173_ (.I0(_02601_),
    .I1(_02602_),
    .S(_01066_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07174_ (.I0(_02600_),
    .I1(_02603_),
    .S(net15),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07175_ (.I0(\dp.rf.rf[8][6] ),
    .I1(\dp.rf.rf[9][6] ),
    .I2(\dp.rf.rf[10][6] ),
    .I3(\dp.rf.rf[11][6] ),
    .S0(net549),
    .S1(net14),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07176_ (.I0(\dp.rf.rf[0][6] ),
    .I1(\dp.rf.rf[1][6] ),
    .I2(\dp.rf.rf[2][6] ),
    .I3(\dp.rf.rf[3][6] ),
    .S0(net13),
    .S1(net14),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07177_ (.I0(_02605_),
    .I1(_02606_),
    .S(_01066_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07178_ (.I0(\dp.rf.rf[12][6] ),
    .I1(\dp.rf.rf[13][6] ),
    .I2(\dp.rf.rf[14][6] ),
    .I3(\dp.rf.rf[15][6] ),
    .S0(net549),
    .S1(net14),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07179_ (.I0(\dp.rf.rf[4][6] ),
    .I1(\dp.rf.rf[5][6] ),
    .I2(\dp.rf.rf[6][6] ),
    .I3(\dp.rf.rf[7][6] ),
    .S0(net550),
    .S1(net14),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07180_ (.I0(_02608_),
    .I1(_02609_),
    .S(_01066_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07181_ (.I0(_02607_),
    .I1(_02610_),
    .S(net15),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _07182_ (.A1(net17),
    .A2(_02604_),
    .B1(_02611_),
    .B2(_01309_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07183_ (.I(_02612_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07184_ (.A1(net19),
    .A2(net527),
    .Z(_05381_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07185_ (.A1(_01311_),
    .A2(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07186_ (.A1(_01311_),
    .A2(_05381_[0]),
    .B(_02613_),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _07187_ (.A1(_01110_),
    .A2(_02614_),
    .Z(_05312_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07188_ (.I(_05312_[0]),
    .ZN(_05316_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07189_ (.I0(\dp.rf.rf[22][6] ),
    .I1(\dp.rf.rf[23][6] ),
    .S(net7),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07190_ (.I(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07191_ (.A1(net537),
    .A2(_02616_),
    .B(net523),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07192_ (.I(\dp.rf.rf[18][6] ),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07193_ (.A1(_02618_),
    .A2(_01030_),
    .A3(_01101_),
    .A4(_01125_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07194_ (.I0(\dp.rf.rf[18][6] ),
    .I1(\dp.rf.rf[19][6] ),
    .S(net7),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07195_ (.I(_02620_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07196_ (.A1(net522),
    .A2(_02619_),
    .A3(_02621_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07197_ (.I0(\dp.rf.rf[17][6] ),
    .I1(\dp.rf.rf[21][6] ),
    .S(net9),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07198_ (.A1(_01148_),
    .A2(_02623_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07199_ (.A1(\dp.rf.rf[20][6] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07200_ (.A1(_02624_),
    .A2(_02625_),
    .B(_01144_),
    .C(net165),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07201_ (.I(\dp.rf.rf[16][6] ),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07202_ (.A1(_02627_),
    .A2(net518),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07203_ (.A1(_02617_),
    .A2(_02622_),
    .B1(_02626_),
    .B2(_02628_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07204_ (.I0(\dp.rf.rf[24][6] ),
    .I1(\dp.rf.rf[25][6] ),
    .I2(\dp.rf.rf[28][6] ),
    .I3(\dp.rf.rf[29][6] ),
    .S0(net7),
    .S1(net9),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07205_ (.A1(_01140_),
    .A2(_02630_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07206_ (.I0(\dp.rf.rf[27][6] ),
    .I1(\dp.rf.rf[31][6] ),
    .S(net9),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07207_ (.I0(\dp.rf.rf[26][6] ),
    .I1(\dp.rf.rf[30][6] ),
    .S(net9),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07208_ (.A1(_01697_),
    .A2(_02632_),
    .B1(_02633_),
    .B2(_01702_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07209_ (.A1(_01580_),
    .A2(_02631_),
    .A3(_02634_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07210_ (.I0(\dp.rf.rf[10][6] ),
    .I1(\dp.rf.rf[11][6] ),
    .I2(\dp.rf.rf[14][6] ),
    .I3(\dp.rf.rf[15][6] ),
    .S0(net7),
    .S1(net9),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07211_ (.I0(\dp.rf.rf[8][6] ),
    .I1(\dp.rf.rf[9][6] ),
    .I2(\dp.rf.rf[12][6] ),
    .I3(\dp.rf.rf[13][6] ),
    .S0(net7),
    .S1(net9),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07212_ (.I0(_02636_),
    .I1(_02637_),
    .S(_01140_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07213_ (.I0(\dp.rf.rf[2][6] ),
    .I1(\dp.rf.rf[3][6] ),
    .I2(\dp.rf.rf[6][6] ),
    .I3(\dp.rf.rf[7][6] ),
    .S0(net7),
    .S1(net9),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07214_ (.I0(\dp.rf.rf[1][6] ),
    .I1(\dp.rf.rf[5][6] ),
    .S(net9),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07215_ (.A1(_01148_),
    .A2(_02640_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07216_ (.A1(\dp.rf.rf[4][6] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07217_ (.A1(_02641_),
    .A2(_02642_),
    .B(net529),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07218_ (.A1(_01440_),
    .A2(_02638_),
    .B1(_02639_),
    .B2(_01535_),
    .C1(_01458_),
    .C2(_02643_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07219_ (.A1(net515),
    .A2(_02629_),
    .A3(_02635_),
    .B(_02644_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _07220_ (.I(_02645_),
    .ZN(_05315_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07221_ (.I0(\dp.rf.rf[24][5] ),
    .I1(\dp.rf.rf[25][5] ),
    .I2(\dp.rf.rf[26][5] ),
    .I3(\dp.rf.rf[27][5] ),
    .S0(net547),
    .S1(net546),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07222_ (.I0(\dp.rf.rf[16][5] ),
    .I1(\dp.rf.rf[17][5] ),
    .I2(\dp.rf.rf[18][5] ),
    .I3(\dp.rf.rf[19][5] ),
    .S0(net547),
    .S1(net546),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07223_ (.I0(_02646_),
    .I1(_02647_),
    .S(_01066_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07224_ (.I0(\dp.rf.rf[28][5] ),
    .I1(\dp.rf.rf[29][5] ),
    .I2(\dp.rf.rf[30][5] ),
    .I3(\dp.rf.rf[31][5] ),
    .S0(net547),
    .S1(net546),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07225_ (.I0(\dp.rf.rf[20][5] ),
    .I1(\dp.rf.rf[21][5] ),
    .I2(\dp.rf.rf[22][5] ),
    .I3(\dp.rf.rf[23][5] ),
    .S0(net547),
    .S1(net546),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07226_ (.I0(_02649_),
    .I1(_02650_),
    .S(_01066_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07227_ (.I0(_02648_),
    .I1(_02651_),
    .S(net15),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07228_ (.I0(\dp.rf.rf[8][5] ),
    .I1(\dp.rf.rf[9][5] ),
    .I2(\dp.rf.rf[10][5] ),
    .I3(\dp.rf.rf[11][5] ),
    .S0(net547),
    .S1(net546),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07229_ (.I0(\dp.rf.rf[0][5] ),
    .I1(\dp.rf.rf[1][5] ),
    .I2(\dp.rf.rf[2][5] ),
    .I3(\dp.rf.rf[3][5] ),
    .S0(net547),
    .S1(net546),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07230_ (.I0(_02653_),
    .I1(_02654_),
    .S(_01066_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07231_ (.I0(\dp.rf.rf[12][5] ),
    .I1(\dp.rf.rf[13][5] ),
    .I2(\dp.rf.rf[14][5] ),
    .I3(\dp.rf.rf[15][5] ),
    .S0(net547),
    .S1(net546),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07232_ (.I0(\dp.rf.rf[4][5] ),
    .I1(\dp.rf.rf[5][5] ),
    .I2(\dp.rf.rf[6][5] ),
    .I3(\dp.rf.rf[7][5] ),
    .S0(net547),
    .S1(net546),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07233_ (.I0(_02656_),
    .I1(_02657_),
    .S(_01066_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07234_ (.I0(_02655_),
    .I1(_02658_),
    .S(net15),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07235_ (.A1(net17),
    .A2(_02652_),
    .B1(_02659_),
    .B2(_01309_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _07236_ (.I(_02660_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07237_ (.A1(net18),
    .A2(net527),
    .Z(_05377_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07238_ (.I0(net160),
    .I1(_05377_[0]),
    .S(_01119_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07239_ (.A1(_01110_),
    .A2(_02661_),
    .ZN(_05320_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07240_ (.I(_05320_[0]),
    .ZN(_05324_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07241_ (.I0(\dp.rf.rf[2][5] ),
    .I1(\dp.rf.rf[3][5] ),
    .I2(\dp.rf.rf[6][5] ),
    .I3(\dp.rf.rf[7][5] ),
    .S0(net539),
    .S1(net534),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07242_ (.I(_02662_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07243_ (.I0(\dp.rf.rf[1][5] ),
    .I1(\dp.rf.rf[5][5] ),
    .S(net534),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07244_ (.A1(\dp.rf.rf[4][5] ),
    .A2(_01245_),
    .B1(_02664_),
    .B2(_01148_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07245_ (.I0(_02663_),
    .I1(_02665_),
    .S(_01140_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07246_ (.I0(\dp.rf.rf[18][5] ),
    .I1(\dp.rf.rf[19][5] ),
    .I2(\dp.rf.rf[22][5] ),
    .I3(\dp.rf.rf[23][5] ),
    .S0(net538),
    .S1(net534),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07247_ (.I0(\dp.rf.rf[17][5] ),
    .I1(\dp.rf.rf[21][5] ),
    .S(net534),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07248_ (.A1(_01148_),
    .A2(_02668_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07249_ (.A1(\dp.rf.rf[20][5] ),
    .A2(net538),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07250_ (.A1(_02669_),
    .A2(_02670_),
    .B(_01144_),
    .C(net526),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07251_ (.I(\dp.rf.rf[16][5] ),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07252_ (.A1(_02672_),
    .A2(net518),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07253_ (.A1(_01284_),
    .A2(_02667_),
    .B1(_02671_),
    .B2(_02673_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07254_ (.I0(\dp.rf.rf[26][5] ),
    .I1(\dp.rf.rf[27][5] ),
    .I2(\dp.rf.rf[30][5] ),
    .I3(\dp.rf.rf[31][5] ),
    .S0(net538),
    .S1(net534),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07255_ (.I0(\dp.rf.rf[24][5] ),
    .I1(\dp.rf.rf[25][5] ),
    .I2(\dp.rf.rf[28][5] ),
    .I3(\dp.rf.rf[29][5] ),
    .S0(net538),
    .S1(net534),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07256_ (.I0(_02675_),
    .I1(_02676_),
    .S(_01140_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07257_ (.A1(_01144_),
    .A2(_02677_),
    .B(_01216_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07258_ (.I0(\dp.rf.rf[10][5] ),
    .I1(\dp.rf.rf[11][5] ),
    .I2(\dp.rf.rf[14][5] ),
    .I3(\dp.rf.rf[15][5] ),
    .S0(net539),
    .S1(net534),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07259_ (.I0(\dp.rf.rf[8][5] ),
    .I1(\dp.rf.rf[9][5] ),
    .I2(\dp.rf.rf[12][5] ),
    .I3(\dp.rf.rf[13][5] ),
    .S0(net539),
    .S1(net534),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07260_ (.I0(_02679_),
    .I1(_02680_),
    .S(_01140_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07261_ (.A1(_01440_),
    .A2(_02681_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _07262_ (.A1(_01242_),
    .A2(_02666_),
    .B1(_02674_),
    .B2(_02678_),
    .C(_02682_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07263_ (.I(_02683_),
    .ZN(_05323_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _07264_ (.I(net3),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07265_ (.I0(_01064_),
    .I1(_02684_),
    .S(net99),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07266_ (.A1(net3),
    .A2(_01112_),
    .B1(_01122_),
    .B2(net17),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _07267_ (.A1(net27),
    .A2(_01030_),
    .A3(_01104_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _07268_ (.A1(_01165_),
    .A2(_01135_),
    .A3(_02685_),
    .B1(_02686_),
    .B2(_02687_),
    .ZN(_05373_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07269_ (.A1(net17),
    .A2(net15),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07270_ (.I0(\dp.rf.rf[22][4] ),
    .I1(\dp.rf.rf[23][4] ),
    .I2(\dp.rf.rf[30][4] ),
    .I3(\dp.rf.rf[31][4] ),
    .S0(net550),
    .S1(net16),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07271_ (.I0(\dp.rf.rf[20][4] ),
    .I1(\dp.rf.rf[21][4] ),
    .I2(\dp.rf.rf[28][4] ),
    .I3(\dp.rf.rf[29][4] ),
    .S0(net550),
    .S1(net16),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07272_ (.I0(_02689_),
    .I1(_02690_),
    .S(_01036_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07273_ (.I0(\dp.rf.rf[24][4] ),
    .I1(\dp.rf.rf[25][4] ),
    .I2(\dp.rf.rf[26][4] ),
    .I3(\dp.rf.rf[27][4] ),
    .S0(net550),
    .S1(net14),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07274_ (.I0(\dp.rf.rf[16][4] ),
    .I1(\dp.rf.rf[17][4] ),
    .I2(\dp.rf.rf[18][4] ),
    .I3(\dp.rf.rf[19][4] ),
    .S0(net13),
    .S1(net14),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07275_ (.I0(_02692_),
    .I1(_02693_),
    .S(_01066_),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07276_ (.A1(_02688_),
    .A2(_02691_),
    .B1(_02694_),
    .B2(_02105_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07277_ (.I0(\dp.rf.rf[12][4] ),
    .I1(\dp.rf.rf[13][4] ),
    .I2(\dp.rf.rf[14][4] ),
    .I3(\dp.rf.rf[15][4] ),
    .S0(net550),
    .S1(net14),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07278_ (.I0(\dp.rf.rf[8][4] ),
    .I1(\dp.rf.rf[9][4] ),
    .I2(\dp.rf.rf[10][4] ),
    .I3(\dp.rf.rf[11][4] ),
    .S0(net550),
    .S1(net14),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07279_ (.I0(_02696_),
    .I1(_02697_),
    .S(_01055_),
    .Z(_02698_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07280_ (.I0(\dp.rf.rf[2][4] ),
    .I1(\dp.rf.rf[3][4] ),
    .I2(\dp.rf.rf[6][4] ),
    .I3(\dp.rf.rf[7][4] ),
    .S0(net550),
    .S1(net15),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07281_ (.I0(\dp.rf.rf[0][4] ),
    .I1(\dp.rf.rf[1][4] ),
    .I2(\dp.rf.rf[4][4] ),
    .I3(\dp.rf.rf[5][4] ),
    .S0(net550),
    .S1(net15),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07282_ (.I0(_02699_),
    .I1(_02700_),
    .S(_01036_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07283_ (.A1(_01084_),
    .A2(_02698_),
    .B1(_02701_),
    .B2(_01067_),
    .C(_01329_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07284_ (.A1(_02695_),
    .A2(_02702_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07285_ (.I(_02703_),
    .ZN(net159));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07286_ (.I0(_05373_[0]),
    .I1(net159),
    .S(_01311_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_308_clk (.I(clknet_6_55__leaf_clk),
    .Z(clknet_leaf_308_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_307_clk (.I(clknet_6_55__leaf_clk),
    .Z(clknet_leaf_307_clk));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07289_ (.A1(_01110_),
    .A2(_02704_),
    .ZN(_05328_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07290_ (.I(_05328_[0]),
    .ZN(_05332_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07291_ (.I0(\dp.rf.rf[22][4] ),
    .I1(\dp.rf.rf[23][4] ),
    .S(net7),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07292_ (.I(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07293_ (.A1(net536),
    .A2(_02708_),
    .B(net523),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07294_ (.I(\dp.rf.rf[18][4] ),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07295_ (.A1(_02710_),
    .A2(net533),
    .A3(net532),
    .A4(_01125_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07296_ (.I0(\dp.rf.rf[18][4] ),
    .I1(\dp.rf.rf[19][4] ),
    .S(net545),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07297_ (.I(_02712_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07298_ (.A1(net521),
    .A2(_02711_),
    .A3(_02713_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07299_ (.I0(\dp.rf.rf[17][4] ),
    .I1(\dp.rf.rf[21][4] ),
    .S(net536),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07300_ (.A1(_01148_),
    .A2(_02715_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07301_ (.A1(\dp.rf.rf[20][4] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07302_ (.A1(_02716_),
    .A2(_02717_),
    .B(_01144_),
    .C(net529),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07303_ (.I(\dp.rf.rf[16][4] ),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07304_ (.A1(_02719_),
    .A2(_01385_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07305_ (.A1(_02709_),
    .A2(_02714_),
    .B1(_02718_),
    .B2(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07306_ (.I0(\dp.rf.rf[24][4] ),
    .I1(\dp.rf.rf[25][4] ),
    .I2(\dp.rf.rf[28][4] ),
    .I3(\dp.rf.rf[29][4] ),
    .S0(net7),
    .S1(net535),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07307_ (.A1(_01140_),
    .A2(_02722_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07308_ (.I0(\dp.rf.rf[27][4] ),
    .I1(\dp.rf.rf[31][4] ),
    .S(net535),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07309_ (.I0(\dp.rf.rf[26][4] ),
    .I1(\dp.rf.rf[30][4] ),
    .S(net535),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07310_ (.A1(_01697_),
    .A2(_02724_),
    .B1(_02725_),
    .B2(_01702_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07311_ (.A1(_01580_),
    .A2(_02723_),
    .A3(_02726_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07312_ (.I0(\dp.rf.rf[8][4] ),
    .I1(\dp.rf.rf[9][4] ),
    .I2(\dp.rf.rf[12][4] ),
    .I3(\dp.rf.rf[13][4] ),
    .S0(net7),
    .S1(net9),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07313_ (.I0(\dp.rf.rf[1][4] ),
    .I1(\dp.rf.rf[5][4] ),
    .S(net535),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07314_ (.A1(_01148_),
    .A2(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07315_ (.A1(\dp.rf.rf[4][4] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07316_ (.A1(_02730_),
    .A2(_02731_),
    .B(net529),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07317_ (.I0(\dp.rf.rf[10][4] ),
    .I1(\dp.rf.rf[11][4] ),
    .I2(\dp.rf.rf[14][4] ),
    .I3(\dp.rf.rf[15][4] ),
    .S0(net7),
    .S1(net9),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07318_ (.I0(\dp.rf.rf[2][4] ),
    .I1(\dp.rf.rf[3][4] ),
    .I2(\dp.rf.rf[6][4] ),
    .I3(\dp.rf.rf[7][4] ),
    .S0(net7),
    .S1(net9),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07319_ (.I0(_02733_),
    .I1(_02734_),
    .S(_01144_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07320_ (.A1(_01279_),
    .A2(_02728_),
    .B1(_02732_),
    .B2(_01458_),
    .C1(_01781_),
    .C2(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07321_ (.A1(_01475_),
    .A2(_02721_),
    .A3(_02727_),
    .B(_02736_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07322_ (.I(net506),
    .ZN(_05331_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07323_ (.A1(_01066_),
    .A2(_01324_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07324_ (.A1(_02687_),
    .A2(_02686_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07325_ (.A1(net2),
    .A2(net527),
    .B(_01324_),
    .C(_02739_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07326_ (.A1(net2),
    .A2(_01112_),
    .B1(_01122_),
    .B2(net16),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _07327_ (.A1(_01135_),
    .A2(_02738_),
    .A3(_02740_),
    .B1(_02741_),
    .B2(_02687_),
    .ZN(_05367_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07328_ (.I0(\dp.rf.rf[24][3] ),
    .I1(\dp.rf.rf[25][3] ),
    .I2(\dp.rf.rf[26][3] ),
    .I3(\dp.rf.rf[27][3] ),
    .S0(net13),
    .S1(net546),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07329_ (.I0(\dp.rf.rf[16][3] ),
    .I1(\dp.rf.rf[17][3] ),
    .I2(\dp.rf.rf[18][3] ),
    .I3(\dp.rf.rf[19][3] ),
    .S0(net13),
    .S1(net546),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07330_ (.I0(\dp.rf.rf[28][3] ),
    .I1(\dp.rf.rf[29][3] ),
    .I2(\dp.rf.rf[30][3] ),
    .I3(\dp.rf.rf[31][3] ),
    .S0(net13),
    .S1(net546),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07331_ (.I0(\dp.rf.rf[20][3] ),
    .I1(\dp.rf.rf[21][3] ),
    .I2(\dp.rf.rf[22][3] ),
    .I3(\dp.rf.rf[23][3] ),
    .S0(net13),
    .S1(net546),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07332_ (.I0(_02742_),
    .I1(_02743_),
    .I2(_02744_),
    .I3(_02745_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07333_ (.I0(\dp.rf.rf[8][3] ),
    .I1(\dp.rf.rf[9][3] ),
    .I2(\dp.rf.rf[10][3] ),
    .I3(\dp.rf.rf[11][3] ),
    .S0(net13),
    .S1(net546),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07334_ (.I0(\dp.rf.rf[0][3] ),
    .I1(\dp.rf.rf[1][3] ),
    .I2(\dp.rf.rf[2][3] ),
    .I3(\dp.rf.rf[3][3] ),
    .S0(net13),
    .S1(net546),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07335_ (.I0(\dp.rf.rf[12][3] ),
    .I1(\dp.rf.rf[13][3] ),
    .I2(\dp.rf.rf[14][3] ),
    .I3(\dp.rf.rf[15][3] ),
    .S0(net13),
    .S1(net546),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07336_ (.I0(\dp.rf.rf[4][3] ),
    .I1(\dp.rf.rf[5][3] ),
    .I2(\dp.rf.rf[6][3] ),
    .I3(\dp.rf.rf[7][3] ),
    .S0(net13),
    .S1(net546),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07337_ (.I0(_02747_),
    .I1(_02748_),
    .I2(_02749_),
    .I3(_02750_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07338_ (.I0(_02746_),
    .I1(_02751_),
    .S(_01064_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07339_ (.A1(_01329_),
    .A2(_02752_),
    .Z(net158));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07340_ (.I0(_05367_[0]),
    .I1(net158),
    .S(_01311_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_296_clk (.I(clknet_6_52__leaf_clk),
    .Z(clknet_leaf_296_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_295_clk (.I(clknet_6_53__leaf_clk),
    .Z(clknet_leaf_295_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_294_clk (.I(clknet_6_55__leaf_clk),
    .Z(clknet_leaf_294_clk));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07344_ (.A1(_01110_),
    .A2(_02753_),
    .ZN(_05336_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07345_ (.I(_05336_[0]),
    .ZN(_05340_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07346_ (.I0(\dp.rf.rf[26][3] ),
    .I1(\dp.rf.rf[27][3] ),
    .I2(\dp.rf.rf[30][3] ),
    .I3(\dp.rf.rf[31][3] ),
    .S0(net542),
    .S1(net534),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07347_ (.I0(\dp.rf.rf[24][3] ),
    .I1(\dp.rf.rf[25][3] ),
    .I2(\dp.rf.rf[28][3] ),
    .I3(\dp.rf.rf[29][3] ),
    .S0(net542),
    .S1(net534),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07348_ (.I0(_02757_),
    .I1(_02758_),
    .S(_01140_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07349_ (.A1(_01144_),
    .A2(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07350_ (.I0(\dp.rf.rf[22][3] ),
    .I1(\dp.rf.rf[23][3] ),
    .S(net542),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07351_ (.A1(\dp.rf.rf[18][3] ),
    .A2(_01368_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07352_ (.A1(\dp.rf.rf[19][3] ),
    .A2(net542),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07353_ (.A1(net522),
    .A2(_02763_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07354_ (.A1(_01167_),
    .A2(_02761_),
    .B1(_02762_),
    .B2(_02764_),
    .C(_01284_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07355_ (.I(\dp.rf.rf[20][3] ),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07356_ (.I0(\dp.rf.rf[17][3] ),
    .I1(\dp.rf.rf[21][3] ),
    .S(net534),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07357_ (.A1(net531),
    .A2(_02767_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07358_ (.A1(_02766_),
    .A2(_01451_),
    .B(_02768_),
    .C(net8),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07359_ (.A1(\dp.rf.rf[16][3] ),
    .A2(_01467_),
    .B1(_02769_),
    .B2(_01177_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07360_ (.A1(_02765_),
    .A2(_02770_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07361_ (.I0(\dp.rf.rf[10][3] ),
    .I1(\dp.rf.rf[11][3] ),
    .I2(\dp.rf.rf[14][3] ),
    .I3(\dp.rf.rf[15][3] ),
    .S0(net542),
    .S1(net534),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07362_ (.I0(\dp.rf.rf[8][3] ),
    .I1(\dp.rf.rf[9][3] ),
    .I2(\dp.rf.rf[12][3] ),
    .I3(\dp.rf.rf[13][3] ),
    .S0(net542),
    .S1(net534),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07363_ (.I0(_02772_),
    .I1(_02773_),
    .S(_01140_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07364_ (.A1(_01273_),
    .A2(_02774_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07365_ (.A1(\dp.rf.rf[2][3] ),
    .A2(_01368_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07366_ (.A1(\dp.rf.rf[3][3] ),
    .A2(net542),
    .B1(net534),
    .B2(net526),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07367_ (.I0(\dp.rf.rf[6][3] ),
    .I1(\dp.rf.rf[7][3] ),
    .S(net542),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07368_ (.A1(_01167_),
    .A2(_02778_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07369_ (.A1(_02776_),
    .A2(_02777_),
    .B(net523),
    .C(_02779_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07370_ (.I(\dp.rf.rf[0][3] ),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07371_ (.I0(\dp.rf.rf[1][3] ),
    .I1(\dp.rf.rf[5][3] ),
    .S(net534),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07372_ (.A1(\dp.rf.rf[4][3] ),
    .A2(_01245_),
    .B1(_02782_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07373_ (.A1(_02781_),
    .A2(net518),
    .B1(_02783_),
    .B2(_01377_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07374_ (.A1(_02780_),
    .A2(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07375_ (.A1(net10),
    .A2(_01197_),
    .B(_01214_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _07376_ (.A1(net514),
    .A2(_02760_),
    .A3(_02771_),
    .B1(_02775_),
    .B2(_02785_),
    .B3(_02786_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _07377_ (.I(net501),
    .ZN(_05339_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07378_ (.A1(_01055_),
    .A2(_01324_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07379_ (.A1(_02687_),
    .A2(_02741_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07380_ (.A1(net32),
    .A2(net527),
    .B(_01324_),
    .C(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07381_ (.A1(net32),
    .A2(_01112_),
    .B1(_01122_),
    .B2(net15),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _07382_ (.A1(_01135_),
    .A2(_02788_),
    .A3(_02790_),
    .B1(_02791_),
    .B2(_02687_),
    .ZN(_05363_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07383_ (.I0(\dp.rf.rf[28][2] ),
    .I1(\dp.rf.rf[29][2] ),
    .I2(\dp.rf.rf[30][2] ),
    .I3(\dp.rf.rf[31][2] ),
    .S0(net13),
    .S1(net14),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07384_ (.I0(\dp.rf.rf[20][2] ),
    .I1(\dp.rf.rf[21][2] ),
    .I2(\dp.rf.rf[22][2] ),
    .I3(\dp.rf.rf[23][2] ),
    .S0(net13),
    .S1(net14),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07385_ (.I0(\dp.rf.rf[24][2] ),
    .I1(\dp.rf.rf[25][2] ),
    .I2(\dp.rf.rf[26][2] ),
    .I3(\dp.rf.rf[27][2] ),
    .S0(net13),
    .S1(net14),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07386_ (.I0(\dp.rf.rf[16][2] ),
    .I1(\dp.rf.rf[17][2] ),
    .I2(\dp.rf.rf[18][2] ),
    .I3(\dp.rf.rf[19][2] ),
    .S0(net13),
    .S1(net14),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07387_ (.I0(_02792_),
    .I1(_02793_),
    .I2(_02794_),
    .I3(_02795_),
    .S0(_01066_),
    .S1(_01055_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07388_ (.I0(\dp.rf.rf[8][2] ),
    .I1(\dp.rf.rf[9][2] ),
    .I2(\dp.rf.rf[10][2] ),
    .I3(\dp.rf.rf[11][2] ),
    .S0(net13),
    .S1(net14),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07389_ (.I0(\dp.rf.rf[0][2] ),
    .I1(\dp.rf.rf[1][2] ),
    .I2(\dp.rf.rf[2][2] ),
    .I3(\dp.rf.rf[3][2] ),
    .S0(net13),
    .S1(net14),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07390_ (.I0(\dp.rf.rf[12][2] ),
    .I1(\dp.rf.rf[13][2] ),
    .I2(\dp.rf.rf[14][2] ),
    .I3(\dp.rf.rf[15][2] ),
    .S0(net13),
    .S1(net14),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07391_ (.I0(\dp.rf.rf[4][2] ),
    .I1(\dp.rf.rf[5][2] ),
    .I2(\dp.rf.rf[6][2] ),
    .I3(\dp.rf.rf[7][2] ),
    .S0(net13),
    .S1(net14),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07392_ (.I0(_02797_),
    .I1(_02798_),
    .I2(_02799_),
    .I3(_02800_),
    .S0(_01066_),
    .S1(net15),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07393_ (.A1(_01329_),
    .A2(_02801_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07394_ (.I0(_02796_),
    .I1(_02802_),
    .S(_01064_),
    .Z(net155));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07395_ (.I0(_05363_[0]),
    .I1(net155),
    .S(_01311_),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_291_clk (.I(clknet_6_53__leaf_clk),
    .Z(clknet_leaf_291_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_290_clk (.I(clknet_6_53__leaf_clk),
    .Z(clknet_leaf_290_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_284_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_284_clk));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07399_ (.A1(_01110_),
    .A2(_02803_),
    .ZN(_05344_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07400_ (.I(_05344_[0]),
    .ZN(_05348_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07401_ (.I0(\dp.rf.rf[8][2] ),
    .I1(\dp.rf.rf[9][2] ),
    .I2(\dp.rf.rf[12][2] ),
    .I3(\dp.rf.rf[13][2] ),
    .S0(net7),
    .S1(net535),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07402_ (.I0(\dp.rf.rf[10][2] ),
    .I1(\dp.rf.rf[11][2] ),
    .I2(\dp.rf.rf[14][2] ),
    .I3(\dp.rf.rf[15][2] ),
    .S0(net7),
    .S1(net535),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07403_ (.I0(\dp.rf.rf[2][2] ),
    .I1(\dp.rf.rf[3][2] ),
    .I2(\dp.rf.rf[6][2] ),
    .I3(\dp.rf.rf[7][2] ),
    .S0(net7),
    .S1(net535),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07404_ (.I0(_02808_),
    .I1(_02809_),
    .S(_01144_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07405_ (.I0(\dp.rf.rf[1][2] ),
    .I1(\dp.rf.rf[5][2] ),
    .S(net535),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07406_ (.A1(\dp.rf.rf[4][2] ),
    .A2(_01245_),
    .B1(_02811_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07407_ (.A1(net165),
    .A2(_02812_),
    .B(_01242_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07408_ (.A1(_01279_),
    .A2(_02807_),
    .B1(_02810_),
    .B2(_01781_),
    .C(_02813_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07409_ (.I0(\dp.rf.rf[26][2] ),
    .I1(\dp.rf.rf[27][2] ),
    .I2(\dp.rf.rf[30][2] ),
    .I3(\dp.rf.rf[31][2] ),
    .S0(net7),
    .S1(net535),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07410_ (.I0(\dp.rf.rf[24][2] ),
    .I1(\dp.rf.rf[25][2] ),
    .I2(\dp.rf.rf[28][2] ),
    .I3(\dp.rf.rf[29][2] ),
    .S0(net7),
    .S1(net535),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07411_ (.I0(_02815_),
    .I1(_02816_),
    .S(_01140_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07412_ (.I0(\dp.rf.rf[22][2] ),
    .I1(\dp.rf.rf[23][2] ),
    .S(net543),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07413_ (.I(_02818_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07414_ (.A1(\dp.rf.rf[18][2] ),
    .A2(_01368_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07415_ (.A1(\dp.rf.rf[19][2] ),
    .A2(net543),
    .B1(net536),
    .B2(net165),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07416_ (.A1(net536),
    .A2(_02819_),
    .B1(_02820_),
    .B2(_02821_),
    .C(net523),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07417_ (.I(\dp.rf.rf[16][2] ),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07418_ (.I0(\dp.rf.rf[17][2] ),
    .I1(\dp.rf.rf[21][2] ),
    .S(net537),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07419_ (.A1(\dp.rf.rf[20][2] ),
    .A2(_01245_),
    .B1(_02824_),
    .B2(_01148_),
    .C(_01140_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07420_ (.A1(_02823_),
    .A2(_01385_),
    .B1(_02825_),
    .B2(_01377_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07421_ (.A1(net519),
    .A2(_02817_),
    .B1(_02822_),
    .B2(_02826_),
    .C(_01216_),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07422_ (.A1(_02814_),
    .A2(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _07423_ (.I(_02828_),
    .ZN(_05347_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07424_ (.A1(_01033_),
    .A2(_01129_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07425_ (.A1(net546),
    .A2(_01318_),
    .B(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _07426_ (.I(net31),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _07427_ (.A1(_02831_),
    .A2(_01165_),
    .A3(_01135_),
    .B1(_02791_),
    .B2(_02687_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07428_ (.A1(net546),
    .A2(_01317_),
    .A3(_01318_),
    .A4(_01165_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07429_ (.A1(_01324_),
    .A2(_02832_),
    .B(_02833_),
    .C(_02004_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07430_ (.A1(_02830_),
    .A2(_02834_),
    .ZN(_05100_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07431_ (.I0(\dp.rf.rf[12][1] ),
    .I1(\dp.rf.rf[13][1] ),
    .I2(\dp.rf.rf[14][1] ),
    .I3(\dp.rf.rf[15][1] ),
    .S0(net550),
    .S1(net14),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07432_ (.I0(\dp.rf.rf[4][1] ),
    .I1(\dp.rf.rf[5][1] ),
    .I2(\dp.rf.rf[6][1] ),
    .I3(\dp.rf.rf[7][1] ),
    .S0(net550),
    .S1(net14),
    .Z(_02836_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07433_ (.I0(\dp.rf.rf[28][1] ),
    .I1(\dp.rf.rf[29][1] ),
    .I2(\dp.rf.rf[30][1] ),
    .I3(\dp.rf.rf[31][1] ),
    .S0(net550),
    .S1(net14),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07434_ (.I0(\dp.rf.rf[20][1] ),
    .I1(\dp.rf.rf[21][1] ),
    .I2(\dp.rf.rf[22][1] ),
    .I3(\dp.rf.rf[23][1] ),
    .S0(net550),
    .S1(net14),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07435_ (.I0(_02835_),
    .I1(_02836_),
    .I2(_02837_),
    .I3(_02838_),
    .S0(_01066_),
    .S1(net17),
    .Z(_02839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07436_ (.A1(net15),
    .A2(_02839_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07437_ (.I0(\dp.rf.rf[2][1] ),
    .I1(\dp.rf.rf[3][1] ),
    .S(net550),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07438_ (.A1(_01036_),
    .A2(net16),
    .A3(_02841_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07439_ (.I0(\dp.rf.rf[0][1] ),
    .I1(\dp.rf.rf[1][1] ),
    .I2(\dp.rf.rf[8][1] ),
    .I3(\dp.rf.rf[9][1] ),
    .S0(net550),
    .S1(net16),
    .Z(_02843_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07440_ (.A1(net14),
    .A2(_02843_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07441_ (.I0(\dp.rf.rf[10][1] ),
    .I1(\dp.rf.rf[11][1] ),
    .S(net550),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07442_ (.A1(_02106_),
    .A2(_02845_),
    .B(_01055_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07443_ (.A1(_02254_),
    .A2(_02842_),
    .A3(_02844_),
    .A4(_02846_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07444_ (.I0(\dp.rf.rf[24][1] ),
    .I1(\dp.rf.rf[25][1] ),
    .S(net550),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07445_ (.A1(net14),
    .A2(_01066_),
    .A3(_02848_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07446_ (.I0(\dp.rf.rf[18][1] ),
    .I1(\dp.rf.rf[19][1] ),
    .S(net13),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07447_ (.A1(_01036_),
    .A2(net16),
    .A3(_02850_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07448_ (.I0(\dp.rf.rf[26][1] ),
    .I1(\dp.rf.rf[27][1] ),
    .S(net550),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07449_ (.I0(\dp.rf.rf[16][1] ),
    .I1(\dp.rf.rf[17][1] ),
    .S(net551),
    .Z(_02853_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07450_ (.A1(_02106_),
    .A2(_02852_),
    .B1(_02853_),
    .B2(_02109_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07451_ (.A1(_02105_),
    .A2(_02849_),
    .A3(_02851_),
    .A4(_02854_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07452_ (.A1(_02840_),
    .A2(_02847_),
    .A3(_02855_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07453_ (.I(_02856_),
    .ZN(net144));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07454_ (.A1(_01119_),
    .A2(_02830_),
    .A3(_02834_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07455_ (.A1(_01311_),
    .A2(_02856_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07456_ (.A1(_02857_),
    .A2(_02858_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_283_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_283_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_282_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_282_clk));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07459_ (.A1(_01110_),
    .A2(_02859_),
    .ZN(_05095_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07460_ (.I(_05095_[0]),
    .ZN(_05354_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07461_ (.I0(\dp.rf.rf[22][1] ),
    .I1(\dp.rf.rf[23][1] ),
    .S(net7),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07462_ (.I(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07463_ (.A1(net536),
    .A2(_02863_),
    .B(net523),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07464_ (.I(\dp.rf.rf[18][1] ),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07465_ (.A1(_02865_),
    .A2(net533),
    .A3(net532),
    .A4(_01125_),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07466_ (.I0(\dp.rf.rf[18][1] ),
    .I1(\dp.rf.rf[19][1] ),
    .S(net7),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07467_ (.I(_02867_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07468_ (.A1(net521),
    .A2(_02866_),
    .A3(_02868_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07469_ (.I0(\dp.rf.rf[17][1] ),
    .I1(\dp.rf.rf[21][1] ),
    .S(net536),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07470_ (.A1(_01148_),
    .A2(_02870_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07471_ (.A1(\dp.rf.rf[20][1] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07472_ (.A1(_02871_),
    .A2(_02872_),
    .B(_01144_),
    .C(net529),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07473_ (.I(\dp.rf.rf[16][1] ),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07474_ (.A1(_02874_),
    .A2(_01385_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07475_ (.A1(_02864_),
    .A2(_02869_),
    .B1(_02873_),
    .B2(_02875_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07476_ (.I0(\dp.rf.rf[24][1] ),
    .I1(\dp.rf.rf[25][1] ),
    .I2(\dp.rf.rf[28][1] ),
    .I3(\dp.rf.rf[29][1] ),
    .S0(net7),
    .S1(net535),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07477_ (.A1(_01140_),
    .A2(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07478_ (.I0(\dp.rf.rf[27][1] ),
    .I1(\dp.rf.rf[31][1] ),
    .S(net535),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07479_ (.I0(\dp.rf.rf[26][1] ),
    .I1(\dp.rf.rf[30][1] ),
    .S(net535),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07480_ (.A1(_01697_),
    .A2(_02879_),
    .B1(_02880_),
    .B2(_01702_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07481_ (.A1(_01580_),
    .A2(_02878_),
    .A3(_02881_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07482_ (.I0(\dp.rf.rf[8][1] ),
    .I1(\dp.rf.rf[9][1] ),
    .I2(\dp.rf.rf[12][1] ),
    .I3(\dp.rf.rf[13][1] ),
    .S0(net7),
    .S1(net9),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07483_ (.I0(\dp.rf.rf[1][1] ),
    .I1(\dp.rf.rf[5][1] ),
    .S(net9),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07484_ (.A1(_01148_),
    .A2(_02884_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07485_ (.A1(\dp.rf.rf[4][1] ),
    .A2(net7),
    .A3(_01167_),
    .B(_01140_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07486_ (.A1(_02885_),
    .A2(_02886_),
    .B(net529),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07487_ (.I0(\dp.rf.rf[10][1] ),
    .I1(\dp.rf.rf[11][1] ),
    .I2(\dp.rf.rf[14][1] ),
    .I3(\dp.rf.rf[15][1] ),
    .S0(net7),
    .S1(net9),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07488_ (.I0(\dp.rf.rf[2][1] ),
    .I1(\dp.rf.rf[3][1] ),
    .I2(\dp.rf.rf[6][1] ),
    .I3(\dp.rf.rf[7][1] ),
    .S0(net7),
    .S1(net9),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07489_ (.I0(_02888_),
    .I1(_02889_),
    .S(_01144_),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07490_ (.A1(_01279_),
    .A2(_02883_),
    .B1(_02887_),
    .B2(_01458_),
    .C1(_01781_),
    .C2(_02890_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _07491_ (.A1(_01475_),
    .A2(_02876_),
    .A3(_02882_),
    .B(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_281_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_281_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07493_ (.I(_02892_),
    .ZN(_05353_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07494_ (.A1(_01128_),
    .A2(_01130_),
    .A3(_01132_),
    .B(_02004_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07495_ (.I0(_01088_),
    .I1(_02893_),
    .S(_01119_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_280_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_280_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07497_ (.A1(_02857_),
    .A2(_02858_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_277_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_277_clk));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07499_ (.A1(net503),
    .A2(_01230_),
    .A3(net499),
    .Z(_02898_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07500_ (.A1(_01311_),
    .A2(net159),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07501_ (.A1(_01119_),
    .A2(_05373_[0]),
    .B(_02899_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_276_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_276_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07503_ (.A1(_01098_),
    .A2(_01092_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07504_ (.A1(_01089_),
    .A2(_02902_),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _07505_ (.A1(net6),
    .A2(net4),
    .A3(_02903_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07506_ (.A1(_02900_),
    .A2(_02904_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07507_ (.A1(_01311_),
    .A2(net158),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07508_ (.A1(_01119_),
    .A2(_05367_[0]),
    .B(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07509_ (.A1(_01119_),
    .A2(net155),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07510_ (.A1(_01311_),
    .A2(_05363_[0]),
    .B(_02908_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_271_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_271_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_270_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_270_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07513_ (.A1(_02907_),
    .A2(net496),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07514_ (.A1(_02905_),
    .A2(_02912_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07515_ (.A1(_01100_),
    .A2(net24),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _07516_ (.A1(net4),
    .A2(net528),
    .A3(_02903_),
    .A4(_02914_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_268_clk (.I(clknet_6_63__leaf_clk),
    .Z(clknet_leaf_268_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_267_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_267_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07519_ (.A1(_02898_),
    .A2(_02913_),
    .B(_02915_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07520_ (.A1(net6),
    .A2(net4),
    .A3(_02903_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_264_clk (.I(clknet_6_63__leaf_clk),
    .Z(clknet_leaf_264_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07522_ (.A1(_02900_),
    .A2(_02919_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07523_ (.I0(_02284_),
    .I1(_02382_),
    .S(net499),
    .Z(_02922_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_261_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_261_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_256_clk (.I(clknet_6_60__leaf_clk),
    .Z(clknet_leaf_256_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_254_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_254_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_253_clk (.I(clknet_6_60__leaf_clk),
    .Z(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07528_ (.I0(_02470_),
    .I1(net507),
    .S(net499),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_251_clk (.I(clknet_6_60__leaf_clk),
    .Z(clknet_leaf_251_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_250_clk (.I(clknet_6_60__leaf_clk),
    .Z(clknet_leaf_250_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07531_ (.I0(_02236_),
    .I1(_02327_),
    .S(net499),
    .Z(_02926_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_249_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_249_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_248_clk (.I(clknet_6_60__leaf_clk),
    .Z(clknet_leaf_248_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07534_ (.I0(_02428_),
    .I1(_02518_),
    .S(net499),
    .Z(_02927_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_246_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_246_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07536_ (.I0(_02922_),
    .I1(_02925_),
    .I2(_02926_),
    .I3(_02927_),
    .S0(net496),
    .S1(net509),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_244_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_243_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_242_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_242_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_238_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_238_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07541_ (.I0(_05303_[0]),
    .I1(_02645_),
    .I2(_02683_),
    .I3(net506),
    .S0(net503),
    .S1(net499),
    .Z(_02931_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_237_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_237_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07543_ (.I0(_01230_),
    .I1(_02828_),
    .S(net500),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_232_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_232_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07545_ (.I0(net501),
    .I1(_02892_),
    .S(net499),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07546_ (.I0(_02932_),
    .I1(_02933_),
    .S(net509),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_231_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07548_ (.I0(_02931_),
    .I1(_02934_),
    .S(net496),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_230_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_228_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_228_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07551_ (.I0(_02929_),
    .I1(_02936_),
    .S(_02907_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_224_clk (.I(clknet_6_39__leaf_clk),
    .Z(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07553_ (.A1(_02704_),
    .A2(_02919_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_223_clk (.I(clknet_6_39__leaf_clk),
    .Z(clknet_leaf_223_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_222_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_222_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_221_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_220_clk (.I(clknet_6_39__leaf_clk),
    .Z(clknet_leaf_220_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07558_ (.I0(_01899_),
    .I1(_01997_),
    .I2(_02086_),
    .I3(net508),
    .S0(_02896_),
    .S1(_02909_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_216_clk (.I(clknet_6_39__leaf_clk),
    .Z(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_215_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07561_ (.I0(_01852_),
    .I1(_01947_),
    .I2(_02044_),
    .I3(_02142_),
    .S0(_02896_),
    .S1(_02909_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07562_ (.I0(_02944_),
    .I1(_02945_),
    .S(net509),
    .Z(_02946_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_211_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_208_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_208_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_205_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_205_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07566_ (.I0(_01287_),
    .I1(_01414_),
    .I2(_05127_[0]),
    .I3(_05135_[0]),
    .S0(_02894_),
    .S1(_02896_),
    .Z(_02948_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_200_clk (.I(clknet_6_32__leaf_clk),
    .Z(clknet_leaf_200_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_198_clk (.I(clknet_6_33__leaf_clk),
    .Z(clknet_leaf_198_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07569_ (.I0(_01602_),
    .I1(_01657_),
    .I2(_05159_[0]),
    .I3(_01786_),
    .S0(_02894_),
    .S1(_02896_),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07570_ (.I0(_02948_),
    .I1(_02951_),
    .S(_02909_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_195_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_195_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07572_ (.I0(_02946_),
    .I1(_02952_),
    .S(net505),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07573_ (.A1(_02921_),
    .A2(_02939_),
    .B1(_02941_),
    .B2(_02954_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07574_ (.A1(_01241_),
    .A2(_01286_),
    .A3(_01312_),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07575_ (.A1(_01241_),
    .A2(_01286_),
    .B(_01312_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07576_ (.A1(net27),
    .A2(_01094_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07577_ (.A1(_01092_),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07578_ (.A1(_01100_),
    .A2(net4),
    .A3(net5),
    .A4(_02959_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07579_ (.A1(_02956_),
    .A2(_02957_),
    .B(_02960_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _07580_ (.A1(net511),
    .A2(_02961_),
    .Z(_02962_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07581_ (.A1(net5),
    .A2(_02902_),
    .B(net4),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07582_ (.A1(_02959_),
    .A2(_02963_),
    .B(_01100_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07583_ (.A1(net6),
    .A2(net4),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07584_ (.A1(_02902_),
    .A2(_02965_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07585_ (.A1(_01089_),
    .A2(_02966_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07586_ (.A1(_01108_),
    .A2(_02964_),
    .A3(_02967_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_194_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_194_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_193_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07589_ (.A1(_01108_),
    .A2(_02959_),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07590_ (.A1(net5),
    .A2(_02965_),
    .Z(_02972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07591_ (.A1(_02971_),
    .A2(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_192_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_192_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07593_ (.A1(_02968_),
    .A2(_02973_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07594_ (.A1(_05114_[0]),
    .A2(_02962_),
    .A3(_02975_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07595_ (.A1(_02968_),
    .A2(_02973_),
    .Z(_02977_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07596_ (.A1(_05113_[0]),
    .A2(_05121_[0]),
    .A3(_02962_),
    .A4(_02977_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07597_ (.I(_05338_[0]),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07598_ (.A1(_05096_[0]),
    .A2(_05346_[0]),
    .B(_05345_[0]),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07599_ (.I(_05337_[0]),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07600_ (.A1(_02979_),
    .A2(_02980_),
    .B(_02981_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _07601_ (.A1(_05313_[0]),
    .A2(_05329_[0]),
    .A3(_05321_[0]),
    .Z(_02983_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07602_ (.A1(_05330_[0]),
    .A2(_02982_),
    .B(_02983_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07603_ (.A1(_05290_[0]),
    .A2(_05298_[0]),
    .A3(_05306_[0]),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07604_ (.I(_05313_[0]),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07605_ (.A1(_05322_[0]),
    .A2(_05321_[0]),
    .B(_05314_[0]),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07606_ (.A1(_02986_),
    .A2(_02987_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07607_ (.A1(_05274_[0]),
    .A2(_05282_[0]),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07608_ (.A1(_02985_),
    .A2(_02988_),
    .A3(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07609_ (.I(_05290_[0]),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07610_ (.A1(_05298_[0]),
    .A2(_05305_[0]),
    .B(_05297_[0]),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07611_ (.I(_05289_[0]),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07612_ (.A1(_02991_),
    .A2(_02992_),
    .B(_02993_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07613_ (.A1(_05281_[0]),
    .A2(_05274_[0]),
    .B1(_02994_),
    .B2(_02989_),
    .C(_05273_[0]),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07614_ (.I(_05265_[0]),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _07615_ (.I(_05257_[0]),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07616_ (.I(_05225_[0]),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07617_ (.I(_05241_[0]),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07618_ (.A1(_05233_[0]),
    .A2(_05226_[0]),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07619_ (.A1(_05249_[0]),
    .A2(_05242_[0]),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _07620_ (.A1(_02998_),
    .A2(_02999_),
    .A3(_03000_),
    .A4(_03001_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07621_ (.A1(_02996_),
    .A2(_02997_),
    .A3(_03002_),
    .Z(_03003_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07622_ (.A1(_02984_),
    .A2(_02990_),
    .B(_02995_),
    .C(_03003_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _07623_ (.I(_05258_[0]),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07624_ (.A1(_05265_[0]),
    .A2(_05266_[0]),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07625_ (.A1(_03005_),
    .A2(_03006_),
    .B(_03002_),
    .C(_02997_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07626_ (.A1(_05249_[0]),
    .A2(_05250_[0]),
    .B(_05242_[0]),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07627_ (.I(_05234_[0]),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07628_ (.A1(_02999_),
    .A2(_03008_),
    .B(_03009_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07629_ (.A1(_05233_[0]),
    .A2(_03010_),
    .B(_05226_[0]),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07630_ (.A1(_02998_),
    .A2(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07631_ (.A1(_05186_[0]),
    .A2(_05194_[0]),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07632_ (.A1(_05218_[0]),
    .A2(_05202_[0]),
    .A3(_05210_[0]),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07633_ (.A1(_03013_),
    .A2(_03014_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _07634_ (.A1(_03004_),
    .A2(_03007_),
    .A3(_03012_),
    .A4(_03015_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07635_ (.A1(_05186_[0]),
    .A2(_05193_[0]),
    .B(_05185_[0]),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07636_ (.A1(_05186_[0]),
    .A2(_05194_[0]),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07637_ (.I(_05209_[0]),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07638_ (.A1(_05217_[0]),
    .A2(_05210_[0]),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07639_ (.A1(_03019_),
    .A2(_03020_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07640_ (.A1(_05202_[0]),
    .A2(_03021_),
    .B(_05201_[0]),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07641_ (.A1(_03018_),
    .A2(_03022_),
    .Z(_03023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07642_ (.A1(_03017_),
    .A2(_03023_),
    .Z(_03024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07643_ (.A1(_05170_[0]),
    .A2(_05178_[0]),
    .Z(_03025_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07644_ (.A1(_05162_[0]),
    .A2(_03025_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07645_ (.A1(_03016_),
    .A2(_03024_),
    .B(_03026_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07646_ (.I(_05162_[0]),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07647_ (.A1(_05170_[0]),
    .A2(_05177_[0]),
    .B(_05169_[0]),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07648_ (.A1(_03028_),
    .A2(_03029_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07649_ (.A1(_05145_[0]),
    .A2(_05153_[0]),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _07650_ (.A1(_05161_[0]),
    .A2(_03027_),
    .A3(_03030_),
    .A4(_03031_),
    .Z(_03032_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07651_ (.A1(_05154_[0]),
    .A2(_05145_[0]),
    .A3(_05153_[0]),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07652_ (.A1(_05146_[0]),
    .A2(_05145_[0]),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _07653_ (.A1(_03032_),
    .A2(_03033_),
    .A3(_03034_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07654_ (.A1(_05130_[0]),
    .A2(_05138_[0]),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07655_ (.A1(_05130_[0]),
    .A2(_05137_[0]),
    .B(_05129_[0]),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07656_ (.A1(_03035_),
    .A2(_03036_),
    .B(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07657_ (.A1(_05122_[0]),
    .A2(_03038_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07658_ (.I0(_02976_),
    .I1(_02978_),
    .S(_03039_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_190_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_189_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_189_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_187_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_187_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07662_ (.A1(net6),
    .A2(_01095_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07663_ (.A1(net5),
    .A2(_03044_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _07664_ (.A1(_02972_),
    .A2(_03045_),
    .B(_01108_),
    .C(_02959_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_185_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_185_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07666_ (.A1(_05105_[0]),
    .A2(net512),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07667_ (.A1(_05109_[0]),
    .A2(_02973_),
    .B(_03048_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07668_ (.A1(_02968_),
    .A2(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07669_ (.A1(_02971_),
    .A2(_02972_),
    .Z(_03051_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07670_ (.A1(_02968_),
    .A2(_03051_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07671_ (.A1(_01110_),
    .A2(_03052_),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07672_ (.A1(_02968_),
    .A2(_03051_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07673_ (.A1(_02971_),
    .A2(_03045_),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07674_ (.A1(_01110_),
    .A2(_03054_),
    .B(_03055_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07675_ (.I0(_03053_),
    .I1(_03056_),
    .S(_05106_[0]),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07676_ (.A1(_05114_[0]),
    .A2(_05113_[0]),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07677_ (.A1(_05114_[0]),
    .A2(_05121_[0]),
    .B(_05113_[0]),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07678_ (.I0(_03058_),
    .I1(_03059_),
    .S(_02962_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07679_ (.A1(_02977_),
    .A2(_03060_),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _07680_ (.A1(_02915_),
    .A2(_03050_),
    .A3(_03057_),
    .A4(_03061_),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07681_ (.A1(_02918_),
    .A2(_02955_),
    .B1(_03040_),
    .B2(_03062_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07682_ (.A1(net28),
    .A2(_02902_),
    .Z(_03063_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _07683_ (.I(_03063_),
    .ZN(net98));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_179_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_179_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_177_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_176_clk (.I(clknet_6_51__leaf_clk),
    .Z(clknet_leaf_176_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_175_clk (.I(clknet_6_50__leaf_clk),
    .Z(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07688_ (.A1(_05097_[0]),
    .A2(_03054_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_174_clk (.I(clknet_6_50__leaf_clk),
    .Z(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_173_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07691_ (.A1(_05351_[0]),
    .A2(net512),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07692_ (.A1(_05355_[0]),
    .A2(_02973_),
    .B(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _07693_ (.A1(net4),
    .A2(net528),
    .A3(_02903_),
    .A4(_02914_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07694_ (.A1(_05352_[0]),
    .A2(_03055_),
    .B1(_03072_),
    .B2(_02968_),
    .C(_03073_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07695_ (.A1(_03068_),
    .A2(_03074_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_172_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_172_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07697_ (.A1(net502),
    .A2(_02919_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07698_ (.I0(_01786_),
    .I1(_01899_),
    .S(_02896_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07699_ (.I0(_01997_),
    .I1(_02086_),
    .S(_02896_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07700_ (.I0(_03078_),
    .I1(_03079_),
    .S(_02909_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_171_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_171_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07702_ (.I0(_02945_),
    .I1(_03080_),
    .S(net509),
    .Z(_03082_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07703_ (.A1(net505),
    .A2(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _07704_ (.I(net24),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07705_ (.I0(_01288_),
    .I1(_05131_[0]),
    .S(_02896_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07706_ (.A1(_01414_),
    .A2(_02896_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07707_ (.I0(_03085_),
    .I1(_03086_),
    .S(net509),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07708_ (.I0(_05139_[0]),
    .I1(_05147_[0]),
    .I2(_05155_[0]),
    .I3(_05163_[0]),
    .S0(_02894_),
    .S1(_02896_),
    .Z(_03088_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07709_ (.A1(_02909_),
    .A2(_03088_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07710_ (.A1(net504),
    .A2(_03087_),
    .B(_03089_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_170_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_170_clk));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07712_ (.A1(net509),
    .A2(_01461_),
    .A3(_01480_),
    .Z(_03092_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07713_ (.A1(net503),
    .A2(_01414_),
    .B(_02896_),
    .C(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07714_ (.A1(_01287_),
    .A2(net500),
    .B(_02909_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07715_ (.A1(_02909_),
    .A2(_03088_),
    .B1(_03093_),
    .B2(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07716_ (.A1(net24),
    .A2(_03095_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_165_clk (.I(clknet_6_33__leaf_clk),
    .Z(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_163_clk (.I(clknet_6_33__leaf_clk),
    .Z(clknet_leaf_163_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07719_ (.A1(_03084_),
    .A2(_03090_),
    .B(_03096_),
    .C(_02907_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07720_ (.I0(_02382_),
    .I1(_02428_),
    .I2(_02470_),
    .I3(_02518_),
    .S0(net503),
    .S1(net499),
    .Z(_03100_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_162_clk (.I(clknet_6_50__leaf_clk),
    .Z(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07722_ (.I0(net508),
    .I1(_02236_),
    .I2(_02284_),
    .I3(_02327_),
    .S0(net503),
    .S1(net499),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07723_ (.I0(_03100_),
    .I1(_03101_),
    .S(net504),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07724_ (.I0(net507),
    .I1(_05303_[0]),
    .I2(_02645_),
    .I3(_02683_),
    .S0(net503),
    .S1(net499),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07725_ (.I0(net506),
    .I1(net501),
    .I2(_02828_),
    .I3(_02892_),
    .S0(net503),
    .S1(net499),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07726_ (.I0(_03103_),
    .I1(_03104_),
    .S(net496),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07727_ (.I0(_03102_),
    .I1(_03105_),
    .S(net497),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07728_ (.I0(_01230_),
    .I1(_02892_),
    .S(net503),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07729_ (.A1(net499),
    .A2(_03107_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07730_ (.A1(_02921_),
    .A2(_03106_),
    .B1(_03108_),
    .B2(_02913_),
    .C(net510),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07731_ (.A1(_03077_),
    .A2(_03083_),
    .A3(_03099_),
    .B(_03109_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07732_ (.A1(_03075_),
    .A2(_03110_),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_161_clk (.I(clknet_6_50__leaf_clk),
    .Z(clknet_leaf_161_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07734_ (.A1(_02968_),
    .A2(_03051_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07735_ (.I(_05349_[0]),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_160_clk (.I(clknet_6_50__leaf_clk),
    .Z(clknet_leaf_160_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_153_clk (.I(clknet_6_32__leaf_clk),
    .Z(clknet_leaf_153_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07738_ (.A1(_05346_[0]),
    .A2(_03055_),
    .B1(_03112_),
    .B2(_03113_),
    .C(_03073_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_150_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _07740_ (.A1(_05096_[0]),
    .A2(_05346_[0]),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07741_ (.I0(_03118_),
    .I1(_05345_[0]),
    .S(_02968_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07742_ (.A1(net512),
    .A2(_03119_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07743_ (.I0(_05127_[0]),
    .I1(_05135_[0]),
    .I2(_01602_),
    .I3(_01657_),
    .S0(_02894_),
    .S1(_02896_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07744_ (.I0(_01287_),
    .I1(_01414_),
    .S(_02894_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07745_ (.A1(net504),
    .A2(_02896_),
    .A3(_03122_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07746_ (.A1(_02909_),
    .A2(_03121_),
    .B(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07747_ (.I0(_05171_[0]),
    .I1(_05187_[0]),
    .S(_02896_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07748_ (.I0(_05203_[0]),
    .I1(_05219_[0]),
    .S(_02896_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07749_ (.I0(_05163_[0]),
    .I1(_05179_[0]),
    .S(_02896_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07750_ (.I0(_05195_[0]),
    .I1(_05211_[0]),
    .S(_02896_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07751_ (.I0(_03125_),
    .I1(_03126_),
    .I2(_03127_),
    .I3(_03128_),
    .S0(_02909_),
    .S1(net509),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07752_ (.A1(_02907_),
    .A2(_03129_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07753_ (.A1(_03084_),
    .A2(_02919_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07754_ (.A1(net505),
    .A2(_03124_),
    .B(_03130_),
    .C(_03131_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07755_ (.A1(_02894_),
    .A2(_02896_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07756_ (.A1(_02894_),
    .A2(_05123_[0]),
    .A3(_02896_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07757_ (.A1(_01288_),
    .A2(_03133_),
    .B(_03134_),
    .C(_02909_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07758_ (.A1(_02909_),
    .A2(_03121_),
    .B(_03135_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07759_ (.A1(net24),
    .A2(_02919_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07760_ (.A1(net505),
    .A2(_03136_),
    .B(_03130_),
    .C(_03137_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _07761_ (.A1(_03132_),
    .A2(_03138_),
    .B(net502),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07762_ (.I0(net508),
    .I1(_02284_),
    .S(_02896_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07763_ (.I0(_02142_),
    .I1(_02236_),
    .S(_02896_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07764_ (.I0(_03140_),
    .I1(_03141_),
    .S(net509),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07765_ (.I0(_02327_),
    .I1(_02382_),
    .I2(_02428_),
    .I3(_02470_),
    .S0(net503),
    .S1(_02896_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07766_ (.I0(_03142_),
    .I1(_03143_),
    .S(net496),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07767_ (.I0(_02518_),
    .I1(net507),
    .I2(_05303_[0]),
    .I3(_02645_),
    .S0(net503),
    .S1(_02896_),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07768_ (.I0(_02683_),
    .I1(net506),
    .I2(net501),
    .I3(_02828_),
    .S0(net503),
    .S1(net499),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07769_ (.I0(_03145_),
    .I1(_03146_),
    .S(net496),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07770_ (.I0(_03144_),
    .I1(_03147_),
    .S(_02907_),
    .Z(_03148_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07771_ (.A1(net499),
    .A2(_02892_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07772_ (.I0(_01230_),
    .I1(_02828_),
    .S(net499),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07773_ (.I0(_03149_),
    .I1(_03150_),
    .S(net503),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07774_ (.A1(_02921_),
    .A2(_03148_),
    .B1(_03151_),
    .B2(_02913_),
    .C(_02915_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _07775_ (.A1(_03116_),
    .A2(_03120_),
    .B1(_03139_),
    .B2(_03152_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07776_ (.A1(_01088_),
    .A2(_01119_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07777_ (.A1(_01128_),
    .A2(_01130_),
    .A3(_01132_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07778_ (.A1(net533),
    .A2(_01118_),
    .A3(_01135_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07779_ (.A1(_01099_),
    .A2(_01109_),
    .B1(_03154_),
    .B2(_03155_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07780_ (.A1(_03153_),
    .A2(_03156_),
    .B1(_05107_[0]),
    .B2(_01137_),
    .ZN(_05093_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07781_ (.I0(_05123_[0]),
    .I1(_05131_[0]),
    .I2(_05139_[0]),
    .I3(_05147_[0]),
    .S0(_02894_),
    .S1(_02896_),
    .Z(_03157_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07782_ (.A1(net496),
    .A2(_03157_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07783_ (.A1(_01288_),
    .A2(net504),
    .B(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _07784_ (.A1(net509),
    .A2(_01288_),
    .A3(net500),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07785_ (.A1(net504),
    .A2(_03160_),
    .B(_03158_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07786_ (.I0(_03159_),
    .I1(_03161_),
    .S(_03084_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07787_ (.I0(_03127_),
    .I1(_03128_),
    .S(_02909_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07788_ (.I0(_05187_[0]),
    .I1(_05203_[0]),
    .S(_02896_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07789_ (.I0(_05155_[0]),
    .I1(_05171_[0]),
    .S(_02896_),
    .Z(_03165_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_145_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_145_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07791_ (.I0(_03164_),
    .I1(_03165_),
    .S(net504),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07792_ (.I0(_03163_),
    .I1(_03167_),
    .S(net509),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07793_ (.A1(net505),
    .A2(_03168_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07794_ (.A1(net505),
    .A2(_03162_),
    .B(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07795_ (.I0(_05219_[0]),
    .I1(_05235_[0]),
    .I2(_05251_[0]),
    .I3(_05267_[0]),
    .S0(_02896_),
    .S1(net496),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07796_ (.I0(_05227_[0]),
    .I1(_05243_[0]),
    .I2(_05259_[0]),
    .I3(_05275_[0]),
    .S0(_02896_),
    .S1(net496),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_143_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_143_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07798_ (.I0(_03171_),
    .I1(_03172_),
    .S(net503),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07799_ (.I0(_02470_),
    .I1(_02518_),
    .I2(net507),
    .I3(_05303_[0]),
    .S0(net503),
    .S1(net499),
    .Z(_03175_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07800_ (.I0(_02645_),
    .I1(_02683_),
    .I2(net506),
    .I3(net501),
    .S0(net503),
    .S1(net499),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07801_ (.I0(_03175_),
    .I1(_03176_),
    .S(net496),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07802_ (.A1(net497),
    .A2(_03177_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07803_ (.A1(net497),
    .A2(_03174_),
    .B(_03178_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_141_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_141_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07805_ (.I0(net501),
    .I1(_02892_),
    .S(net500),
    .Z(_03181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07806_ (.I0(_03150_),
    .I1(_03181_),
    .S(net503),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07807_ (.A1(_02921_),
    .A2(_03179_),
    .B1(_03182_),
    .B2(_02913_),
    .C(_02915_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07808_ (.A1(_03077_),
    .A2(_03170_),
    .B(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07809_ (.A1(_01088_),
    .A2(_01119_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _07810_ (.A1(net29),
    .A2(net533),
    .A3(_01032_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07811_ (.A1(net4),
    .A2(net5),
    .A3(_01094_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07812_ (.A1(net5),
    .A2(_01094_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07813_ (.A1(_03186_),
    .A2(_03187_),
    .B(_03188_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07814_ (.A1(net5),
    .A2(_03186_),
    .B1(_03189_),
    .B2(net27),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07815_ (.A1(_01100_),
    .A2(_01108_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _07816_ (.A1(_03190_),
    .A2(_03191_),
    .B1(_01311_),
    .B2(_02893_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07817_ (.A1(_05352_[0]),
    .A2(_05346_[0]),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _07818_ (.A1(_03185_),
    .A2(_03192_),
    .B1(_01230_),
    .B2(_02894_),
    .C(_03193_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07819_ (.A1(_05351_[0]),
    .A2(_05346_[0]),
    .B(_05345_[0]),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07820_ (.A1(_03194_),
    .A2(_03195_),
    .Z(_03196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07821_ (.A1(_03054_),
    .A2(_03196_),
    .B(_03055_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_139_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_137_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_137_clk));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07824_ (.A1(_05338_[0]),
    .A2(_03052_),
    .A3(_03196_),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_136_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_134_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_134_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07827_ (.A1(_05337_[0]),
    .A2(net512),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07828_ (.A1(_05341_[0]),
    .A2(_02973_),
    .B(_03203_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07829_ (.A1(_02968_),
    .A2(_03204_),
    .B(_03073_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07830_ (.A1(_02979_),
    .A2(_03197_),
    .B(_03200_),
    .C(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07831_ (.A1(_03184_),
    .A2(_03206_),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07832_ (.A1(net505),
    .A2(_02951_),
    .B(net504),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07833_ (.I0(_05179_[0]),
    .I1(_05195_[0]),
    .S(_02896_),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07834_ (.I0(_05147_[0]),
    .I1(_05163_[0]),
    .S(_02896_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07835_ (.I0(_03164_),
    .I1(_03208_),
    .I2(_03165_),
    .I3(_03209_),
    .S0(net509),
    .S1(net504),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07836_ (.A1(net496),
    .A2(_02948_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07837_ (.I0(_03210_),
    .I1(_03211_),
    .S(net505),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07838_ (.A1(_03084_),
    .A2(_01288_),
    .A3(_03207_),
    .B(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07839_ (.I0(_02428_),
    .I1(_02470_),
    .I2(_02518_),
    .I3(net507),
    .S0(net503),
    .S1(net499),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07840_ (.I0(_02931_),
    .I1(_03214_),
    .S(net504),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07841_ (.I0(net506),
    .I1(net501),
    .I2(_02828_),
    .I3(_02892_),
    .S0(net509),
    .S1(net500),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07842_ (.I0(_02898_),
    .I1(_03216_),
    .S(net496),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07843_ (.I0(_03215_),
    .I1(_03217_),
    .S(_02904_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07844_ (.I0(_02086_),
    .I1(net508),
    .I2(_02284_),
    .I3(_02382_),
    .S0(_02896_),
    .S1(net496),
    .Z(_03219_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07845_ (.I0(_02044_),
    .I1(_02142_),
    .I2(_02236_),
    .I3(_02327_),
    .S0(_02896_),
    .S1(net496),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07846_ (.I0(_03219_),
    .I1(_03220_),
    .S(net509),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07847_ (.A1(_02919_),
    .A2(_03221_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07848_ (.I0(_03218_),
    .I1(_03222_),
    .S(net505),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_131_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_131_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07850_ (.A1(_02941_),
    .A2(_03213_),
    .B1(_03223_),
    .B2(_02900_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _07851_ (.A1(_05330_[0]),
    .A2(_02982_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07852_ (.I0(_03226_),
    .I1(_05329_[0]),
    .S(_02968_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07853_ (.I(_05333_[0]),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07854_ (.A1(_05330_[0]),
    .A2(_03055_),
    .B1(net512),
    .B2(_03227_),
    .C1(_03112_),
    .C2(_03228_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07855_ (.I0(_03225_),
    .I1(_03229_),
    .S(_02915_),
    .Z(_03230_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07856_ (.I(_03230_),
    .ZN(net92));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07857_ (.I0(_01414_),
    .I1(_05127_[0]),
    .S(_02894_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07858_ (.A1(_02909_),
    .A2(_02896_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07859_ (.A1(_02909_),
    .A2(_02896_),
    .B(_01288_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07860_ (.A1(_03231_),
    .A2(_03232_),
    .B(_03233_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _07861_ (.A1(net504),
    .A2(_03087_),
    .A3(_03131_),
    .B1(_03137_),
    .B2(_03234_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07862_ (.I0(_05139_[0]),
    .I1(_05155_[0]),
    .S(_02896_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07863_ (.I0(_03208_),
    .I1(_03209_),
    .I2(_03125_),
    .I3(_03236_),
    .S0(net504),
    .S1(net509),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07864_ (.A1(net505),
    .A2(_02904_),
    .A3(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07865_ (.A1(net505),
    .A2(_03235_),
    .B(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_127_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_126_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07868_ (.I0(_02683_),
    .I1(net506),
    .I2(net501),
    .I3(_02828_),
    .S0(net509),
    .S1(net500),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07869_ (.I0(_03108_),
    .I1(_03242_),
    .S(net496),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07870_ (.I0(_03100_),
    .I1(_03103_),
    .S(net496),
    .Z(_03244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07871_ (.I0(_03243_),
    .I1(_03244_),
    .S(_02919_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07872_ (.I0(_01997_),
    .I1(_02086_),
    .I2(net508),
    .I3(_02284_),
    .S0(_02896_),
    .S1(net496),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07873_ (.I0(_03220_),
    .I1(_03246_),
    .S(net509),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07874_ (.A1(net505),
    .A2(_02919_),
    .A3(_03247_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07875_ (.A1(net497),
    .A2(_03245_),
    .B(_03248_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07876_ (.I0(_03239_),
    .I1(_03249_),
    .S(_02900_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07877_ (.A1(_05337_[0]),
    .A2(_05330_[0]),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07878_ (.A1(_05329_[0]),
    .A2(_03251_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07879_ (.A1(_05345_[0]),
    .A2(_05351_[0]),
    .A3(_03252_),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07880_ (.A1(_05352_[0]),
    .A2(_05093_[0]),
    .B(_03253_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07881_ (.A1(_05330_[0]),
    .A2(_05338_[0]),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07882_ (.A1(_05345_[0]),
    .A2(_05346_[0]),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07883_ (.A1(_03255_),
    .A2(_03256_),
    .B(_03252_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07884_ (.A1(_03254_),
    .A2(_03257_),
    .Z(_03258_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07885_ (.A1(_05322_[0]),
    .A2(_03258_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07886_ (.A1(_05321_[0]),
    .A2(net512),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07887_ (.A1(_05325_[0]),
    .A2(_02973_),
    .B(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _07888_ (.A1(_05322_[0]),
    .A2(_03055_),
    .B1(_03054_),
    .B2(_03259_),
    .C1(_03261_),
    .C2(_02968_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07889_ (.I0(_03250_),
    .I1(_03262_),
    .S(_02915_),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07890_ (.I(_03263_),
    .ZN(net93));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07891_ (.A1(_02896_),
    .A2(_02892_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07892_ (.I0(_05107_[0]),
    .I1(_05347_[0]),
    .S(_02896_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07893_ (.I0(_05323_[0]),
    .I1(_05339_[0]),
    .S(net500),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07894_ (.I0(_05315_[0]),
    .I1(_05331_[0]),
    .S(net500),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07895_ (.I0(_03264_),
    .I1(_03265_),
    .I2(_03266_),
    .I3(_03267_),
    .S0(_02894_),
    .S1(_02909_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07896_ (.A1(_02919_),
    .A2(_03268_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07897_ (.I0(_03143_),
    .I1(_03145_),
    .S(net496),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07898_ (.A1(_02919_),
    .A2(_03270_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07899_ (.A1(_03269_),
    .A2(_03271_),
    .B(net505),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07900_ (.I0(_01947_),
    .I1(_02044_),
    .S(_02896_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _07901_ (.I0(_03079_),
    .I1(_03140_),
    .I2(_03273_),
    .I3(_03141_),
    .S0(net496),
    .S1(net509),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _07902_ (.A1(net505),
    .A2(_02919_),
    .A3(_03274_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_125_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07904_ (.A1(_03272_),
    .A2(_03275_),
    .B(_02900_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07905_ (.A1(_03122_),
    .A2(_03232_),
    .B(_02907_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07906_ (.A1(net24),
    .A2(_03233_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07907_ (.I0(_05159_[0]),
    .I1(_01786_),
    .I2(_01852_),
    .I3(_01899_),
    .S0(_02894_),
    .S1(_02896_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07908_ (.I0(_03280_),
    .I1(_03121_),
    .S(net504),
    .Z(_03281_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07909_ (.A1(net505),
    .A2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _07910_ (.A1(_03278_),
    .A2(_03279_),
    .B(_03077_),
    .C(_03282_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _07911_ (.A1(net510),
    .A2(_03283_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07912_ (.A1(_05313_[0]),
    .A2(net512),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07913_ (.A1(_05317_[0]),
    .A2(_02973_),
    .B(_03285_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07914_ (.A1(_02968_),
    .A2(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07915_ (.A1(_05330_[0]),
    .A2(_02982_),
    .Z(_03288_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _07916_ (.A1(_05329_[0]),
    .A2(_03288_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07917_ (.A1(_05322_[0]),
    .A2(_03289_),
    .B(_05321_[0]),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07918_ (.A1(_03290_),
    .A2(_03054_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07919_ (.A1(_03055_),
    .A2(_03291_),
    .B(_05314_[0]),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_121_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _07921_ (.A1(_05314_[0]),
    .A2(_03290_),
    .A3(_03052_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _07922_ (.A1(_02915_),
    .A2(_03287_),
    .A3(_03292_),
    .A4(_03294_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _07923_ (.A1(_03277_),
    .A2(_03284_),
    .B(_03295_),
    .ZN(net94));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07924_ (.A1(_05305_[0]),
    .A2(net512),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07925_ (.A1(_05309_[0]),
    .A2(_02973_),
    .B(_03296_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07926_ (.A1(_05314_[0]),
    .A2(_05322_[0]),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07927_ (.A1(_05314_[0]),
    .A2(_05321_[0]),
    .B(_05313_[0]),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07928_ (.A1(_03254_),
    .A2(_03257_),
    .A3(_03298_),
    .B(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07929_ (.A1(_03054_),
    .A2(_03300_),
    .Z(_03301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07930_ (.A1(_02971_),
    .A2(_03045_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07931_ (.A1(_03052_),
    .A2(_03300_),
    .B(_03302_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07932_ (.I0(_03301_),
    .I1(_03303_),
    .S(_05306_[0]),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07933_ (.A1(_02968_),
    .A2(_03297_),
    .B(_03304_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07934_ (.I0(_02327_),
    .I1(_02428_),
    .S(net499),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07935_ (.I0(_02922_),
    .I1(_03306_),
    .S(net503),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07936_ (.I0(_03175_),
    .I1(_03307_),
    .S(net504),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07937_ (.I0(_05303_[0]),
    .I1(_02683_),
    .I2(net501),
    .I3(_02892_),
    .S0(net500),
    .S1(net504),
    .Z(_03309_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07938_ (.I0(_01230_),
    .I1(net506),
    .I2(_02828_),
    .I3(_02645_),
    .S0(_02909_),
    .S1(_02896_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07939_ (.I0(_03309_),
    .I1(_03310_),
    .S(net509),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_118_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07941_ (.I0(_03308_),
    .I1(_03311_),
    .S(_02904_),
    .Z(_03313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07942_ (.I0(_03273_),
    .I1(_03141_),
    .S(net496),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07943_ (.I0(_02944_),
    .I1(_03314_),
    .S(net503),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07944_ (.A1(_02919_),
    .A2(_03315_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07945_ (.I0(_03313_),
    .I1(_03316_),
    .S(net505),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07946_ (.I0(_05155_[0]),
    .I1(_05163_[0]),
    .I2(_05171_[0]),
    .I3(_05179_[0]),
    .S0(_02894_),
    .S1(_02896_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07947_ (.I0(_03157_),
    .I1(_03318_),
    .S(_02909_),
    .Z(_03319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07948_ (.A1(_02907_),
    .A2(_03319_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07949_ (.A1(net504),
    .A2(_03133_),
    .B(_03084_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07950_ (.A1(_01287_),
    .A2(_03321_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07951_ (.A1(net505),
    .A2(_03322_),
    .B(_03077_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _07952_ (.A1(_02900_),
    .A2(_03317_),
    .B1(_03320_),
    .B2(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07953_ (.I0(_03305_),
    .I1(_03324_),
    .S(_03073_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07954_ (.I(_03325_),
    .ZN(net95));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07955_ (.I0(net507),
    .I1(_02645_),
    .I2(net506),
    .I3(_02828_),
    .S0(net500),
    .S1(net504),
    .Z(_03326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07956_ (.I0(_03309_),
    .I1(_03326_),
    .S(net503),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07957_ (.A1(net496),
    .A2(_02898_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07958_ (.I0(_02929_),
    .I1(_02946_),
    .I2(_03327_),
    .I3(_03328_),
    .S0(net505),
    .S1(_02904_),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07959_ (.A1(_03084_),
    .A2(_02919_),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07960_ (.A1(_02907_),
    .A2(_03330_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07961_ (.A1(net24),
    .A2(_02919_),
    .Z(_03332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07962_ (.A1(_01288_),
    .A2(net505),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _07963_ (.A1(_03332_),
    .A2(_03333_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07964_ (.A1(net505),
    .A2(_02952_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07965_ (.A1(_03331_),
    .A2(_03334_),
    .B(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07966_ (.I0(_03329_),
    .I1(_03336_),
    .S(_02704_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07967_ (.A1(_05297_[0]),
    .A2(net512),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07968_ (.A1(_05301_[0]),
    .A2(_02973_),
    .B(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _07969_ (.A1(_03288_),
    .A2(_02983_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07970_ (.A1(_05306_[0]),
    .A2(_03340_),
    .A3(_02988_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _07971_ (.A1(_05305_[0]),
    .A2(_03052_),
    .A3(_03341_),
    .B(_03302_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07972_ (.A1(_05305_[0]),
    .A2(_03341_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _07973_ (.A1(_05298_[0]),
    .A2(_03052_),
    .A3(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07974_ (.A1(_02968_),
    .A2(_03339_),
    .B1(_03342_),
    .B2(_05298_[0]),
    .C(_03344_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07975_ (.I(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_117_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07977_ (.I0(_03337_),
    .I1(_03346_),
    .S(_02915_),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07978_ (.A1(net496),
    .A2(_03108_),
    .Z(_03348_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07979_ (.I0(_02518_),
    .I1(_05303_[0]),
    .I2(_02683_),
    .I3(net501),
    .S0(net500),
    .S1(net504),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07980_ (.I0(_03326_),
    .I1(_03349_),
    .S(net503),
    .Z(_03350_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _07981_ (.I0(_03082_),
    .I1(_03102_),
    .I2(_03348_),
    .I3(_03350_),
    .S0(net497),
    .S1(_02904_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _07982_ (.A1(net504),
    .A2(_03087_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _07983_ (.A1(net505),
    .A2(_03095_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _07984_ (.A1(_03089_),
    .A2(_03352_),
    .A3(_03331_),
    .B1(_03334_),
    .B2(_03353_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _07985_ (.I0(_03351_),
    .I1(_03354_),
    .S(_02704_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07986_ (.A1(_05352_[0]),
    .A2(_05346_[0]),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _07987_ (.A1(_03153_),
    .A2(_03156_),
    .B1(_05107_[0]),
    .B2(net509),
    .C(_03356_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07988_ (.I(_03195_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _07989_ (.A1(_05306_[0]),
    .A2(_05314_[0]),
    .A3(_05322_[0]),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _07990_ (.A1(_03357_),
    .A2(_03358_),
    .B(_03255_),
    .C(_03359_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _07991_ (.I(_03299_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07992_ (.A1(_05306_[0]),
    .A2(_03361_),
    .B(_05305_[0]),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07993_ (.A1(_03252_),
    .A2(_03359_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _07994_ (.A1(_03362_),
    .A2(_03363_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07995_ (.A1(_03360_),
    .A2(_03364_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _07996_ (.A1(_05298_[0]),
    .A2(_03365_),
    .B(_05297_[0]),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _07997_ (.A1(_02991_),
    .A2(_03366_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _07998_ (.A1(_05289_[0]),
    .A2(net512),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _07999_ (.A1(_05293_[0]),
    .A2(_02973_),
    .B(_03368_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08000_ (.A1(_05290_[0]),
    .A2(_03055_),
    .B1(_03369_),
    .B2(_02968_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08001_ (.A1(_03052_),
    .A2(_03367_),
    .B(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08002_ (.I0(_03355_),
    .I1(_03371_),
    .S(_02915_),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08003_ (.A1(_05281_[0]),
    .A2(net512),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08004_ (.A1(_05285_[0]),
    .A2(_02973_),
    .B(_03372_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08005_ (.A1(_02985_),
    .A2(_03340_),
    .A3(_02988_),
    .Z(_03374_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08006_ (.A1(_03374_),
    .A2(_02994_),
    .A3(_03052_),
    .B(_03302_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08007_ (.A1(_03374_),
    .A2(_02994_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08008_ (.A1(_05282_[0]),
    .A2(_03376_),
    .A3(_03052_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08009_ (.A1(_02968_),
    .A2(_03373_),
    .B1(_03375_),
    .B2(_05282_[0]),
    .C(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08010_ (.I0(_02470_),
    .I1(net507),
    .I2(_02645_),
    .I3(net506),
    .S0(net500),
    .S1(net504),
    .Z(_03379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08011_ (.I0(_03349_),
    .I1(_03379_),
    .S(net503),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08012_ (.A1(net505),
    .A2(net496),
    .Z(_03381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08013_ (.A1(_02907_),
    .A2(_03380_),
    .B1(_03381_),
    .B2(_03151_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08014_ (.I(_03382_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08015_ (.I(_03129_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08016_ (.I0(_03384_),
    .I1(_03144_),
    .S(_02907_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08017_ (.I0(_03383_),
    .I1(_03385_),
    .S(_02919_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08018_ (.A1(_02909_),
    .A2(_03121_),
    .B(_03135_),
    .C(net505),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08019_ (.A1(_03124_),
    .A2(_03331_),
    .B1(_03334_),
    .B2(_03387_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08020_ (.I0(_03386_),
    .I1(_03388_),
    .S(net502),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08021_ (.A1(_02915_),
    .A2(_03389_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08022_ (.A1(_02915_),
    .A2(_03378_),
    .B(_03390_),
    .ZN(net67));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08023_ (.I0(_02428_),
    .I1(_02518_),
    .I2(_05303_[0]),
    .I3(_02683_),
    .S0(net500),
    .S1(net504),
    .Z(_03391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08024_ (.I0(_03379_),
    .I1(_03391_),
    .S(net503),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08025_ (.A1(_03182_),
    .A2(_03381_),
    .B1(_03392_),
    .B2(net498),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08026_ (.I0(_03163_),
    .I1(_03167_),
    .I2(_03172_),
    .I3(_03171_),
    .S0(net509),
    .S1(net498),
    .Z(_03394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08027_ (.I0(_03393_),
    .I1(_03394_),
    .S(_02919_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08028_ (.A1(net498),
    .A2(_03330_),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08029_ (.A1(net498),
    .A2(net496),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08030_ (.A1(_01288_),
    .A2(_03397_),
    .B(_03137_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08031_ (.A1(_02912_),
    .A2(_03157_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08032_ (.A1(_03161_),
    .A2(_03396_),
    .B1(_03398_),
    .B2(_03399_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08033_ (.I0(_03395_),
    .I1(_03400_),
    .S(net502),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08034_ (.A1(_03073_),
    .A2(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08035_ (.I(_05282_[0]),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08036_ (.A1(_02985_),
    .A2(_03300_),
    .B(_02994_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08037_ (.I(_05281_[0]),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08038_ (.A1(_03403_),
    .A2(_03404_),
    .B(_03405_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08039_ (.A1(_05274_[0]),
    .A2(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08040_ (.A1(_05273_[0]),
    .A2(net512),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08041_ (.A1(_05277_[0]),
    .A2(_02973_),
    .B(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08042_ (.A1(_05274_[0]),
    .A2(_03055_),
    .B1(_03409_),
    .B2(_02968_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08043_ (.A1(_03052_),
    .A2(_03407_),
    .B(_03410_),
    .C(_02915_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08044_ (.A1(_03402_),
    .A2(_03411_),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08045_ (.A1(_05265_[0]),
    .A2(net512),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08046_ (.A1(_05269_[0]),
    .A2(_02973_),
    .B(_03412_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08047_ (.A1(_02984_),
    .A2(_02990_),
    .B(_02995_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08048_ (.A1(_03414_),
    .A2(_03054_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08049_ (.A1(_03414_),
    .A2(_03052_),
    .B(_03302_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08050_ (.I0(_03415_),
    .I1(_03416_),
    .S(_05266_[0]),
    .Z(_03417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08051_ (.A1(_02968_),
    .A2(_03413_),
    .B(_03417_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08052_ (.A1(_03397_),
    .A2(_02948_),
    .B(_03398_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08053_ (.A1(_03211_),
    .A2(_03331_),
    .B(_03419_),
    .C(net502),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08054_ (.A1(_02900_),
    .A2(_02904_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _08055_ (.I0(_02382_),
    .I1(_02470_),
    .I2(net507),
    .I3(_02645_),
    .S0(net500),
    .S1(net504),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08056_ (.I0(_03391_),
    .I1(_03422_),
    .S(net503),
    .Z(_03423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08057_ (.I0(_03217_),
    .I1(_03423_),
    .S(net498),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08058_ (.A1(_03421_),
    .A2(_03424_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08059_ (.A1(net498),
    .A2(_03221_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08060_ (.A1(net498),
    .A2(_03210_),
    .B(_03426_),
    .C(_02921_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08061_ (.A1(_03073_),
    .A2(_03420_),
    .A3(_03425_),
    .A4(_03427_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08062_ (.A1(_03073_),
    .A2(_03418_),
    .B(_03428_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08063_ (.I0(_05259_[0]),
    .I1(_05275_[0]),
    .I2(_05291_[0]),
    .I3(_05307_[0]),
    .S0(net500),
    .S1(net504),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08064_ (.A1(net503),
    .A2(_03422_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08065_ (.A1(net503),
    .A2(_03429_),
    .B(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08066_ (.A1(net498),
    .A2(_02904_),
    .Z(_03432_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08067_ (.A1(net505),
    .A2(_02904_),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08068_ (.A1(_03431_),
    .A2(_03432_),
    .B1(_03433_),
    .B2(_03243_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08069_ (.A1(net498),
    .A2(_02919_),
    .A3(_03247_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08070_ (.A1(net498),
    .A2(_02904_),
    .A3(_03237_),
    .Z(_03436_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08071_ (.A1(_02900_),
    .A2(_03073_),
    .A3(_03435_),
    .A4(_03436_),
    .Z(_03437_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08072_ (.A1(_05266_[0]),
    .A2(_05290_[0]),
    .A3(_02989_),
    .Z(_03438_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08073_ (.A1(_05298_[0]),
    .A2(_03438_),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08074_ (.I(_05274_[0]),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08075_ (.A1(_05282_[0]),
    .A2(_05289_[0]),
    .B(_05281_[0]),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08076_ (.I(_05273_[0]),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08077_ (.A1(_03440_),
    .A2(_03441_),
    .B(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08078_ (.A1(_05266_[0]),
    .A2(_03443_),
    .B1(_03438_),
    .B2(_05297_[0]),
    .C(_05265_[0]),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08079_ (.I(_03444_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08080_ (.A1(_03365_),
    .A2(_03439_),
    .B(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08081_ (.A1(_05258_[0]),
    .A2(_03446_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08082_ (.A1(_05257_[0]),
    .A2(net512),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08083_ (.A1(_05261_[0]),
    .A2(_02973_),
    .B(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08084_ (.A1(_05258_[0]),
    .A2(_03055_),
    .B1(_03449_),
    .B2(_02968_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08085_ (.A1(_02915_),
    .A2(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08086_ (.A1(_03054_),
    .A2(_03447_),
    .B(_03451_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08087_ (.A1(net505),
    .A2(net504),
    .A3(_03131_),
    .Z(_03453_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08088_ (.A1(_03087_),
    .A2(_03453_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08089_ (.A1(_02907_),
    .A2(_03234_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08090_ (.A1(_03334_),
    .A2(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _08091_ (.A1(_02900_),
    .A2(net510),
    .A3(_03454_),
    .A4(_03456_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08092_ (.A1(_03434_),
    .A2(_03437_),
    .B(_03452_),
    .C(_03457_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08093_ (.A1(net505),
    .A2(_03233_),
    .B(_03333_),
    .C(_03332_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08094_ (.A1(_03122_),
    .A2(_03232_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08095_ (.A1(_03331_),
    .A2(_03334_),
    .B1(_03458_),
    .B2(_03459_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08096_ (.I0(_03274_),
    .I1(_03281_),
    .S(net505),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08097_ (.A1(_02900_),
    .A2(_02919_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_116_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08099_ (.I0(_05251_[0]),
    .I1(_05267_[0]),
    .I2(_05283_[0]),
    .I3(_05299_[0]),
    .S0(net500),
    .S1(net504),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08100_ (.I0(_03429_),
    .I1(_03464_),
    .S(net503),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08101_ (.I0(_03268_),
    .I1(_03465_),
    .S(net498),
    .Z(_03466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08102_ (.A1(_02905_),
    .A2(_03466_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08103_ (.A1(_02900_),
    .A2(_03460_),
    .B1(_03461_),
    .B2(_03462_),
    .C(_03467_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08104_ (.A1(_05249_[0]),
    .A2(net512),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08105_ (.A1(_05253_[0]),
    .A2(_02973_),
    .B(_03469_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08106_ (.A1(_05266_[0]),
    .A2(_03414_),
    .B(_05265_[0]),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08107_ (.A1(_03005_),
    .A2(_03471_),
    .B(_02997_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08108_ (.A1(_03472_),
    .A2(_03054_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08109_ (.A1(_03472_),
    .A2(_03052_),
    .B(_03302_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08110_ (.I0(_03473_),
    .I1(_03474_),
    .S(_05250_[0]),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08111_ (.A1(_02968_),
    .A2(_03470_),
    .B(_03475_),
    .C(_03073_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08112_ (.A1(_03073_),
    .A2(_03468_),
    .B(_03476_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08113_ (.A1(_05250_[0]),
    .A2(_05258_[0]),
    .A3(_03438_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08114_ (.A1(_05298_[0]),
    .A2(_03477_),
    .Z(_03478_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08115_ (.A1(_03005_),
    .A2(_03444_),
    .B(_02997_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08116_ (.A1(_05250_[0]),
    .A2(_03479_),
    .Z(_03480_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08117_ (.A1(_05249_[0]),
    .A2(_03480_),
    .Z(_03481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08118_ (.A1(_03365_),
    .A2(_03478_),
    .B(_03481_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08119_ (.A1(_05242_[0]),
    .A2(_03482_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08120_ (.A1(_03054_),
    .A2(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08121_ (.A1(_05241_[0]),
    .A2(net512),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08122_ (.A1(_05245_[0]),
    .A2(_02973_),
    .B(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08123_ (.A1(_05242_[0]),
    .A2(_03055_),
    .B1(_03486_),
    .B2(_02968_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08124_ (.A1(_02915_),
    .A2(_03484_),
    .A3(_03487_),
    .Z(_03488_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08125_ (.I(_03319_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08126_ (.I0(_03315_),
    .I1(_03489_),
    .S(net505),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08127_ (.A1(_01287_),
    .A2(_03332_),
    .Z(_03491_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08128_ (.A1(_02921_),
    .A2(_03491_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08129_ (.A1(_03160_),
    .A2(_03453_),
    .B(_03492_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08130_ (.A1(net502),
    .A2(_03490_),
    .B(_03493_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08131_ (.I0(_02236_),
    .I1(_02327_),
    .I2(_02428_),
    .I3(_02518_),
    .S0(net500),
    .S1(net504),
    .Z(_03495_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08132_ (.I0(_02284_),
    .I1(_02382_),
    .I2(_02470_),
    .I3(net507),
    .S0(net500),
    .S1(net504),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _08133_ (.I0(_03309_),
    .I1(_03310_),
    .I2(_03495_),
    .I3(_03496_),
    .S0(net509),
    .S1(_02907_),
    .Z(_03497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08134_ (.A1(_02905_),
    .A2(_03497_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08135_ (.A1(_03073_),
    .A2(_03494_),
    .A3(_03498_),
    .Z(_03499_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08136_ (.A1(_03488_),
    .A2(_03499_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08137_ (.A1(_05250_[0]),
    .A2(_03472_),
    .B(_05249_[0]),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08138_ (.I(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08139_ (.A1(_05242_[0]),
    .A2(_03501_),
    .B(_05241_[0]),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08140_ (.A1(_03054_),
    .A2(_03502_),
    .B(_03055_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08141_ (.A1(_03052_),
    .A2(_03502_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08142_ (.I0(_03503_),
    .I1(_03504_),
    .S(_03009_),
    .Z(_03505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08143_ (.A1(_05233_[0]),
    .A2(net512),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08144_ (.A1(_05237_[0]),
    .A2(_02973_),
    .B(_03506_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08145_ (.A1(_02968_),
    .A2(_03507_),
    .B(_03073_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08146_ (.I0(net508),
    .I1(_02284_),
    .I2(_02382_),
    .I3(_02470_),
    .S0(net500),
    .S1(net504),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08147_ (.I0(_03495_),
    .I1(_03509_),
    .S(net503),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08148_ (.I0(_03327_),
    .I1(_03510_),
    .S(net497),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08149_ (.A1(net502),
    .A2(_02904_),
    .Z(_03512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08150_ (.A1(_02912_),
    .A2(_03512_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08151_ (.A1(_02905_),
    .A2(_03511_),
    .B1(_03513_),
    .B2(_02898_),
    .C(net510),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08152_ (.I(_03492_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08153_ (.A1(net502),
    .A2(_02954_),
    .B(_03515_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08154_ (.A1(_03505_),
    .A2(_03508_),
    .B1(_03514_),
    .B2(_03516_),
    .ZN(net73));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08155_ (.A1(_01288_),
    .A2(net502),
    .B(_03137_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _08156_ (.I(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08157_ (.A1(net505),
    .A2(_03095_),
    .B(net502),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08158_ (.I0(_02142_),
    .I1(_02236_),
    .I2(_02327_),
    .I3(_02428_),
    .S0(net500),
    .S1(net504),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08159_ (.I0(_03509_),
    .I1(_03520_),
    .S(net503),
    .Z(_03521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08160_ (.I0(_03350_),
    .I1(_03521_),
    .S(_02907_),
    .Z(_03522_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08161_ (.A1(_02900_),
    .A2(_03330_),
    .Z(_03523_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08162_ (.A1(net505),
    .A2(_03090_),
    .A3(_03523_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08163_ (.A1(_02907_),
    .A2(_03082_),
    .A3(_03515_),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08164_ (.A1(_02905_),
    .A2(_03522_),
    .B(_03524_),
    .C(_03525_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08165_ (.A1(_03108_),
    .A2(_03513_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08166_ (.A1(_03518_),
    .A2(_03519_),
    .B(_03526_),
    .C(_03527_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08167_ (.A1(_03255_),
    .A2(_03359_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08168_ (.A1(_03194_),
    .A2(_03195_),
    .B(_03529_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08169_ (.A1(_03362_),
    .A2(_03363_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08170_ (.A1(_03530_),
    .A2(_03531_),
    .B(_03478_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08171_ (.A1(_05233_[0]),
    .A2(_05241_[0]),
    .A3(_03481_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08172_ (.A1(_05242_[0]),
    .A2(_05241_[0]),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08173_ (.A1(_05234_[0]),
    .A2(_03534_),
    .B(_05233_[0]),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08174_ (.A1(_03532_),
    .A2(_03533_),
    .B(_03535_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08175_ (.A1(_05226_[0]),
    .A2(_03536_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08176_ (.A1(_05225_[0]),
    .A2(net512),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08177_ (.A1(_05229_[0]),
    .A2(_02973_),
    .B(_03538_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08178_ (.A1(_05226_[0]),
    .A2(_03055_),
    .B1(_03539_),
    .B2(_02968_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08179_ (.A1(_03052_),
    .A2(_03537_),
    .B(_03540_),
    .C(net510),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08180_ (.A1(net510),
    .A2(_03528_),
    .B(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08181_ (.I(_03542_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08182_ (.A1(net505),
    .A2(_03136_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08183_ (.A1(_03130_),
    .A2(_03543_),
    .B(_02900_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08184_ (.A1(_03517_),
    .A2(_03544_),
    .Z(_03545_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08185_ (.I0(_02086_),
    .I1(net508),
    .I2(_02284_),
    .I3(_02382_),
    .S0(net500),
    .S1(net504),
    .Z(_03546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08186_ (.I0(_03520_),
    .I1(_03546_),
    .S(net503),
    .Z(_03547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08187_ (.I0(_03380_),
    .I1(_03547_),
    .S(_02907_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08188_ (.A1(_02905_),
    .A2(_03548_),
    .Z(_03549_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08189_ (.A1(_03151_),
    .A2(_03513_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08190_ (.A1(net510),
    .A2(_03549_),
    .A3(_03550_),
    .Z(_03551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08191_ (.A1(_02900_),
    .A2(_03132_),
    .B(_03545_),
    .C(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08192_ (.A1(_05217_[0]),
    .A2(net512),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08193_ (.A1(_05221_[0]),
    .A2(_02973_),
    .B(_03553_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08194_ (.A1(_03004_),
    .A2(_03007_),
    .A3(_03012_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08195_ (.A1(_03555_),
    .A2(_03054_),
    .Z(_03556_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08196_ (.A1(_03555_),
    .A2(_03052_),
    .B(_03302_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08197_ (.I0(_03556_),
    .I1(_03557_),
    .S(_05218_[0]),
    .Z(_03558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08198_ (.A1(_02968_),
    .A2(_03554_),
    .B(_03558_),
    .C(_03073_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08199_ (.A1(_03552_),
    .A2(_03559_),
    .ZN(net75));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08200_ (.A1(net505),
    .A2(_03159_),
    .Z(_03560_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08201_ (.A1(net502),
    .A2(_03169_),
    .A3(_03560_),
    .B(_03517_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08202_ (.I0(_02044_),
    .I1(_02142_),
    .I2(_02236_),
    .I3(_02327_),
    .S0(net500),
    .S1(net504),
    .Z(_03562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08203_ (.I0(_03546_),
    .I1(_03562_),
    .S(net503),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08204_ (.I0(_03392_),
    .I1(_03563_),
    .S(net498),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08205_ (.A1(_02905_),
    .A2(_03564_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08206_ (.A1(net505),
    .A2(_03161_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08207_ (.A1(_03169_),
    .A2(_03566_),
    .B(_03523_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08208_ (.A1(_03182_),
    .A2(_03513_),
    .B(net510),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08209_ (.A1(_03561_),
    .A2(_03565_),
    .A3(_03567_),
    .A4(_03568_),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08210_ (.A1(_05209_[0]),
    .A2(net512),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08211_ (.A1(_05213_[0]),
    .A2(_02973_),
    .B(_03570_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08212_ (.A1(_02968_),
    .A2(_03571_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08213_ (.A1(net510),
    .A2(_03572_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08214_ (.A1(_05210_[0]),
    .A2(_03052_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08215_ (.A1(_05210_[0]),
    .A2(_03054_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08216_ (.I(_05226_[0]),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08217_ (.A1(_03532_),
    .A2(_03533_),
    .B(_03535_),
    .C(_03576_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08218_ (.A1(_05217_[0]),
    .A2(_05218_[0]),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08219_ (.A1(_05217_[0]),
    .A2(_05225_[0]),
    .A3(_03577_),
    .B(_03578_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08220_ (.I0(_03574_),
    .I1(_03575_),
    .S(_03579_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08221_ (.A1(_05210_[0]),
    .A2(_03055_),
    .B(_03573_),
    .C(_03580_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08222_ (.A1(_03569_),
    .A2(_03581_),
    .Z(_03582_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08223_ (.I(_03582_),
    .ZN(net76));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08224_ (.A1(_05201_[0]),
    .A2(net512),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08225_ (.A1(_05205_[0]),
    .A2(_02973_),
    .B(_03583_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08226_ (.A1(_05218_[0]),
    .A2(_05210_[0]),
    .A3(_03555_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08227_ (.A1(_03021_),
    .A2(_03585_),
    .A3(_03052_),
    .B(_03302_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08228_ (.A1(_03021_),
    .A2(_03585_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08229_ (.A1(_05202_[0]),
    .A2(_03587_),
    .A3(_03052_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08230_ (.A1(_02968_),
    .A2(_03584_),
    .B1(_03586_),
    .B2(_05202_[0]),
    .C(_03588_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08231_ (.A1(_03212_),
    .A2(_03492_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08232_ (.I0(_01997_),
    .I1(_02044_),
    .I2(_02086_),
    .I3(_02142_),
    .S0(net509),
    .S1(net500),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08233_ (.I0(net508),
    .I1(_02236_),
    .I2(_02284_),
    .I3(_02327_),
    .S0(net509),
    .S1(net500),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08234_ (.I0(_03591_),
    .I1(_03592_),
    .S(net504),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08235_ (.A1(_02900_),
    .A2(_03593_),
    .Z(_03594_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08236_ (.A1(net502),
    .A2(_03217_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08237_ (.A1(_03594_),
    .A2(_03595_),
    .B(_03432_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08238_ (.A1(_02900_),
    .A2(_03207_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08239_ (.A1(net505),
    .A2(_02905_),
    .A3(_03423_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08240_ (.A1(_03491_),
    .A2(_03597_),
    .B(_03598_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08241_ (.A1(_03073_),
    .A2(_03590_),
    .A3(_03596_),
    .A4(_03599_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08242_ (.A1(net510),
    .A2(_03589_),
    .B(_03600_),
    .ZN(net78));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08243_ (.I0(_01947_),
    .I1(_02044_),
    .I2(_02142_),
    .I3(_02236_),
    .S0(net500),
    .S1(net504),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08244_ (.I0(_01997_),
    .I1(_02086_),
    .I2(net508),
    .I3(_02284_),
    .S0(net500),
    .S1(net504),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08245_ (.I0(_03601_),
    .I1(_03602_),
    .S(net509),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08246_ (.A1(_03431_),
    .A2(_03433_),
    .B1(_03603_),
    .B2(_03432_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08247_ (.A1(_02900_),
    .A2(_03239_),
    .A3(_03604_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08248_ (.A1(_03243_),
    .A2(_03432_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08249_ (.A1(_02900_),
    .A2(_03517_),
    .A3(_03606_),
    .Z(_03607_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08250_ (.A1(_03605_),
    .A2(_03607_),
    .B(net510),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08251_ (.A1(_05242_[0]),
    .A2(_03481_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08252_ (.A1(_05241_[0]),
    .A2(_03609_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08253_ (.A1(_05242_[0]),
    .A2(_05298_[0]),
    .A3(_03477_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08254_ (.A1(_03360_),
    .A2(_03364_),
    .B(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08255_ (.A1(_05226_[0]),
    .A2(_03014_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08256_ (.A1(_03610_),
    .A2(_03612_),
    .B(_03613_),
    .C(_05234_[0]),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08257_ (.A1(_05218_[0]),
    .A2(_05225_[0]),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08258_ (.A1(_05217_[0]),
    .A2(_03615_),
    .B(_05210_[0]),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08259_ (.A1(_03019_),
    .A2(_03616_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08260_ (.A1(_05202_[0]),
    .A2(_03617_),
    .Z(_03618_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08261_ (.A1(_05201_[0]),
    .A2(_03618_),
    .Z(_03619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08262_ (.A1(_05233_[0]),
    .A2(_03613_),
    .B(_03619_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08263_ (.A1(_03614_),
    .A2(_03620_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08264_ (.A1(_05194_[0]),
    .A2(_03052_),
    .A3(_03621_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08265_ (.A1(_05194_[0]),
    .A2(_03054_),
    .A3(_03621_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08266_ (.A1(_05193_[0]),
    .A2(_03046_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08267_ (.A1(_05197_[0]),
    .A2(_02973_),
    .B(_03624_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08268_ (.A1(_05194_[0]),
    .A2(_03055_),
    .B1(_03625_),
    .B2(_02968_),
    .C(_03073_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08269_ (.A1(_03622_),
    .A2(_03623_),
    .A3(_03626_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08270_ (.A1(_03608_),
    .A2(_03627_),
    .ZN(net79));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08271_ (.I(_05186_[0]),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08272_ (.A1(_03555_),
    .A2(_03014_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08273_ (.A1(_03022_),
    .A2(_03629_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08274_ (.A1(_05194_[0]),
    .A2(_03630_),
    .B(_05193_[0]),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08275_ (.A1(_03054_),
    .A2(_03631_),
    .B(_03055_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08276_ (.A1(_05186_[0]),
    .A2(_03052_),
    .A3(_03631_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08277_ (.A1(_05185_[0]),
    .A2(_03046_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08278_ (.A1(_05189_[0]),
    .A2(_02973_),
    .B(_03634_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08279_ (.A1(_02968_),
    .A2(_03635_),
    .B(_03073_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08280_ (.A1(_03628_),
    .A2(_03632_),
    .B(_03633_),
    .C(_03636_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08281_ (.A1(net505),
    .A2(_02919_),
    .A3(_03268_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08282_ (.A1(_03518_),
    .A2(_03638_),
    .B(_02900_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08283_ (.I0(_05187_[0]),
    .I1(_05195_[0]),
    .I2(_05203_[0]),
    .I3(_05211_[0]),
    .S0(net509),
    .S1(net500),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08284_ (.I0(_05219_[0]),
    .I1(_05227_[0]),
    .I2(_05235_[0]),
    .I3(_05243_[0]),
    .S0(net509),
    .S1(net500),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08285_ (.I0(_03640_),
    .I1(_03641_),
    .S(net504),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08286_ (.I0(_03465_),
    .I1(_03642_),
    .S(_02907_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08287_ (.A1(_03233_),
    .A2(_03517_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08288_ (.A1(_03278_),
    .A2(_03644_),
    .Z(_03645_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08289_ (.A1(_03282_),
    .A2(_03492_),
    .A3(_03645_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08290_ (.A1(_03421_),
    .A2(_03643_),
    .B(_03646_),
    .C(_03073_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08291_ (.A1(_03639_),
    .A2(_03647_),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08292_ (.A1(_03637_),
    .A2(_03648_),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08293_ (.A1(_05226_[0]),
    .A2(_03013_),
    .A3(_03014_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08294_ (.A1(_03532_),
    .A2(_03533_),
    .B(_03649_),
    .C(_03535_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08295_ (.A1(_03013_),
    .A2(_03619_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08296_ (.A1(_03017_),
    .A2(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08297_ (.A1(_03052_),
    .A2(_03650_),
    .A3(_03652_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08298_ (.A1(_03055_),
    .A2(_03653_),
    .B(_05178_[0]),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08299_ (.A1(_05177_[0]),
    .A2(_03046_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08300_ (.A1(_05181_[0]),
    .A2(_02973_),
    .B(_03655_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08301_ (.A1(_02968_),
    .A2(_03656_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08302_ (.I(_05178_[0]),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08303_ (.A1(_03650_),
    .A2(_03652_),
    .B(_03658_),
    .C(_03054_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08304_ (.A1(net510),
    .A2(_03657_),
    .A3(_03659_),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08305_ (.A1(_03333_),
    .A2(_03517_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08306_ (.A1(net504),
    .A2(_03160_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08307_ (.A1(_02900_),
    .A2(_03330_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08308_ (.A1(net505),
    .A2(_03662_),
    .B(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08309_ (.A1(net505),
    .A2(_03489_),
    .B1(_03661_),
    .B2(_03664_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08310_ (.A1(net502),
    .A2(_03491_),
    .B(net510),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08311_ (.A1(_02907_),
    .A2(_03311_),
    .A3(_03512_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08312_ (.I0(_03496_),
    .I1(_03495_),
    .S(net503),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08313_ (.I0(_01852_),
    .I1(_01899_),
    .I2(_01947_),
    .I3(_01997_),
    .S0(net509),
    .S1(net500),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08314_ (.I0(_02044_),
    .I1(_02086_),
    .I2(_02142_),
    .I3(net508),
    .S0(net509),
    .S1(net500),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08315_ (.I0(_03669_),
    .I1(_03670_),
    .S(net504),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08316_ (.I0(_03668_),
    .I1(_03671_),
    .S(_02907_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08317_ (.A1(_02905_),
    .A2(_03672_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08318_ (.A1(_03665_),
    .A2(_03666_),
    .A3(_03667_),
    .A4(_03673_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08319_ (.A1(_03654_),
    .A2(_03660_),
    .B(_03674_),
    .ZN(net81));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08320_ (.I0(_03328_),
    .I1(_03327_),
    .S(net497),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08321_ (.A1(_02904_),
    .A2(_03675_),
    .B(_03491_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08322_ (.I0(_01786_),
    .I1(_01852_),
    .I2(_01899_),
    .I3(_01947_),
    .S0(net509),
    .S1(net500),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08323_ (.I0(_03591_),
    .I1(_03677_),
    .S(_02909_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08324_ (.I0(_03510_),
    .I1(_03678_),
    .S(net497),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08325_ (.A1(_02904_),
    .A2(_03679_),
    .B(_03336_),
    .C(_02704_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08326_ (.A1(_02704_),
    .A2(_03676_),
    .B(_03680_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08327_ (.A1(_03016_),
    .A2(_03024_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08328_ (.A1(_05178_[0]),
    .A2(_03682_),
    .B(_05177_[0]),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08329_ (.A1(_03054_),
    .A2(_03683_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08330_ (.A1(_03055_),
    .A2(_03684_),
    .B(_05170_[0]),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08331_ (.A1(_05170_[0]),
    .A2(_03052_),
    .A3(_03683_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08332_ (.A1(_05169_[0]),
    .A2(_03046_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08333_ (.A1(_05173_[0]),
    .A2(_02973_),
    .B(_03687_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08334_ (.A1(_02968_),
    .A2(_03688_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08335_ (.A1(_03685_),
    .A2(_03686_),
    .A3(_03689_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08336_ (.I0(_03681_),
    .I1(_03690_),
    .S(net510),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08337_ (.A1(_03333_),
    .A2(_03517_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08338_ (.A1(_02907_),
    .A2(_03523_),
    .Z(_03692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08339_ (.A1(_03090_),
    .A2(_03692_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08340_ (.A1(_03353_),
    .A2(_03691_),
    .B(_03666_),
    .C(_03693_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08341_ (.I0(_05159_[0]),
    .I1(_01786_),
    .I2(_01852_),
    .I3(_01899_),
    .S0(net509),
    .S1(net500),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08342_ (.I0(_01947_),
    .I1(_01997_),
    .I2(_02044_),
    .I3(_02086_),
    .S0(net509),
    .S1(net500),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08343_ (.I0(_03695_),
    .I1(_03696_),
    .S(net504),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08344_ (.I0(_03348_),
    .I1(_03350_),
    .I2(_03521_),
    .I3(_03697_),
    .S0(_02907_),
    .S1(_02900_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08345_ (.A1(_02904_),
    .A2(_03698_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08346_ (.A1(_03694_),
    .A2(_03699_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08347_ (.I(_05177_[0]),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08348_ (.A1(_03658_),
    .A2(_03017_),
    .B(_03701_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08349_ (.A1(_05170_[0]),
    .A2(_03702_),
    .B(_05169_[0]),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08350_ (.A1(_05241_[0]),
    .A2(_03609_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08351_ (.A1(_05242_[0]),
    .A2(_05298_[0]),
    .A3(_03477_),
    .Z(_03705_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08352_ (.A1(_03530_),
    .A2(_03531_),
    .B(_03705_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08353_ (.A1(_05234_[0]),
    .A2(_03613_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08354_ (.A1(_03704_),
    .A2(_03706_),
    .B(_03707_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _08355_ (.I(_03620_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08356_ (.A1(_03708_),
    .A2(_03709_),
    .B(_03013_),
    .C(_03025_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08357_ (.A1(_03028_),
    .A2(_03703_),
    .A3(_03710_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08358_ (.A1(_03703_),
    .A2(_03710_),
    .B(_03028_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08359_ (.A1(_05161_[0]),
    .A2(_03046_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08360_ (.A1(_05165_[0]),
    .A2(_02973_),
    .B(_03713_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08361_ (.A1(_05162_[0]),
    .A2(_03055_),
    .B1(_03714_),
    .B2(_02968_),
    .C(_03073_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08362_ (.A1(_03052_),
    .A2(_03711_),
    .A3(_03712_),
    .B(_03715_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08363_ (.A1(_03700_),
    .A2(_03716_),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08364_ (.A1(net505),
    .A2(_03547_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08365_ (.I0(_05155_[0]),
    .I1(_05163_[0]),
    .I2(_05171_[0]),
    .I3(_05179_[0]),
    .S0(net509),
    .S1(net500),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08366_ (.I0(_03640_),
    .I1(_03718_),
    .S(_02909_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08367_ (.A1(net505),
    .A2(_03719_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08368_ (.A1(_03717_),
    .A2(_03720_),
    .B(_02919_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08369_ (.A1(_01288_),
    .A2(_03137_),
    .B1(_03382_),
    .B2(_02919_),
    .C(net502),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08370_ (.A1(net502),
    .A2(_03388_),
    .A3(_03721_),
    .B(_03722_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08371_ (.A1(_05161_[0]),
    .A2(_03027_),
    .A3(_03030_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08372_ (.A1(_03724_),
    .A2(_03052_),
    .B(_03302_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08373_ (.A1(_05154_[0]),
    .A2(_03725_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08374_ (.A1(_05153_[0]),
    .A2(_03046_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08375_ (.A1(_05157_[0]),
    .A2(_02973_),
    .B(_03727_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08376_ (.A1(_05154_[0]),
    .A2(_03052_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08377_ (.A1(_02968_),
    .A2(_03728_),
    .B1(_03729_),
    .B2(_03724_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08378_ (.A1(net510),
    .A2(_03726_),
    .A3(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08379_ (.A1(_03073_),
    .A2(_03723_),
    .B(_03731_),
    .ZN(net84));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08380_ (.A1(_05162_[0]),
    .A2(_03025_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08381_ (.A1(_05154_[0]),
    .A2(_03732_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08382_ (.A1(_03708_),
    .A2(_03709_),
    .B(_03733_),
    .C(_03013_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08383_ (.A1(_05154_[0]),
    .A2(_03732_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08384_ (.A1(_05161_[0]),
    .A2(_03030_),
    .B(_05154_[0]),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08385_ (.A1(_03017_),
    .A2(_03735_),
    .B(_03736_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08386_ (.A1(_05153_[0]),
    .A2(_03737_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08387_ (.A1(_03734_),
    .A2(_03738_),
    .B(_03052_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08388_ (.A1(_05145_[0]),
    .A2(_03046_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08389_ (.A1(_05149_[0]),
    .A2(_02973_),
    .B(_03740_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08390_ (.A1(_02968_),
    .A2(_03741_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08391_ (.A1(net510),
    .A2(_03742_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08392_ (.A1(_05146_[0]),
    .A2(_03743_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08393_ (.A1(_03614_),
    .A2(_03620_),
    .B(_03735_),
    .C(_03018_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08394_ (.I(_03738_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08395_ (.A1(_05146_[0]),
    .A2(net510),
    .A3(_03302_),
    .A4(_03742_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08396_ (.A1(_03052_),
    .A2(_03745_),
    .A3(_03746_),
    .B(_03747_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08397_ (.A1(net502),
    .A2(_03393_),
    .Z(_03749_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08398_ (.I0(_01602_),
    .I1(_01657_),
    .I2(_05159_[0]),
    .I3(_01786_),
    .S0(net509),
    .S1(net500),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08399_ (.I0(_03669_),
    .I1(_03750_),
    .S(_02909_),
    .Z(_03751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08400_ (.I0(_03563_),
    .I1(_03751_),
    .S(net498),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08401_ (.A1(net502),
    .A2(_03752_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08402_ (.I0(_01288_),
    .I1(_03157_),
    .S(net496),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08403_ (.A1(_02900_),
    .A2(_02907_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08404_ (.A1(_01287_),
    .A2(_03755_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08405_ (.A1(_03754_),
    .A2(_03755_),
    .B(_03756_),
    .C(_03137_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08406_ (.A1(_03161_),
    .A2(_03692_),
    .B(_03757_),
    .C(net510),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08407_ (.A1(_02919_),
    .A2(_03749_),
    .A3(_03753_),
    .B(_03758_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08408_ (.A1(_03739_),
    .A2(_03744_),
    .B(_03748_),
    .C(_03759_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08409_ (.I(_03760_),
    .ZN(net85));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08410_ (.A1(_03035_),
    .A2(_03052_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08411_ (.A1(_03035_),
    .A2(_03054_),
    .B(_03055_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08412_ (.I0(_03761_),
    .I1(_03762_),
    .S(_05138_[0]),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08413_ (.A1(_05137_[0]),
    .A2(_03046_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08414_ (.A1(_05141_[0]),
    .A2(_02973_),
    .B(_03764_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08415_ (.A1(_02968_),
    .A2(_03765_),
    .B(_03073_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08416_ (.A1(_03763_),
    .A2(_03766_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08417_ (.A1(_02904_),
    .A2(_03424_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08418_ (.A1(_02900_),
    .A2(_03419_),
    .B1(_03518_),
    .B2(_03768_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08419_ (.I0(_05135_[0]),
    .I1(_01602_),
    .I2(_01657_),
    .I3(_05159_[0]),
    .S0(net509),
    .S1(net500),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08420_ (.I0(_03677_),
    .I1(_03770_),
    .S(_02909_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08421_ (.I0(_03593_),
    .I1(_03771_),
    .S(net497),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08422_ (.A1(_02905_),
    .A2(_03772_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08423_ (.A1(_02909_),
    .A2(_02948_),
    .A3(_03692_),
    .Z(_03774_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08424_ (.A1(net510),
    .A2(_03769_),
    .A3(_03773_),
    .A4(_03774_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08425_ (.A1(_03767_),
    .A2(_03775_),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08426_ (.A1(_05129_[0]),
    .A2(_03046_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08427_ (.A1(_05133_[0]),
    .A2(_02973_),
    .B(_03776_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08428_ (.A1(_05130_[0]),
    .A2(_03055_),
    .B1(_03777_),
    .B2(_02968_),
    .C(_03073_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08429_ (.A1(_05138_[0]),
    .A2(_03034_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08430_ (.A1(_03018_),
    .A2(_03735_),
    .A3(_03779_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08431_ (.A1(_03614_),
    .A2(_03620_),
    .B(_03780_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08432_ (.I(_05153_[0]),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08433_ (.A1(_05145_[0]),
    .A2(_03737_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08434_ (.A1(_03782_),
    .A2(_03783_),
    .B(_03779_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08435_ (.A1(_05130_[0]),
    .A2(_05137_[0]),
    .A3(_03781_),
    .A4(_03784_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08436_ (.A1(_05137_[0]),
    .A2(_03781_),
    .A3(_03784_),
    .B(_05130_[0]),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08437_ (.A1(_03054_),
    .A2(_03785_),
    .A3(_03786_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08438_ (.A1(_03455_),
    .A2(_03691_),
    .B(_03666_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08439_ (.I0(_05127_[0]),
    .I1(_05135_[0]),
    .I2(_01602_),
    .I3(_01657_),
    .S0(net509),
    .S1(net500),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08440_ (.I0(_03695_),
    .I1(_03789_),
    .S(_02909_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08441_ (.A1(_03433_),
    .A2(_03603_),
    .B1(_03790_),
    .B2(_03432_),
    .C(_03454_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08442_ (.A1(_02900_),
    .A2(_03791_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08443_ (.A1(net502),
    .A2(_03434_),
    .B(_03792_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08444_ (.A1(_03788_),
    .A2(_03793_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08445_ (.A1(_03778_),
    .A2(_03787_),
    .B(_03794_),
    .ZN(net87));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08446_ (.I0(_05123_[0]),
    .I1(_05131_[0]),
    .I2(_05139_[0]),
    .I3(_05147_[0]),
    .S0(net509),
    .S1(net500),
    .Z(_03795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08447_ (.I0(_03718_),
    .I1(_03795_),
    .S(_02909_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08448_ (.I0(_03268_),
    .I1(_03465_),
    .I2(_03642_),
    .I3(_03796_),
    .S0(_02907_),
    .S1(_02900_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08449_ (.A1(_03661_),
    .A2(_03692_),
    .B(_03122_),
    .C(_03232_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08450_ (.A1(_03232_),
    .A2(_03755_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08451_ (.A1(_03491_),
    .A2(_03799_),
    .B(net510),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08452_ (.A1(_02919_),
    .A2(_03797_),
    .B(_03798_),
    .C(_03800_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08453_ (.A1(_05121_[0]),
    .A2(_03046_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08454_ (.A1(_05125_[0]),
    .A2(_02973_),
    .B(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08455_ (.A1(_02968_),
    .A2(_03803_),
    .B(_03073_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08456_ (.A1(_03037_),
    .A2(_03052_),
    .B(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08457_ (.A1(_05122_[0]),
    .A2(_03805_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08458_ (.A1(_03036_),
    .A2(_03761_),
    .B(_03806_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08459_ (.A1(_05122_[0]),
    .A2(_03302_),
    .A3(_03804_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08460_ (.I(_05129_[0]),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08461_ (.A1(_05138_[0]),
    .A2(_05137_[0]),
    .B(_05130_[0]),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08462_ (.A1(_03809_),
    .A2(_03054_),
    .A3(_03810_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08463_ (.I(_05137_[0]),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08464_ (.A1(_03809_),
    .A2(_03812_),
    .A3(_03035_),
    .A4(_03054_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08465_ (.A1(_03808_),
    .A2(_03811_),
    .A3(_03813_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08466_ (.A1(_03801_),
    .A2(_03807_),
    .A3(_03814_),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08467_ (.A1(_05113_[0]),
    .A2(_03046_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08468_ (.A1(_05117_[0]),
    .A2(_02973_),
    .B(_03815_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08469_ (.A1(_05114_[0]),
    .A2(_03055_),
    .B1(_03816_),
    .B2(_02968_),
    .C(_03073_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08470_ (.A1(_05138_[0]),
    .A2(_05145_[0]),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08471_ (.A1(_05137_[0]),
    .A2(_03818_),
    .B(_05130_[0]),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08472_ (.A1(_03809_),
    .A2(_03819_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08473_ (.A1(_05122_[0]),
    .A2(_03820_),
    .B(_05121_[0]),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08474_ (.A1(_05114_[0]),
    .A2(_03052_),
    .A3(_03821_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08475_ (.I0(_01287_),
    .I1(_01414_),
    .I2(_05127_[0]),
    .I3(_05135_[0]),
    .S0(net509),
    .S1(net500),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _08476_ (.I0(_03669_),
    .I1(_03670_),
    .I2(_03823_),
    .I3(_03750_),
    .S0(net504),
    .S1(_02907_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08477_ (.A1(_01287_),
    .A2(_03332_),
    .B(_02915_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08478_ (.A1(net502),
    .A2(_03160_),
    .A3(_03453_),
    .B(_03825_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08479_ (.A1(_03497_),
    .A2(_03512_),
    .B1(_03824_),
    .B2(_02905_),
    .C(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08480_ (.A1(_03817_),
    .A2(_03822_),
    .B(_03827_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08481_ (.I(_03827_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08482_ (.A1(_05130_[0]),
    .A2(_05138_[0]),
    .A3(_05146_[0]),
    .A4(_05122_[0]),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08483_ (.A1(_03013_),
    .A2(_03733_),
    .A3(_03830_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08484_ (.A1(_03708_),
    .A2(_03709_),
    .B(_03831_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08485_ (.A1(_05153_[0]),
    .A2(_03737_),
    .B(_03830_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08486_ (.A1(_05114_[0]),
    .A2(_03054_),
    .A3(_03821_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08487_ (.A1(_03829_),
    .A2(_03832_),
    .A3(_03833_),
    .A4(_03834_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08488_ (.A1(_05114_[0]),
    .A2(_03052_),
    .A3(_03827_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08489_ (.A1(_03832_),
    .A2(_03833_),
    .B(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08490_ (.A1(_03828_),
    .A2(_03835_),
    .A3(_03837_),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _08491_ (.I(net65),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08492_ (.A1(_01029_),
    .A2(_01165_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08493_ (.A1(_02004_),
    .A2(_03838_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_114_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08495_ (.I0(net100),
    .I1(_01230_),
    .S(_03839_),
    .Z(_05357_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08496_ (.I0(net111),
    .I1(_02892_),
    .S(_03839_),
    .Z(_05099_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08497_ (.I0(net122),
    .I1(_02828_),
    .S(_03839_),
    .Z(_05362_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08498_ (.I0(net125),
    .I1(_02787_),
    .S(_03839_),
    .Z(_05366_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08499_ (.I0(net126),
    .I1(_02737_),
    .S(_03839_),
    .Z(_05372_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08500_ (.I0(net127),
    .I1(_02683_),
    .S(_03839_),
    .Z(_05376_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08501_ (.I0(net128),
    .I1(_02645_),
    .S(_03839_),
    .Z(_05380_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08502_ (.I0(net129),
    .I1(_05303_[0]),
    .S(_03839_),
    .Z(_05384_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08503_ (.I0(net130),
    .I1(_02560_),
    .S(_03839_),
    .Z(_05388_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08504_ (.I0(net131),
    .I1(_02518_),
    .S(_03839_),
    .Z(_05392_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_113_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08506_ (.I0(net101),
    .I1(_02470_),
    .S(_03839_),
    .Z(_05396_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08507_ (.I0(net102),
    .I1(_02428_),
    .S(_03839_),
    .Z(_05400_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08508_ (.I0(net103),
    .I1(_02382_),
    .S(_03839_),
    .Z(_05404_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08509_ (.I0(net104),
    .I1(_02327_),
    .S(_03839_),
    .Z(_05408_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08510_ (.I0(net105),
    .I1(_02284_),
    .S(_03839_),
    .Z(_05412_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08511_ (.I0(net106),
    .I1(_02236_),
    .S(_03839_),
    .Z(_05416_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08512_ (.I0(net107),
    .I1(_02192_),
    .S(_03839_),
    .Z(_05420_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08513_ (.I0(net108),
    .I1(_02142_),
    .S(_03839_),
    .Z(_05424_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08514_ (.I0(net109),
    .I1(_02086_),
    .S(_03839_),
    .Z(_05428_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08515_ (.I0(net110),
    .I1(_02044_),
    .S(_03839_),
    .Z(_05432_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_112_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08517_ (.I0(net112),
    .I1(_01997_),
    .S(_03839_),
    .Z(_05436_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08518_ (.I0(net113),
    .I1(_01947_),
    .S(_03839_),
    .Z(_05440_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08519_ (.I0(net114),
    .I1(_01899_),
    .S(_03839_),
    .Z(_05444_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08520_ (.I0(net115),
    .I1(_01852_),
    .S(_03839_),
    .Z(_05448_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08521_ (.I0(net116),
    .I1(_01786_),
    .S(_03839_),
    .Z(_05452_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08522_ (.I0(net117),
    .I1(_05159_[0]),
    .S(_03839_),
    .Z(_05456_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08523_ (.I0(net118),
    .I1(_01657_),
    .S(_03839_),
    .Z(_05460_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08524_ (.I0(net119),
    .I1(_01602_),
    .S(_03839_),
    .Z(_05464_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08525_ (.I0(net120),
    .I1(_05135_[0]),
    .S(_03839_),
    .Z(_05468_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08526_ (.I0(net121),
    .I1(_05127_[0]),
    .S(_03839_),
    .Z(_05472_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08527_ (.I0(net123),
    .I1(_01414_),
    .S(_03839_),
    .Z(_05476_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08528_ (.I(_02893_),
    .ZN(_05358_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08529_ (.I(_02387_),
    .ZN(_05401_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08530_ (.A1(_02383_),
    .A2(_02384_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08531_ (.A1(net5),
    .A2(_02385_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08532_ (.A1(_01310_),
    .A2(_03844_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08533_ (.A1(_01310_),
    .A2(_03844_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08534_ (.I0(_03845_),
    .I1(_03846_),
    .S(_01288_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08535_ (.A1(_01329_),
    .A2(_01349_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08536_ (.A1(_01437_),
    .A2(_05131_[0]),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08537_ (.A1(_01437_),
    .A2(_05131_[0]),
    .B1(_01500_),
    .B2(_05139_[0]),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08538_ (.A1(_01287_),
    .A2(_01310_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08539_ (.A1(_03848_),
    .A2(_01414_),
    .B1(_03849_),
    .B2(_03850_),
    .C(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08540_ (.A1(_01288_),
    .A2(_01310_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08541_ (.A1(_01350_),
    .A2(_05123_[0]),
    .A3(_03853_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08542_ (.A1(_03847_),
    .A2(_03852_),
    .A3(_03854_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08543_ (.A1(_03843_),
    .A2(_03044_),
    .A3(_03855_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08544_ (.A1(_01693_),
    .A2(_05163_[0]),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08545_ (.I(_01693_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08546_ (.A1(_01735_),
    .A2(_01742_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08547_ (.A1(_03858_),
    .A2(_05159_[0]),
    .B(_03859_),
    .C(_01786_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08548_ (.A1(_01566_),
    .A2(_01602_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08549_ (.A1(_01625_),
    .A2(_01657_),
    .A3(_03861_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08550_ (.A1(_01625_),
    .A2(_01657_),
    .B(_03861_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08551_ (.A1(_03857_),
    .A2(_03860_),
    .A3(_03862_),
    .B(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08552_ (.A1(_01523_),
    .A2(_01533_),
    .B(_01500_),
    .C(_01549_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08553_ (.A1(_05127_[0]),
    .A2(_03865_),
    .B(_01414_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08554_ (.A1(_01461_),
    .A2(_01480_),
    .B(_03865_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08555_ (.A1(_01437_),
    .A2(_03867_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08556_ (.A1(_03866_),
    .A2(_03868_),
    .B(_01350_),
    .C(_03853_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08557_ (.A1(_01329_),
    .A2(_01436_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08558_ (.A1(_01461_),
    .A2(_01480_),
    .A3(_03865_),
    .B(_03870_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08559_ (.A1(_05123_[0]),
    .A2(_03867_),
    .A3(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08560_ (.A1(_01566_),
    .A2(_01602_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08561_ (.A1(_03853_),
    .A2(_03872_),
    .B(_03873_),
    .C(_03847_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08562_ (.A1(_03864_),
    .A2(_03869_),
    .A3(_03874_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08563_ (.I(_02060_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08564_ (.A1(_03876_),
    .A2(_02072_),
    .A3(_02085_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _08565_ (.I(_02015_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08566_ (.A1(_03878_),
    .A2(_03876_),
    .A3(_02072_),
    .A4(_02085_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08567_ (.A1(_02015_),
    .A2(_02028_),
    .A3(_02043_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08568_ (.A1(_05211_[0]),
    .A2(_03877_),
    .B(_03879_),
    .C(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08569_ (.A1(_02066_),
    .A2(_02068_),
    .A3(_02071_),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08570_ (.A1(net523),
    .A2(_02077_),
    .A3(_02079_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08571_ (.I(\dp.rf.rf[20][18] ),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08572_ (.A1(_01148_),
    .A2(_02082_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08573_ (.A1(_03884_),
    .A2(_01451_),
    .B(_03885_),
    .C(net8),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08574_ (.A1(\dp.rf.rf[16][18] ),
    .A2(_01467_),
    .B1(_03886_),
    .B2(net524),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08575_ (.A1(_01273_),
    .A2(_02075_),
    .B(_01216_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08576_ (.A1(_03883_),
    .A2(_03887_),
    .B(_03888_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08577_ (.A1(_03882_),
    .A2(_03889_),
    .B(_02060_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08578_ (.A1(_02142_),
    .A2(_02164_),
    .A3(net508),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08579_ (.A1(_02112_),
    .A2(_02164_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08580_ (.A1(_02112_),
    .A2(_02142_),
    .B1(net508),
    .B2(_03892_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08581_ (.A1(_05211_[0]),
    .A2(_03890_),
    .A3(_03891_),
    .A4(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08582_ (.A1(_03878_),
    .A2(_03890_),
    .A3(_03891_),
    .A4(_03893_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08583_ (.A1(_03881_),
    .A2(_03894_),
    .A3(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08584_ (.A1(_01868_),
    .A2(_01899_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _08585_ (.A1(_01954_),
    .A2(_01959_),
    .A3(_01964_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08586_ (.A1(_01947_),
    .A2(_03898_),
    .A3(_01997_),
    .B(_01916_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08587_ (.A1(_01868_),
    .A2(_01899_),
    .B1(_03898_),
    .B2(_01997_),
    .C(_01947_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08588_ (.A1(_01868_),
    .A2(_01899_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08589_ (.A1(_03897_),
    .A2(_03899_),
    .B(_03900_),
    .C(_03901_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08590_ (.A1(_01852_),
    .A2(_03902_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _08591_ (.A1(_01868_),
    .A2(_01899_),
    .B1(_01916_),
    .B2(_01947_),
    .C1(_03898_),
    .C2(_01997_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08592_ (.A1(_01868_),
    .A2(_01899_),
    .B(_01916_),
    .C(_01947_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08593_ (.A1(_03897_),
    .A2(_03904_),
    .A3(_03905_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08594_ (.A1(_01852_),
    .A2(_03906_),
    .B(_01821_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08595_ (.A1(_01625_),
    .A2(_01657_),
    .A3(_03861_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08596_ (.A1(_03859_),
    .A2(_01786_),
    .B(_01713_),
    .C(_01725_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08597_ (.A1(_01566_),
    .A2(_01602_),
    .B(_01639_),
    .C(_01656_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08598_ (.A1(_01566_),
    .A2(_01602_),
    .B(_01625_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08599_ (.A1(_01713_),
    .A2(_01725_),
    .B(_03859_),
    .C(_01786_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08600_ (.A1(_01693_),
    .A2(_03909_),
    .B1(_03910_),
    .B2(_03911_),
    .C(_03912_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _08601_ (.A1(_01566_),
    .A2(_01602_),
    .B(_03908_),
    .C(_03913_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08602_ (.A1(_03896_),
    .A2(_03903_),
    .B(_03907_),
    .C(_03914_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08603_ (.A1(_03897_),
    .A2(_03899_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08604_ (.A1(_03901_),
    .A2(_03900_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08605_ (.A1(_03916_),
    .A2(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08606_ (.A1(_01852_),
    .A2(_03906_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08607_ (.A1(_03918_),
    .A2(_03896_),
    .B(_03919_),
    .C(_03914_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08608_ (.A1(_03875_),
    .A2(_03915_),
    .A3(_03920_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08609_ (.A1(_02402_),
    .A2(_02428_),
    .B(_02443_),
    .C(_02470_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08610_ (.A1(_02402_),
    .A2(_02428_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08611_ (.A1(_03922_),
    .A2(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08612_ (.A1(_02265_),
    .A2(_02273_),
    .B(_02255_),
    .C(_02283_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08613_ (.A1(_02219_),
    .A2(_02235_),
    .A3(_03925_),
    .B(_02207_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08614_ (.A1(_02219_),
    .A2(_02235_),
    .B(_03925_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08615_ (.A1(_03926_),
    .A2(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08616_ (.A1(_02360_),
    .A2(_02368_),
    .B(_02343_),
    .C(_02381_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08617_ (.A1(_02310_),
    .A2(_02326_),
    .A3(_03929_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08618_ (.A1(_02310_),
    .A2(_02326_),
    .B(_03929_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08619_ (.A1(_02297_),
    .A2(_03930_),
    .B(_03931_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08620_ (.A1(_02532_),
    .A2(net507),
    .B(_02518_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08621_ (.A1(_02518_),
    .A2(_02532_),
    .A3(net507),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08622_ (.A1(_02402_),
    .A2(_02428_),
    .B1(_02443_),
    .B2(_02470_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08623_ (.A1(_02486_),
    .A2(_03933_),
    .B(_03934_),
    .C(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08624_ (.A1(_03924_),
    .A2(_03928_),
    .A3(_03932_),
    .A4(_03936_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08625_ (.I(_02207_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08626_ (.A1(_03938_),
    .A2(_05243_[0]),
    .B1(_02255_),
    .B2(_05251_[0]),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08627_ (.A1(_02331_),
    .A2(_02335_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08628_ (.A1(_03940_),
    .A2(_02342_),
    .B(_02382_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08629_ (.A1(_05259_[0]),
    .A2(_03941_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08630_ (.A1(_05259_[0]),
    .A2(_03941_),
    .B(_02297_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08631_ (.A1(_03939_),
    .A2(_03942_),
    .A3(_03943_),
    .B(_03928_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08632_ (.A1(_03937_),
    .A2(_03944_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08633_ (.A1(_02612_),
    .A2(_02645_),
    .B(_02582_),
    .C(_02597_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08634_ (.A1(_02582_),
    .A2(_02597_),
    .B(_02612_),
    .C(_02645_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08635_ (.A1(net162),
    .A2(_03946_),
    .B(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08636_ (.A1(_02703_),
    .A2(net506),
    .B(_02683_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08637_ (.A1(_02683_),
    .A2(_02703_),
    .A3(net506),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08638_ (.A1(net158),
    .A2(_05339_[0]),
    .B1(_03949_),
    .B2(net160),
    .C(_03950_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08639_ (.A1(_03948_),
    .A2(_03951_),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08640_ (.A1(net155),
    .A2(_05347_[0]),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08641_ (.A1(net158),
    .A2(_05339_[0]),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08642_ (.A1(_02856_),
    .A2(_02892_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08643_ (.A1(_02856_),
    .A2(_02892_),
    .B(_01088_),
    .C(_01230_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08644_ (.A1(net155),
    .A2(_05347_[0]),
    .B1(_03955_),
    .B2(_03956_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08645_ (.A1(_03953_),
    .A2(_03954_),
    .A3(_03957_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08646_ (.A1(net161),
    .A2(_05315_[0]),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08647_ (.A1(_02612_),
    .A2(_02645_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08648_ (.A1(_02703_),
    .A2(net506),
    .B(_02683_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08649_ (.A1(_02683_),
    .A2(_02703_),
    .A3(net506),
    .B(_02660_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08650_ (.A1(_03960_),
    .A2(_03961_),
    .A3(_03962_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08651_ (.A1(_03959_),
    .A2(_03963_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08652_ (.A1(net162),
    .A2(_05307_[0]),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08653_ (.A1(net162),
    .A2(_05307_[0]),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _08654_ (.A1(_03952_),
    .A2(_03958_),
    .B1(_03964_),
    .B2(_03965_),
    .C(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08655_ (.A1(_03939_),
    .A2(_03942_),
    .A3(_03943_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08656_ (.A1(_02518_),
    .A2(_02532_),
    .A3(net507),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08657_ (.A1(_02532_),
    .A2(net507),
    .B(_02518_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08658_ (.A1(_02486_),
    .A2(_03969_),
    .B(_03970_),
    .C(_03935_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08659_ (.A1(_03924_),
    .A2(_03971_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08660_ (.A1(_03968_),
    .A2(_03972_),
    .B1(_03932_),
    .B2(_03939_),
    .C(_03928_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08661_ (.A1(_03945_),
    .A2(_03967_),
    .B(_03973_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08662_ (.A1(_03921_),
    .A2(_03974_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08663_ (.A1(_03856_),
    .A2(_03975_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08664_ (.A1(_03961_),
    .A2(_03962_),
    .B1(_03959_),
    .B2(_05307_[0]),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08665_ (.A1(_05307_[0]),
    .A2(_03959_),
    .B(net162),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08666_ (.A1(_03977_),
    .A2(_03978_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08667_ (.A1(net160),
    .A2(_03949_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08668_ (.A1(_03980_),
    .A2(_03950_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08669_ (.A1(_01088_),
    .A2(_01230_),
    .B1(_02856_),
    .B2(_02892_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08670_ (.A1(net155),
    .A2(_05347_[0]),
    .B1(_03955_),
    .B2(_03982_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08671_ (.A1(_03953_),
    .A2(_03983_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08672_ (.A1(_05339_[0]),
    .A2(_03981_),
    .A3(_03984_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08673_ (.A1(_05339_[0]),
    .A2(_03984_),
    .B(_03981_),
    .C(net158),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08674_ (.A1(_03979_),
    .A2(_03985_),
    .A3(_03986_),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08675_ (.A1(_03937_),
    .A2(_03944_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08676_ (.A1(_03948_),
    .A2(_03855_),
    .A3(_03973_),
    .A4(_03988_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08677_ (.A1(_01100_),
    .A2(net4),
    .A3(_01089_),
    .A4(_02385_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08678_ (.A1(_03987_),
    .A2(_03989_),
    .B(_03990_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08679_ (.A1(_03843_),
    .A2(_02965_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08680_ (.A1(net23),
    .A2(_02003_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08681_ (.A1(_03855_),
    .A2(_03992_),
    .B(_03993_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08682_ (.A1(_03843_),
    .A2(_03044_),
    .A3(_03855_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08683_ (.A1(_02142_),
    .A2(_02164_),
    .A3(net508),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08684_ (.A1(_02112_),
    .A2(_02164_),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08685_ (.A1(_02112_),
    .A2(_02142_),
    .B1(net508),
    .B2(_03997_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08686_ (.A1(_03878_),
    .A2(_05211_[0]),
    .B1(_03996_),
    .B2(_03998_),
    .C(_03890_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08687_ (.A1(_01821_),
    .A2(_01852_),
    .B1(_03881_),
    .B2(_03999_),
    .C(_03906_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08688_ (.A1(_01821_),
    .A2(_01852_),
    .B(_03902_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08689_ (.A1(_01820_),
    .A2(_05179_[0]),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08690_ (.A1(_04000_),
    .A2(_04001_),
    .A3(_04002_),
    .B(_03914_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08691_ (.A1(_03875_),
    .A2(_04003_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08692_ (.A1(_03990_),
    .A2(_03995_),
    .B(_04004_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08693_ (.A1(_03992_),
    .A2(_03875_),
    .A3(_04003_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08694_ (.A1(_03921_),
    .A2(_03974_),
    .B(_04006_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _08695_ (.A1(_03991_),
    .A2(_03994_),
    .A3(_04005_),
    .A4(_04007_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08696_ (.A1(_03987_),
    .A2(_03989_),
    .A3(_04004_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08697_ (.A1(_01100_),
    .A2(_01089_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08698_ (.A1(net4),
    .A2(_03843_),
    .A3(_04010_),
    .A4(_03967_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08699_ (.A1(_03921_),
    .A2(_03967_),
    .B(_03990_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _08700_ (.A1(_03921_),
    .A2(_04009_),
    .A3(_04011_),
    .B(_04012_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _08701_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_109_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08703_ (.I0(_05359_[0]),
    .I1(net100),
    .S(net486),
    .Z(_00001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08704_ (.I0(_05102_[0]),
    .I1(net111),
    .S(net486),
    .Z(_00002_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_107_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_103_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_102_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_99_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_98_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_96_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_95_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_94_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_92_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_89_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_88_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_87_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_85_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_84_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_81_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_79_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place480 (.I(_04384_),
    .Z(net480));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place513 (.I(_03838_),
    .Z(net513));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place510 (.I(_02915_),
    .Z(net510));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place543 (.I(net7),
    .Z(net543));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place542 (.I(net7),
    .Z(net542));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place509 (.I(_01137_),
    .Z(net509));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place490 (.I(_04998_),
    .Z(net490));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place489 (.I(_05012_),
    .Z(net489));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place486 (.I(_04014_),
    .Z(net486));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place484 (.I(_04325_),
    .Z(net484));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place483 (.I(_04199_),
    .Z(net483));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place545 (.I(net7),
    .Z(net545));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place479 (.I(_04425_),
    .Z(net479));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk (.I(clknet_6_11__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk (.I(clknet_6_10__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk (.I(clknet_6_11__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place478 (.I(_04025_),
    .Z(net478));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08739_ (.A1(net66),
    .A2(_03063_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08740_ (.A1(net23),
    .A2(_02003_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place527 (.I(_01126_),
    .Z(net527));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08742_ (.A1(net513),
    .A2(_04019_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08744_ (.A1(net33),
    .A2(net98),
    .B(_04021_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08745_ (.A1(_05359_[0]),
    .A2(net513),
    .B1(_04019_),
    .B2(net100),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08746_ (.A1(_04018_),
    .A2(_04023_),
    .B(_04024_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _08748_ (.I(net32),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08749_ (.A1(_02684_),
    .A2(_04027_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08750_ (.A1(net2),
    .A2(_04028_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08751_ (.A1(net23),
    .A2(net28),
    .B(_01098_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08752_ (.A1(net23),
    .A2(_02384_),
    .B1(_01116_),
    .B2(_04030_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08753_ (.A1(_01030_),
    .A2(_04031_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08754_ (.A1(net31),
    .A2(_04032_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08755_ (.A1(net30),
    .A2(_04033_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08756_ (.A1(_04029_),
    .A2(_04034_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place529 (.I(net167),
    .Z(net529));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08759_ (.I0(\dp.rf.rf[10][0] ),
    .I1(net478),
    .S(_04035_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08760_ (.A1(net5),
    .A2(net99),
    .A3(_02902_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08761_ (.A1(net4),
    .A2(_04038_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08762_ (.A1(_01100_),
    .A2(net62),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _08763_ (.A1(_04039_),
    .A2(_04040_),
    .B(net98),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08764_ (.A1(net34),
    .A2(_04039_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08765_ (.A1(net513),
    .A2(_04019_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08767_ (.A1(net510),
    .A2(_03063_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08768_ (.A1(_03378_),
    .A2(_04045_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08769_ (.A1(_04041_),
    .A2(_04042_),
    .B(_04043_),
    .C(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08770_ (.I(_05399_[0]),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08771_ (.A1(_05101_[0]),
    .A2(_05365_[0]),
    .B(_05364_[0]),
    .C(_05368_[0]),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08772_ (.A1(_05369_[0]),
    .A2(_05368_[0]),
    .B(_05375_[0]),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08773_ (.A1(_05374_[0]),
    .A2(_05378_[0]),
    .A3(_05382_[0]),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08774_ (.A1(_04049_),
    .A2(_04050_),
    .B(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08775_ (.A1(_05379_[0]),
    .A2(_05378_[0]),
    .A3(_05382_[0]),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08776_ (.A1(_05383_[0]),
    .A2(_05382_[0]),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08777_ (.A1(_04053_),
    .A2(_04054_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08778_ (.A1(_04052_),
    .A2(_04055_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08779_ (.A1(_05387_[0]),
    .A2(_05391_[0]),
    .A3(_05395_[0]),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08780_ (.I(_05395_[0]),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08781_ (.A1(_05391_[0]),
    .A2(_05386_[0]),
    .B(_05390_[0]),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08782_ (.I(_05394_[0]),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08783_ (.A1(_04058_),
    .A2(_04059_),
    .B(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08784_ (.A1(_04056_),
    .A2(_04057_),
    .B(_04061_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08785_ (.A1(_04048_),
    .A2(_04062_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08786_ (.A1(net128),
    .A2(net129),
    .A3(net130),
    .A4(net131),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08787_ (.A1(net126),
    .A2(_05370_[0]),
    .A3(net127),
    .Z(_04065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08788_ (.A1(_04064_),
    .A2(_04065_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place528 (.I(net527),
    .Z(net528));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08790_ (.A1(net101),
    .A2(_04066_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_4 _08791_ (.A1(_03390_),
    .A2(_04047_),
    .B1(_04063_),
    .B2(net513),
    .C1(_04068_),
    .C2(_04019_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08793_ (.I0(\dp.rf.rf[10][10] ),
    .I1(_04069_),
    .S(_04035_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place516 (.I(_01242_),
    .Z(net516));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08795_ (.A1(net35),
    .A2(_04039_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08796_ (.A1(_03052_),
    .A2(_03407_),
    .B(_03410_),
    .C(_04045_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08797_ (.A1(_04041_),
    .A2(_04072_),
    .B(_04073_),
    .C(_03402_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08798_ (.A1(net122),
    .A2(net125),
    .A3(net126),
    .A4(net127),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08799_ (.A1(_04064_),
    .A2(_04075_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08801_ (.A1(net101),
    .A2(_04076_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08802_ (.A1(net102),
    .A2(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08803_ (.A1(_05374_[0]),
    .A2(_05378_[0]),
    .A3(_05382_[0]),
    .Z(_04080_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08804_ (.A1(_05098_[0]),
    .A2(_05361_[0]),
    .B(_05360_[0]),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08805_ (.A1(_05365_[0]),
    .A2(_05369_[0]),
    .A3(_05375_[0]),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08806_ (.A1(_05375_[0]),
    .A2(_05368_[0]),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08807_ (.A1(_05369_[0]),
    .A2(_05375_[0]),
    .A3(_05364_[0]),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08808_ (.A1(_04081_),
    .A2(_04082_),
    .B(_04083_),
    .C(_04084_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08809_ (.A1(_05399_[0]),
    .A2(_04057_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _08810_ (.A1(_04080_),
    .A2(_04085_),
    .B(_04086_),
    .C(_04055_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08811_ (.A1(_05399_[0]),
    .A2(_04061_),
    .B(_05398_[0]),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08812_ (.A1(_04087_),
    .A2(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08813_ (.A1(_05403_[0]),
    .A2(_04089_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _08814_ (.A1(_04019_),
    .A2(_04079_),
    .B1(_04090_),
    .B2(net513),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _08815_ (.A1(_04043_),
    .A2(_04074_),
    .B(_04091_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place548 (.I(net13),
    .Z(net548));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08817_ (.I0(\dp.rf.rf[10][11] ),
    .I1(_04092_),
    .S(_04035_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08818_ (.A1(net36),
    .A2(_04039_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08819_ (.A1(net98),
    .A2(net69),
    .B1(_04041_),
    .B2(_04094_),
    .C(_04043_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08820_ (.A1(_01029_),
    .A2(_01165_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place522 (.I(_01187_),
    .Z(net522));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08822_ (.I(_05398_[0]),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08823_ (.A1(_04048_),
    .A2(_04062_),
    .B(_04098_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08824_ (.A1(_05403_[0]),
    .A2(_04099_),
    .B(_05402_[0]),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08825_ (.A1(_05407_[0]),
    .A2(_04100_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08826_ (.A1(net101),
    .A2(net102),
    .A3(_04066_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08827_ (.A1(net103),
    .A2(_04102_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place526 (.I(net168),
    .Z(net526));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08829_ (.A1(_04096_),
    .A2(_04101_),
    .B1(_04103_),
    .B2(_03993_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08830_ (.A1(_04095_),
    .A2(_04105_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place520 (.I(_01245_),
    .Z(net520));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08832_ (.I0(\dp.rf.rf[10][12] ),
    .I1(_04106_),
    .S(_04035_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08833_ (.A1(net37),
    .A2(_04039_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08834_ (.A1(net98),
    .A2(net70),
    .B1(_04041_),
    .B2(_04108_),
    .C(_04043_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08835_ (.I(_05411_[0]),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08836_ (.I(_05407_[0]),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08837_ (.A1(_05403_[0]),
    .A2(_04089_),
    .B(_05402_[0]),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08838_ (.I(_05406_[0]),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08839_ (.A1(_04111_),
    .A2(_04112_),
    .B(_04113_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08840_ (.A1(_04110_),
    .A2(_04114_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08841_ (.A1(net101),
    .A2(net102),
    .A3(net103),
    .A4(_04076_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08842_ (.A1(net104),
    .A2(_04116_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08843_ (.A1(_04096_),
    .A2(_04115_),
    .B1(_04117_),
    .B2(_03993_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08844_ (.A1(_04109_),
    .A2(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place519 (.I(_01273_),
    .Z(net519));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08846_ (.I0(\dp.rf.rf[10][13] ),
    .I1(_04119_),
    .S(_04035_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08847_ (.A1(net38),
    .A2(_04039_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _08848_ (.A1(net98),
    .A2(net71),
    .B1(_04041_),
    .B2(_04121_),
    .C(_04043_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08849_ (.A1(_05403_[0]),
    .A2(_05398_[0]),
    .B(_05402_[0]),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08850_ (.A1(_04111_),
    .A2(_04123_),
    .B(_04113_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08851_ (.A1(_05411_[0]),
    .A2(_04124_),
    .B(_05410_[0]),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08852_ (.A1(_05403_[0]),
    .A2(_05407_[0]),
    .A3(_05411_[0]),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08853_ (.A1(_05399_[0]),
    .A2(_04057_),
    .A3(_04126_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08854_ (.A1(_04052_),
    .A2(_04055_),
    .A3(_04127_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08855_ (.A1(_05399_[0]),
    .A2(_04061_),
    .A3(_04126_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _08856_ (.A1(_04125_),
    .A2(_04128_),
    .A3(_04129_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08857_ (.A1(_05415_[0]),
    .A2(_04130_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08858_ (.A1(net101),
    .A2(net102),
    .A3(net103),
    .A4(net104),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08859_ (.A1(_04066_),
    .A2(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08860_ (.A1(net105),
    .A2(_04133_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _08861_ (.A1(_04096_),
    .A2(_04131_),
    .B1(_04134_),
    .B2(_03993_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08862_ (.A1(_04122_),
    .A2(_04135_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place518 (.I(_01385_),
    .Z(net518));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08864_ (.I0(\dp.rf.rf[10][14] ),
    .I1(_04136_),
    .S(_04035_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place551 (.I(net13),
    .Z(net551));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _08866_ (.A1(_03484_),
    .A2(_03487_),
    .A3(_04045_),
    .Z(_04139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08867_ (.A1(net39),
    .A2(_04039_),
    .B(_04041_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _08868_ (.A1(_03499_),
    .A2(_04021_),
    .A3(_04139_),
    .A4(_04140_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08869_ (.A1(_05407_[0]),
    .A2(_05402_[0]),
    .B(_05406_[0]),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08870_ (.I(_05410_[0]),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08871_ (.A1(_04110_),
    .A2(_04142_),
    .B(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08872_ (.A1(_04089_),
    .A2(_04126_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _08873_ (.A1(_04144_),
    .A2(_04145_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08874_ (.A1(_05415_[0]),
    .A2(_04146_),
    .B(_05414_[0]),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08875_ (.A1(_05419_[0]),
    .A2(_04147_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08876_ (.A1(net105),
    .A2(_04076_),
    .A3(_04132_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08877_ (.A1(net106),
    .A2(_04149_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _08878_ (.A1(_04096_),
    .A2(_04148_),
    .B1(_04150_),
    .B2(_03993_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08879_ (.A1(_04141_),
    .A2(_04151_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place544 (.I(net7),
    .Z(net544));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08881_ (.I0(\dp.rf.rf[10][15] ),
    .I1(_04152_),
    .S(_04035_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place541 (.I(net7),
    .Z(net541));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _08883_ (.A1(_04029_),
    .A2(_04034_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place525 (.I(net166),
    .Z(net525));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place537 (.I(net9),
    .Z(net537));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08886_ (.I0(net62),
    .I1(net39),
    .S(net4),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08887_ (.A1(_01100_),
    .A2(_04158_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _08888_ (.A1(_04038_),
    .A2(_04159_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place540 (.I(net7),
    .Z(net540));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08890_ (.A1(net40),
    .A2(_04038_),
    .B(_04160_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08891_ (.A1(_03063_),
    .A2(_04162_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08892_ (.A1(_03063_),
    .A2(net73),
    .B(_04021_),
    .C(_04163_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08893_ (.A1(_03856_),
    .A2(_03975_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08894_ (.A1(_03991_),
    .A2(_03994_),
    .A3(_04005_),
    .A4(_04007_),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08895_ (.A1(net105),
    .A2(net106),
    .A3(_04066_),
    .A4(_04132_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08896_ (.A1(net107),
    .A2(_04167_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08897_ (.A1(_04021_),
    .A2(_04168_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08898_ (.A1(_04165_),
    .A2(_04166_),
    .B(_04169_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08899_ (.I(_05423_[0]),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08900_ (.I(_05418_[0]),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08901_ (.A1(_05415_[0]),
    .A2(_04130_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08902_ (.A1(_05414_[0]),
    .A2(_04173_),
    .B(_05419_[0]),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08903_ (.A1(_04172_),
    .A2(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08904_ (.A1(_04171_),
    .A2(_04175_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _08905_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04043_),
    .A4(_04176_),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08906_ (.A1(_04164_),
    .A2(_04170_),
    .A3(_04177_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08907_ (.A1(\dp.rf.rf[10][16] ),
    .A2(_04155_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08908_ (.A1(_04155_),
    .A2(_04178_),
    .B(_04179_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08909_ (.A1(_03063_),
    .A2(_04043_),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08910_ (.A1(_05419_[0]),
    .A2(_05414_[0]),
    .B(_05418_[0]),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08911_ (.I(_05422_[0]),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08912_ (.A1(_04171_),
    .A2(_04181_),
    .B(_04182_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08913_ (.A1(_05427_[0]),
    .A2(_04183_),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08914_ (.A1(_05415_[0]),
    .A2(_05419_[0]),
    .A3(_05423_[0]),
    .A4(_05427_[0]),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08915_ (.A1(_04144_),
    .A2(_04185_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08916_ (.A1(_04184_),
    .A2(_04186_),
    .Z(_04187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08917_ (.I(_04126_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _08918_ (.A1(_05415_[0]),
    .A2(_05419_[0]),
    .A3(_05423_[0]),
    .A4(_05427_[0]),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08919_ (.A1(_04087_),
    .A2(_04088_),
    .B(_04188_),
    .C(_04189_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08920_ (.A1(_05415_[0]),
    .A2(_05419_[0]),
    .A3(_05423_[0]),
    .A4(_04146_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _08921_ (.A1(_05427_[0]),
    .A2(_04183_),
    .A3(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08922_ (.A1(_04187_),
    .A2(_04190_),
    .A3(_04192_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08923_ (.A1(net41),
    .A2(_04038_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08924_ (.A1(net105),
    .A2(net106),
    .A3(net107),
    .A4(_04132_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08925_ (.A1(_04076_),
    .A2(_04195_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08926_ (.A1(net108),
    .A2(_04196_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _08927_ (.A1(_03063_),
    .A2(_04160_),
    .A3(_04194_),
    .B1(_04197_),
    .B2(_04019_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08928_ (.A1(_03542_),
    .A2(_04180_),
    .B1(_04193_),
    .B2(_04096_),
    .C(_04198_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place515 (.I(_01475_),
    .Z(net515));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08930_ (.I0(\dp.rf.rf[10][17] ),
    .I1(net483),
    .S(_04035_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08931_ (.A1(_03063_),
    .A2(_04043_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08932_ (.A1(net108),
    .A2(_04195_),
    .Z(_04202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08933_ (.A1(_04066_),
    .A2(_04202_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08934_ (.A1(net109),
    .A2(_04203_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08935_ (.I(_05427_[0]),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08936_ (.A1(_05423_[0]),
    .A2(_04175_),
    .B(_05422_[0]),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08937_ (.I(_05426_[0]),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08938_ (.A1(_04205_),
    .A2(_04206_),
    .B(_04207_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08939_ (.A1(_05431_[0]),
    .A2(_04208_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08940_ (.A1(net42),
    .A2(_04038_),
    .B(_04160_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08941_ (.A1(_03063_),
    .A2(_04210_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _08942_ (.A1(_03993_),
    .A2(_04204_),
    .B1(_04209_),
    .B2(_04096_),
    .C(_04211_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08943_ (.A1(_03552_),
    .A2(_03559_),
    .A3(_04201_),
    .B(_04212_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place521 (.I(_01187_),
    .Z(net521));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08945_ (.I0(\dp.rf.rf[10][18] ),
    .I1(net482),
    .S(_04035_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08946_ (.A1(net43),
    .A2(_04038_),
    .B(_04160_),
    .C(_03063_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08947_ (.A1(_05426_[0]),
    .A2(_04187_),
    .A3(_04190_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08948_ (.A1(_05431_[0]),
    .A2(_04216_),
    .B(_05430_[0]),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08949_ (.A1(_05435_[0]),
    .A2(_04217_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08950_ (.A1(net109),
    .A2(_04076_),
    .A3(_04202_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08951_ (.A1(net110),
    .A2(_04219_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _08952_ (.A1(net513),
    .A2(_04218_),
    .B1(_04220_),
    .B2(_04019_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08953_ (.A1(_03582_),
    .A2(_04180_),
    .B(_04215_),
    .C(_04221_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place514 (.I(_01475_),
    .Z(net514));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08955_ (.I0(\dp.rf.rf[10][19] ),
    .I1(_04222_),
    .S(_04035_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08956_ (.I(_05102_[0]),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08957_ (.A1(net44),
    .A2(net98),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08958_ (.A1(_03063_),
    .A2(net77),
    .B(_04021_),
    .C(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08959_ (.A1(net111),
    .A2(_04019_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _08960_ (.A1(_04224_),
    .A2(_04096_),
    .B(_04226_),
    .C(_04227_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place534 (.I(net9),
    .Z(net534));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place533 (.I(_01030_),
    .Z(net533));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _08963_ (.I0(\dp.rf.rf[10][1] ),
    .I1(_04228_),
    .S(_04035_),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08964_ (.A1(net45),
    .A2(_04038_),
    .B(_04160_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08965_ (.A1(_03063_),
    .A2(_04231_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08966_ (.A1(_03063_),
    .A2(net78),
    .B(_04021_),
    .C(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _08967_ (.A1(net108),
    .A2(net109),
    .A3(net110),
    .A4(_04195_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _08968_ (.A1(_04066_),
    .A2(_04234_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08969_ (.A1(net112),
    .A2(_04235_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08970_ (.A1(_04021_),
    .A2(_04236_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08971_ (.A1(_04165_),
    .A2(_04166_),
    .B(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08972_ (.I(_05439_[0]),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _08973_ (.A1(_05415_[0]),
    .A2(_05419_[0]),
    .A3(_05423_[0]),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08974_ (.A1(_04171_),
    .A2(_04181_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08975_ (.A1(_05422_[0]),
    .A2(_05426_[0]),
    .A3(_05430_[0]),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _08976_ (.A1(_04130_),
    .A2(_04240_),
    .B(_04241_),
    .C(_04242_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _08977_ (.A1(_05431_[0]),
    .A2(_05430_[0]),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08978_ (.A1(_05427_[0]),
    .A2(_05426_[0]),
    .A3(_05430_[0]),
    .B(_04244_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _08979_ (.A1(_04243_),
    .A2(_04245_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08980_ (.A1(_05435_[0]),
    .A2(_04246_),
    .B(_05434_[0]),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08981_ (.A1(_04239_),
    .A2(_04247_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _08982_ (.A1(_04165_),
    .A2(_04166_),
    .A3(_04021_),
    .A4(_04248_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _08983_ (.A1(_04233_),
    .A2(_04238_),
    .A3(_04249_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08984_ (.A1(\dp.rf.rf[10][20] ),
    .A2(_04155_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08985_ (.A1(_04155_),
    .A2(_04250_),
    .B(_04251_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08986_ (.A1(net46),
    .A2(_04038_),
    .B(_04160_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _08987_ (.A1(_03608_),
    .A2(_03627_),
    .A3(_04201_),
    .B1(_04252_),
    .B2(_03063_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _08988_ (.A1(net112),
    .A2(_04234_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08989_ (.A1(_04076_),
    .A2(_04254_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _08990_ (.A1(net113),
    .A2(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _08991_ (.A1(_04021_),
    .A2(_04256_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08992_ (.A1(_04165_),
    .A2(_04166_),
    .B(_04257_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _08993_ (.A1(_05426_[0]),
    .A2(_05430_[0]),
    .A3(_05434_[0]),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _08994_ (.A1(_05435_[0]),
    .A2(_04244_),
    .B(_05434_[0]),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08995_ (.I(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _08996_ (.A1(_04187_),
    .A2(_04190_),
    .A3(_04259_),
    .B(_04261_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _08997_ (.I(_05438_[0]),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _08998_ (.A1(_04239_),
    .A2(_04262_),
    .B(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _08999_ (.A1(_05443_[0]),
    .A2(_04264_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09000_ (.A1(_04165_),
    .A2(_04166_),
    .A3(_04021_),
    .A4(_04265_),
    .Z(_04266_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09001_ (.A1(_04253_),
    .A2(_04258_),
    .A3(_04266_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place523 (.I(_01180_),
    .Z(net523));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09003_ (.I0(\dp.rf.rf[10][21] ),
    .I1(_04267_),
    .S(_04035_),
    .Z(_00048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09004_ (.A1(_04165_),
    .A2(_04166_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09005_ (.A1(net113),
    .A2(_04066_),
    .A3(_04254_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09006_ (.A1(net114),
    .A2(_04270_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09007_ (.A1(_04043_),
    .A2(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09008_ (.A1(_05435_[0]),
    .A2(_05439_[0]),
    .A3(_05443_[0]),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09009_ (.A1(_05439_[0]),
    .A2(_05443_[0]),
    .A3(_05434_[0]),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09010_ (.A1(_05443_[0]),
    .A2(_05438_[0]),
    .B(_04274_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _09011_ (.A1(_04243_),
    .A2(_04245_),
    .A3(_04273_),
    .B(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09012_ (.A1(_05442_[0]),
    .A2(_04276_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09013_ (.A1(_05447_[0]),
    .A2(_04277_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _09014_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04043_),
    .A4(_04278_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09015_ (.A1(_03063_),
    .A2(_03637_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09016_ (.A1(net47),
    .A2(_04038_),
    .B(_04160_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09017_ (.A1(_03063_),
    .A2(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09018_ (.A1(_03648_),
    .A2(_04280_),
    .B(_04282_),
    .C(_04021_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09019_ (.A1(_04269_),
    .A2(_04272_),
    .B(_04279_),
    .C(_04283_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place524 (.I(_01177_),
    .Z(net524));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09021_ (.I0(\dp.rf.rf[10][22] ),
    .I1(net481),
    .S(_04035_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09022_ (.I(\dp.rf.rf[10][23] ),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09023_ (.A1(net113),
    .A2(net114),
    .A3(_04076_),
    .A4(_04254_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09024_ (.A1(net115),
    .A2(_04287_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09025_ (.A1(_04021_),
    .A2(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09026_ (.A1(_05439_[0]),
    .A2(_05443_[0]),
    .A3(_05447_[0]),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09027_ (.A1(_05443_[0]),
    .A2(_05447_[0]),
    .A3(_05438_[0]),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09028_ (.A1(_05447_[0]),
    .A2(_05442_[0]),
    .B(_04291_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09029_ (.I(_05446_[0]),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09030_ (.A1(_04262_),
    .A2(_04290_),
    .B(_04292_),
    .C(_04293_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09031_ (.A1(_05451_[0]),
    .A2(_04294_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09032_ (.A1(_04021_),
    .A2(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09033_ (.I0(_04289_),
    .I1(_04296_),
    .S(_04014_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place511 (.I(_01110_),
    .Z(net511));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09035_ (.A1(net48),
    .A2(_04038_),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09036_ (.A1(_03063_),
    .A2(_04160_),
    .A3(_04299_),
    .Z(_04300_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09037_ (.A1(net98),
    .A2(net81),
    .B(_04043_),
    .C(_04300_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09038_ (.A1(_04035_),
    .A2(_04301_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09039_ (.A1(_04286_),
    .A2(_04155_),
    .B1(net485),
    .B2(_04302_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _09040_ (.A1(net113),
    .A2(net114),
    .A3(net115),
    .A4(_04254_),
    .Z(_04303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09041_ (.A1(_04066_),
    .A2(_04303_),
    .Z(_04304_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09042_ (.A1(net116),
    .A2(_04304_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09043_ (.A1(_05442_[0]),
    .A2(_05446_[0]),
    .A3(_05450_[0]),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _09044_ (.A1(_05447_[0]),
    .A2(_05446_[0]),
    .A3(_05450_[0]),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _09045_ (.A1(_05451_[0]),
    .A2(_05450_[0]),
    .B1(_04276_),
    .B2(_04306_),
    .C(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09046_ (.A1(_05455_[0]),
    .A2(_04308_),
    .Z(_04309_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09047_ (.A1(_03685_),
    .A2(_03686_),
    .A3(_03689_),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09048_ (.A1(net49),
    .A2(_04038_),
    .B(_04160_),
    .C(_03063_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09049_ (.A1(_04310_),
    .A2(_04045_),
    .B(_04311_),
    .C(_04021_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09050_ (.A1(net510),
    .A2(_03681_),
    .B(_04312_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _09051_ (.A1(_04019_),
    .A2(_04305_),
    .B1(_04309_),
    .B2(net513),
    .C(_04313_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place539 (.I(net7),
    .Z(net539));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09053_ (.I0(\dp.rf.rf[10][24] ),
    .I1(_04314_),
    .S(_04035_),
    .Z(_00051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09054_ (.I(\dp.rf.rf[10][25] ),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09055_ (.A1(net116),
    .A2(_04076_),
    .A3(_04303_),
    .Z(_04317_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09056_ (.A1(net117),
    .A2(_04317_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place536 (.I(net9),
    .Z(net536));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09058_ (.A1(_05451_[0]),
    .A2(_05455_[0]),
    .A3(_04294_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09059_ (.A1(_05455_[0]),
    .A2(_05450_[0]),
    .Z(_04321_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09060_ (.A1(_05454_[0]),
    .A2(_04320_),
    .A3(_04321_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09061_ (.A1(_05459_[0]),
    .A2(_04322_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09062_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04013_),
    .A4(_04323_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09063_ (.A1(_04014_),
    .A2(_04318_),
    .B(_04324_),
    .C(_04021_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place508 (.I(_02192_),
    .Z(net508));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _09065_ (.A1(_03700_),
    .A2(_03716_),
    .A3(_04180_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09066_ (.A1(net50),
    .A2(_04038_),
    .Z(_04328_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09067_ (.A1(_04160_),
    .A2(_04328_),
    .B(net98),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09068_ (.A1(_04035_),
    .A2(_04327_),
    .A3(_04329_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09069_ (.A1(_04316_),
    .A2(_04155_),
    .B1(_04325_),
    .B2(_04330_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09070_ (.A1(_05455_[0]),
    .A2(_05459_[0]),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09071_ (.A1(_05459_[0]),
    .A2(_05454_[0]),
    .B(_05458_[0]),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09072_ (.A1(_04308_),
    .A2(_04331_),
    .B(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09073_ (.A1(_05463_[0]),
    .A2(_04333_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09074_ (.A1(_04096_),
    .A2(_04334_),
    .Z(_04335_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09075_ (.A1(net84),
    .A2(_04180_),
    .Z(_04336_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09076_ (.A1(net116),
    .A2(net117),
    .A3(_04303_),
    .Z(_04337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09077_ (.A1(_04066_),
    .A2(_04337_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09078_ (.A1(net118),
    .A2(_04338_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09079_ (.A1(_03993_),
    .A2(_04339_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09080_ (.A1(net51),
    .A2(_04038_),
    .B(_04160_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09081_ (.A1(_03063_),
    .A2(_04341_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09082_ (.A1(_04335_),
    .A2(_04336_),
    .A3(_04340_),
    .A4(_04342_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place507 (.I(_02560_),
    .Z(net507));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09084_ (.I0(\dp.rf.rf[10][26] ),
    .I1(_04343_),
    .S(_04035_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09085_ (.A1(net52),
    .A2(_04038_),
    .B(_04160_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09086_ (.I0(_03760_),
    .I1(_04345_),
    .S(net98),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09087_ (.A1(net118),
    .A2(_04337_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09088_ (.A1(_04076_),
    .A2(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09089_ (.A1(net119),
    .A2(_04348_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09090_ (.A1(_05459_[0]),
    .A2(_04322_),
    .Z(_04350_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09091_ (.A1(_05458_[0]),
    .A2(_04350_),
    .Z(_04351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09092_ (.A1(_05463_[0]),
    .A2(_04351_),
    .B(_05462_[0]),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09093_ (.A1(_05467_[0]),
    .A2(_04352_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _09094_ (.A1(_04019_),
    .A2(_04349_),
    .B1(_04353_),
    .B2(net513),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09095_ (.A1(_04043_),
    .A2(_04346_),
    .B(_04354_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place535 (.I(net9),
    .Z(net535));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09097_ (.I0(\dp.rf.rf[10][27] ),
    .I1(_04355_),
    .S(_04035_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09098_ (.A1(_05463_[0]),
    .A2(_04333_),
    .Z(_04357_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09099_ (.A1(_05462_[0]),
    .A2(_04357_),
    .Z(_04358_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09100_ (.A1(_05467_[0]),
    .A2(_04358_),
    .B(_05466_[0]),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09101_ (.A1(_05471_[0]),
    .A2(_04359_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _09102_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04043_),
    .A4(_04360_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09103_ (.A1(net119),
    .A2(_04347_),
    .Z(_04362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09104_ (.A1(_04066_),
    .A2(_04362_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09105_ (.A1(net120),
    .A2(_04363_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09106_ (.A1(_04021_),
    .A2(_04364_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09107_ (.A1(_04165_),
    .A2(_04166_),
    .B(_04365_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09108_ (.A1(_03767_),
    .A2(_03775_),
    .A3(_04180_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09109_ (.A1(net53),
    .A2(_04038_),
    .B(_04160_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _09110_ (.A1(_03063_),
    .A2(_04368_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09111_ (.A1(_04361_),
    .A2(_04366_),
    .A3(_04367_),
    .A4(_04369_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place530 (.I(_01208_),
    .Z(net530));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09113_ (.I0(\dp.rf.rf[10][28] ),
    .I1(_04370_),
    .S(_04035_),
    .Z(_00055_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09114_ (.I(\dp.rf.rf[10][29] ),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09115_ (.A1(net120),
    .A2(_04362_),
    .Z(_04373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09116_ (.A1(_04076_),
    .A2(_04373_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09117_ (.A1(net121),
    .A2(_04374_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _09118_ (.A1(_05463_[0]),
    .A2(_05467_[0]),
    .A3(_05471_[0]),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09119_ (.I(_05470_[0]),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09120_ (.A1(_05467_[0]),
    .A2(_05462_[0]),
    .Z(_04378_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09121_ (.A1(_05466_[0]),
    .A2(_04378_),
    .B(_05471_[0]),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09122_ (.A1(_04377_),
    .A2(_04379_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09123_ (.A1(_04351_),
    .A2(_04376_),
    .B(_04380_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09124_ (.A1(_05475_[0]),
    .A2(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09125_ (.A1(_03976_),
    .A2(_04008_),
    .A3(net487),
    .A4(_04382_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09126_ (.A1(net486),
    .A2(_04375_),
    .B(_04383_),
    .C(_04021_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place538 (.I(net7),
    .Z(net538));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09128_ (.I(_03778_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _09129_ (.A1(_03054_),
    .A2(_03785_),
    .A3(_03786_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _09130_ (.A1(_03788_),
    .A2(_03793_),
    .B1(_04386_),
    .B2(_04387_),
    .C(_04180_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09131_ (.A1(net54),
    .A2(_04038_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _09132_ (.A1(_04160_),
    .A2(_04389_),
    .B(net98),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09133_ (.A1(_04035_),
    .A2(_04388_),
    .A3(_04390_),
    .Z(_04391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09134_ (.A1(_04372_),
    .A2(_04155_),
    .B1(net480),
    .B2(_04391_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09135_ (.A1(_05101_[0]),
    .A2(_05365_[0]),
    .Z(_04392_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09136_ (.I(net122),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _09137_ (.A1(net55),
    .A2(net98),
    .B1(_04096_),
    .B2(_04392_),
    .C1(_03993_),
    .C2(_04393_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09138_ (.A1(net88),
    .A2(_04180_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09139_ (.A1(_04394_),
    .A2(_04395_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place506 (.I(_02737_),
    .Z(net506));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09141_ (.I0(\dp.rf.rf[10][2] ),
    .I1(_04396_),
    .S(_04035_),
    .Z(_00057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09142_ (.A1(net121),
    .A2(_04373_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09143_ (.A1(_04066_),
    .A2(_04398_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09144_ (.A1(net123),
    .A2(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09145_ (.A1(_04021_),
    .A2(_04400_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09146_ (.I(_05475_[0]),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09147_ (.A1(_04333_),
    .A2(_04376_),
    .B(_04380_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09148_ (.I(_05474_[0]),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09149_ (.A1(_04402_),
    .A2(_04403_),
    .B(_04404_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09150_ (.A1(_05479_[0]),
    .A2(_04405_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09151_ (.A1(_04021_),
    .A2(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09152_ (.A1(net56),
    .A2(_04038_),
    .Z(_04408_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09153_ (.A1(_04160_),
    .A2(_04408_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09154_ (.I0(net89),
    .I1(_04409_),
    .S(net98),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _09155_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04407_),
    .B1(_04410_),
    .B2(_04021_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09156_ (.A1(_04269_),
    .A2(_04401_),
    .B(_04411_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place505 (.I(_02753_),
    .Z(net505));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09158_ (.I0(\dp.rf.rf[10][30] ),
    .I1(net477),
    .S(_04035_),
    .Z(_00058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09159_ (.I(\dp.rf.rf[10][31] ),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09160_ (.A1(net123),
    .A2(_04076_),
    .A3(_04398_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09161_ (.A1(net124),
    .A2(_04415_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09162_ (.I0(net124),
    .I1(_01287_),
    .S(_03839_),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09163_ (.A1(_05459_[0]),
    .A2(_05475_[0]),
    .A3(_04322_),
    .A4(_04376_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09164_ (.A1(_05475_[0]),
    .A2(_04380_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09165_ (.A1(_05475_[0]),
    .A2(_05458_[0]),
    .A3(_04376_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _09166_ (.A1(_05474_[0]),
    .A2(_04418_),
    .A3(_04419_),
    .A4(_04420_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09167_ (.A1(_05479_[0]),
    .A2(_04421_),
    .B(_05478_[0]),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _09168_ (.A1(net25),
    .A2(_04417_),
    .A3(_04422_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _09169_ (.A1(_03976_),
    .A2(_04008_),
    .A3(net487),
    .A4(_04423_),
    .Z(_04424_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09170_ (.A1(net486),
    .A2(_04416_),
    .B(_04424_),
    .C(_04021_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place532 (.I(_01101_),
    .Z(net532));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09172_ (.A1(net57),
    .A2(_04038_),
    .Z(_04427_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09173_ (.A1(_03063_),
    .A2(_04160_),
    .A3(_04427_),
    .Z(_04428_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _09174_ (.A1(net98),
    .A2(net90),
    .B(_04043_),
    .C(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09175_ (.A1(_04035_),
    .A2(_04429_),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09176_ (.A1(_04414_),
    .A2(_04155_),
    .B1(net479),
    .B2(_04430_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09177_ (.I(_04081_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09178_ (.A1(_05365_[0]),
    .A2(_04431_),
    .B(_05364_[0]),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09179_ (.A1(_05369_[0]),
    .A2(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _09180_ (.A1(net58),
    .A2(net98),
    .B1(_04096_),
    .B2(_04433_),
    .C1(_03993_),
    .C2(_05371_[0]),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _09181_ (.A1(_03184_),
    .A2(_03206_),
    .A3(_04180_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09182_ (.A1(_04434_),
    .A2(_04435_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place512 (.I(_03046_),
    .Z(net512));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09184_ (.I0(\dp.rf.rf[10][3] ),
    .I1(_04436_),
    .S(_04035_),
    .Z(_00060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09185_ (.A1(net59),
    .A2(net98),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09186_ (.A1(net98),
    .A2(_03230_),
    .B(_04043_),
    .C(_04438_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09187_ (.A1(net126),
    .A2(_05370_[0]),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09188_ (.A1(_05101_[0]),
    .A2(_05365_[0]),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09189_ (.A1(_05364_[0]),
    .A2(_04441_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09190_ (.A1(_05369_[0]),
    .A2(_04442_),
    .B(_05368_[0]),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09191_ (.A1(_05375_[0]),
    .A2(_04443_),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09192_ (.A1(_03993_),
    .A2(_04440_),
    .B1(_04444_),
    .B2(_04096_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09193_ (.A1(_04439_),
    .A2(_04445_),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place531 (.I(_01148_),
    .Z(net531));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09195_ (.I0(\dp.rf.rf[10][4] ),
    .I1(_04446_),
    .S(_04035_),
    .Z(_00061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09196_ (.A1(net60),
    .A2(net98),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _09197_ (.A1(net98),
    .A2(_03263_),
    .B(_04043_),
    .C(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09198_ (.A1(net122),
    .A2(net125),
    .A3(net126),
    .Z(_04450_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09199_ (.A1(net127),
    .A2(_04450_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09200_ (.A1(_05374_[0]),
    .A2(_04085_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09201_ (.A1(_05379_[0]),
    .A2(_04452_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _09202_ (.A1(_03993_),
    .A2(_04451_),
    .B1(_04453_),
    .B2(_04096_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09203_ (.A1(_04449_),
    .A2(_04454_),
    .Z(_04455_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place504 (.I(_02803_),
    .Z(net504));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09205_ (.I0(\dp.rf.rf[10][5] ),
    .I1(_04455_),
    .S(_04035_),
    .Z(_00062_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09206_ (.A1(net128),
    .A2(_04065_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09207_ (.A1(_04165_),
    .A2(_04166_),
    .B(_04043_),
    .C(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09208_ (.I(_05374_[0]),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09209_ (.A1(_04049_),
    .A2(_04050_),
    .B(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09210_ (.A1(_05379_[0]),
    .A2(_04460_),
    .B(_05378_[0]),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09211_ (.A1(_05383_[0]),
    .A2(_04461_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _09212_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04043_),
    .A4(_04462_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09213_ (.A1(net61),
    .A2(net98),
    .Z(_04464_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09214_ (.A1(_03063_),
    .A2(net94),
    .B(_04021_),
    .C(_04464_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09215_ (.A1(_04458_),
    .A2(_04463_),
    .A3(_04465_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09216_ (.A1(\dp.rf.rf[10][6] ),
    .A2(_04155_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09217_ (.A1(_04155_),
    .A2(_04466_),
    .B(_04467_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09218_ (.A1(_04080_),
    .A2(_04085_),
    .B(_04055_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09219_ (.A1(_05387_[0]),
    .A2(_04468_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09220_ (.A1(net128),
    .A2(_04075_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09221_ (.A1(net129),
    .A2(_04470_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_4 _09222_ (.A1(net62),
    .A2(_03063_),
    .B1(net513),
    .B2(_04469_),
    .C1(_04471_),
    .C2(_04019_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _09223_ (.A1(_03325_),
    .A2(_04180_),
    .B(_04472_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place550 (.I(net13),
    .Z(net550));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09225_ (.I0(\dp.rf.rf[10][7] ),
    .I1(_04473_),
    .S(_04035_),
    .Z(_00064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09226_ (.A1(net63),
    .A2(_04039_),
    .B(_04041_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09227_ (.A1(_03345_),
    .A2(_04045_),
    .B(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09228_ (.A1(_02915_),
    .A2(_03337_),
    .B(_04476_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09229_ (.A1(_04043_),
    .A2(_04477_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09230_ (.A1(net128),
    .A2(net129),
    .A3(_04065_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09231_ (.A1(net130),
    .A2(_04479_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _09232_ (.A1(_04165_),
    .A2(_04166_),
    .B(_04043_),
    .C(_04480_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09233_ (.A1(_05387_[0]),
    .A2(_04056_),
    .B(_05386_[0]),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09234_ (.A1(_05391_[0]),
    .A2(_04482_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _09235_ (.A1(_03976_),
    .A2(_04008_),
    .A3(_04043_),
    .A4(_04483_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09236_ (.A1(_04478_),
    .A2(_04481_),
    .A3(_04484_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09237_ (.A1(\dp.rf.rf[10][8] ),
    .A2(_04155_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09238_ (.A1(_04155_),
    .A2(_04485_),
    .B(_04486_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09239_ (.A1(net64),
    .A2(_04039_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _09240_ (.A1(net98),
    .A2(net97),
    .B1(_04041_),
    .B2(_04487_),
    .C(_04043_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _09241_ (.A1(net128),
    .A2(net129),
    .A3(net130),
    .A4(_04075_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _09242_ (.A1(net131),
    .A2(_04489_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09243_ (.I(_04468_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09244_ (.A1(_05387_[0]),
    .A2(_04491_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _09245_ (.A1(_05386_[0]),
    .A2(_04492_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _09246_ (.A1(_05391_[0]),
    .A2(_04493_),
    .B(_05390_[0]),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _09247_ (.A1(_05395_[0]),
    .A2(_04494_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09248_ (.A1(_03993_),
    .A2(_04490_),
    .B1(_04495_),
    .B2(_04096_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09249_ (.A1(_04488_),
    .A2(_04496_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place503 (.I(_02894_),
    .Z(net503));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09251_ (.I0(\dp.rf.rf[10][9] ),
    .I1(_04497_),
    .S(_04035_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09252_ (.A1(_01131_),
    .A2(_04033_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09253_ (.A1(_04029_),
    .A2(_04499_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place502 (.I(_02704_),
    .Z(net502));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place549 (.I(net13),
    .Z(net549));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09256_ (.I0(\dp.rf.rf[11][0] ),
    .I1(net478),
    .S(_04500_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09257_ (.I0(\dp.rf.rf[11][10] ),
    .I1(_04069_),
    .S(_04500_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09258_ (.I0(\dp.rf.rf[11][11] ),
    .I1(_04092_),
    .S(_04500_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09259_ (.I0(\dp.rf.rf[11][12] ),
    .I1(_04106_),
    .S(_04500_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09260_ (.I0(\dp.rf.rf[11][13] ),
    .I1(_04119_),
    .S(_04500_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09261_ (.I0(\dp.rf.rf[11][14] ),
    .I1(_04136_),
    .S(_04500_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09262_ (.I0(\dp.rf.rf[11][15] ),
    .I1(_04152_),
    .S(_04500_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place501 (.I(_02787_),
    .Z(net501));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place495 (.I(_04611_),
    .Z(net495));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09265_ (.A1(_04029_),
    .A2(_04499_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place494 (.I(_04626_),
    .Z(net494));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09267_ (.A1(\dp.rf.rf[11][16] ),
    .A2(_04505_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09268_ (.A1(_04178_),
    .A2(_04505_),
    .B(_04507_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09269_ (.I0(\dp.rf.rf[11][17] ),
    .I1(net483),
    .S(_04500_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09270_ (.I0(\dp.rf.rf[11][18] ),
    .I1(net482),
    .S(_04500_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09271_ (.I0(\dp.rf.rf[11][19] ),
    .I1(_04222_),
    .S(_04500_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place493 (.I(_04641_),
    .Z(net493));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09273_ (.I0(\dp.rf.rf[11][1] ),
    .I1(_04228_),
    .S(_04500_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place492 (.I(_04656_),
    .Z(net492));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09275_ (.A1(\dp.rf.rf[11][20] ),
    .A2(_04505_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09276_ (.A1(_04250_),
    .A2(_04505_),
    .B(_04510_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09277_ (.I0(\dp.rf.rf[11][21] ),
    .I1(_04267_),
    .S(_04500_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09278_ (.I0(\dp.rf.rf[11][22] ),
    .I1(net481),
    .S(_04500_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09279_ (.I(\dp.rf.rf[11][23] ),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place491 (.I(_04984_),
    .Z(net491));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09281_ (.A1(_04301_),
    .A2(_04500_),
    .Z(_04513_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09282_ (.A1(_04511_),
    .A2(_04505_),
    .B1(_04513_),
    .B2(net485),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09283_ (.I0(\dp.rf.rf[11][24] ),
    .I1(_04314_),
    .S(_04500_),
    .Z(_00083_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09284_ (.I(\dp.rf.rf[11][25] ),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place496 (.I(_02909_),
    .Z(net496));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place498 (.I(_02907_),
    .Z(net498));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09287_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04500_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09288_ (.A1(_04514_),
    .A2(_04505_),
    .B1(_04517_),
    .B2(_04325_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09289_ (.I0(\dp.rf.rf[11][26] ),
    .I1(_04343_),
    .S(_04500_),
    .Z(_00085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09290_ (.I0(\dp.rf.rf[11][27] ),
    .I1(_04355_),
    .S(_04500_),
    .Z(_00086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09291_ (.I0(\dp.rf.rf[11][28] ),
    .I1(_04370_),
    .S(_04500_),
    .Z(_00087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09292_ (.I(\dp.rf.rf[11][29] ),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place499 (.I(_02896_),
    .Z(net499));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place500 (.I(_02859_),
    .Z(net500));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09295_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04500_),
    .Z(_04521_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09296_ (.A1(_04518_),
    .A2(_04505_),
    .B1(_04521_),
    .B2(net480),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09297_ (.I0(\dp.rf.rf[11][2] ),
    .I1(_04396_),
    .S(_04500_),
    .Z(_00089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09298_ (.I0(\dp.rf.rf[11][30] ),
    .I1(net477),
    .S(_04500_),
    .Z(_00090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09299_ (.I(\dp.rf.rf[11][31] ),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place547 (.I(net13),
    .Z(net547));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09301_ (.A1(_04429_),
    .A2(_04500_),
    .Z(_04524_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09302_ (.A1(_04522_),
    .A2(_04505_),
    .B1(_04524_),
    .B2(net479),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09303_ (.I0(\dp.rf.rf[11][3] ),
    .I1(_04436_),
    .S(_04500_),
    .Z(_00092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09304_ (.I0(\dp.rf.rf[11][4] ),
    .I1(_04446_),
    .S(_04500_),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09305_ (.I0(\dp.rf.rf[11][5] ),
    .I1(_04455_),
    .S(_04500_),
    .Z(_00094_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place517 (.I(_01216_),
    .Z(net517));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09307_ (.A1(\dp.rf.rf[11][6] ),
    .A2(_04505_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09308_ (.A1(_04466_),
    .A2(_04505_),
    .B(_04526_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09309_ (.I0(\dp.rf.rf[11][7] ),
    .I1(_04473_),
    .S(_04500_),
    .Z(_00096_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place488 (.I(_05027_),
    .Z(net488));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09311_ (.A1(\dp.rf.rf[11][8] ),
    .A2(_04505_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09312_ (.A1(_04485_),
    .A2(_04505_),
    .B(_04528_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09313_ (.I0(\dp.rf.rf[11][9] ),
    .I1(_04497_),
    .S(_04500_),
    .Z(_00098_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _09314_ (.A1(_02684_),
    .A2(net2),
    .A3(net32),
    .Z(_04529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09315_ (.A1(_02831_),
    .A2(_04032_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09316_ (.I(net2),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09317_ (.A1(_04531_),
    .A2(_04028_),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _09318_ (.A1(net30),
    .A2(_04530_),
    .A3(_04532_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09319_ (.A1(_04529_),
    .A2(_04533_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place477 (.I(_04412_),
    .Z(net477));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place482 (.I(_04213_),
    .Z(net482));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09322_ (.I0(\dp.rf.rf[12][0] ),
    .I1(net478),
    .S(_04534_),
    .Z(_00099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09323_ (.I0(\dp.rf.rf[12][10] ),
    .I1(_04069_),
    .S(_04534_),
    .Z(_00100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09324_ (.I0(\dp.rf.rf[12][11] ),
    .I1(_04092_),
    .S(_04534_),
    .Z(_00101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09325_ (.I0(\dp.rf.rf[12][12] ),
    .I1(_04106_),
    .S(_04534_),
    .Z(_00102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09326_ (.I0(\dp.rf.rf[12][13] ),
    .I1(_04119_),
    .S(_04534_),
    .Z(_00103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09327_ (.I0(\dp.rf.rf[12][14] ),
    .I1(_04136_),
    .S(_04534_),
    .Z(_00104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09328_ (.I0(\dp.rf.rf[12][15] ),
    .I1(_04152_),
    .S(_04534_),
    .Z(_00105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09329_ (.A1(_04529_),
    .A2(_04533_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_26_clk (.I(clknet_6_10__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09331_ (.A1(\dp.rf.rf[12][16] ),
    .A2(_04537_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09332_ (.A1(_04178_),
    .A2(_04537_),
    .B(_04539_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09333_ (.I0(\dp.rf.rf[12][17] ),
    .I1(net483),
    .S(_04534_),
    .Z(_00107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09334_ (.I0(\dp.rf.rf[12][18] ),
    .I1(net482),
    .S(_04534_),
    .Z(_00108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09335_ (.I0(\dp.rf.rf[12][19] ),
    .I1(_04222_),
    .S(_04534_),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place497 (.I(_02907_),
    .Z(net497));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09337_ (.I0(\dp.rf.rf[12][1] ),
    .I1(_04228_),
    .S(_04534_),
    .Z(_00110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09338_ (.A1(\dp.rf.rf[12][20] ),
    .A2(_04537_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09339_ (.A1(_04250_),
    .A2(_04537_),
    .B(_04541_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09340_ (.I0(\dp.rf.rf[12][21] ),
    .I1(_04267_),
    .S(_04534_),
    .Z(_00112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09341_ (.I0(\dp.rf.rf[12][22] ),
    .I1(net481),
    .S(_04534_),
    .Z(_00113_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09342_ (.I(\dp.rf.rf[12][23] ),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09343_ (.A1(_04301_),
    .A2(_04534_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09344_ (.A1(_04542_),
    .A2(_04537_),
    .B1(_04543_),
    .B2(net485),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09345_ (.I0(\dp.rf.rf[12][24] ),
    .I1(_04314_),
    .S(_04534_),
    .Z(_00115_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09346_ (.I(\dp.rf.rf[12][25] ),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09347_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04534_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09348_ (.A1(_04544_),
    .A2(_04537_),
    .B1(_04545_),
    .B2(_04325_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09349_ (.I0(\dp.rf.rf[12][26] ),
    .I1(_04343_),
    .S(_04534_),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09350_ (.I0(\dp.rf.rf[12][27] ),
    .I1(_04355_),
    .S(_04534_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09351_ (.I0(\dp.rf.rf[12][28] ),
    .I1(_04370_),
    .S(_04534_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09352_ (.I(\dp.rf.rf[12][29] ),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09353_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04534_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09354_ (.A1(_04546_),
    .A2(_04537_),
    .B1(_04547_),
    .B2(net480),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09355_ (.I0(\dp.rf.rf[12][2] ),
    .I1(_04396_),
    .S(_04534_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09356_ (.I0(\dp.rf.rf[12][30] ),
    .I1(net477),
    .S(_04534_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09357_ (.I(\dp.rf.rf[12][31] ),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09358_ (.A1(_04429_),
    .A2(_04534_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09359_ (.A1(_04548_),
    .A2(_04537_),
    .B1(_04549_),
    .B2(net479),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09360_ (.I0(\dp.rf.rf[12][3] ),
    .I1(_04436_),
    .S(_04534_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09361_ (.I0(\dp.rf.rf[12][4] ),
    .I1(_04446_),
    .S(_04534_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09362_ (.I0(\dp.rf.rf[12][5] ),
    .I1(_04455_),
    .S(_04534_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09363_ (.A1(\dp.rf.rf[12][6] ),
    .A2(_04537_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09364_ (.A1(_04466_),
    .A2(_04537_),
    .B(_04550_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09365_ (.I0(\dp.rf.rf[12][7] ),
    .I1(_04473_),
    .S(_04534_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09366_ (.A1(\dp.rf.rf[12][8] ),
    .A2(_04537_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09367_ (.A1(_04485_),
    .A2(_04537_),
    .B(_04551_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09368_ (.I0(\dp.rf.rf[12][9] ),
    .I1(_04497_),
    .S(_04534_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09369_ (.A1(_01131_),
    .A2(_04530_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_27_clk (.I(clknet_6_10__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09371_ (.A1(_04529_),
    .A2(_04552_),
    .Z(_04554_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_28_clk (.I(clknet_6_10__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_42_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09374_ (.I0(\dp.rf.rf[13][0] ),
    .I1(net478),
    .S(_04554_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09375_ (.I0(\dp.rf.rf[13][10] ),
    .I1(_04069_),
    .S(_04554_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09376_ (.I0(\dp.rf.rf[13][11] ),
    .I1(_04092_),
    .S(_04554_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09377_ (.I0(\dp.rf.rf[13][12] ),
    .I1(_04106_),
    .S(_04554_),
    .Z(_00134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09378_ (.I0(\dp.rf.rf[13][13] ),
    .I1(_04119_),
    .S(_04554_),
    .Z(_00135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09379_ (.I0(\dp.rf.rf[13][14] ),
    .I1(_04136_),
    .S(_04554_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09380_ (.I0(\dp.rf.rf[13][15] ),
    .I1(_04152_),
    .S(_04554_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09381_ (.A1(_04529_),
    .A2(_04552_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_56_clk (.I(clknet_6_40__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09383_ (.A1(\dp.rf.rf[13][16] ),
    .A2(_04557_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09384_ (.A1(_04178_),
    .A2(_04557_),
    .B(_04559_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09385_ (.I0(\dp.rf.rf[13][17] ),
    .I1(net483),
    .S(_04554_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09386_ (.I0(\dp.rf.rf[13][18] ),
    .I1(net482),
    .S(_04554_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09387_ (.I0(\dp.rf.rf[13][19] ),
    .I1(_04222_),
    .S(_04554_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place546 (.I(net14),
    .Z(net546));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09389_ (.I0(\dp.rf.rf[13][1] ),
    .I1(_04228_),
    .S(_04554_),
    .Z(_00142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09390_ (.A1(\dp.rf.rf[13][20] ),
    .A2(_04557_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09391_ (.A1(_04250_),
    .A2(_04557_),
    .B(_04561_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09392_ (.I0(\dp.rf.rf[13][21] ),
    .I1(_04267_),
    .S(_04554_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09393_ (.I0(\dp.rf.rf[13][22] ),
    .I1(net481),
    .S(_04554_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09394_ (.I(\dp.rf.rf[13][23] ),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09395_ (.A1(_04301_),
    .A2(_04554_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09396_ (.A1(_04562_),
    .A2(_04557_),
    .B1(_04563_),
    .B2(net485),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09397_ (.I0(\dp.rf.rf[13][24] ),
    .I1(_04314_),
    .S(_04554_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09398_ (.I(\dp.rf.rf[13][25] ),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09399_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04554_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09400_ (.A1(_04564_),
    .A2(_04557_),
    .B1(_04565_),
    .B2(_04325_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09401_ (.I0(\dp.rf.rf[13][26] ),
    .I1(_04343_),
    .S(_04554_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09402_ (.I0(\dp.rf.rf[13][27] ),
    .I1(_04355_),
    .S(_04554_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09403_ (.I0(\dp.rf.rf[13][28] ),
    .I1(_04370_),
    .S(_04554_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09404_ (.I(\dp.rf.rf[13][29] ),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09405_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04554_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09406_ (.A1(_04566_),
    .A2(_04557_),
    .B1(_04567_),
    .B2(net480),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09407_ (.I0(\dp.rf.rf[13][2] ),
    .I1(_04396_),
    .S(_04554_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09408_ (.I0(\dp.rf.rf[13][30] ),
    .I1(net477),
    .S(_04554_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09409_ (.I(\dp.rf.rf[13][31] ),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09410_ (.A1(_04429_),
    .A2(_04554_),
    .Z(_04569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09411_ (.A1(_04568_),
    .A2(_04557_),
    .B1(_04569_),
    .B2(net479),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09412_ (.I0(\dp.rf.rf[13][3] ),
    .I1(_04436_),
    .S(_04554_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09413_ (.I0(\dp.rf.rf[13][4] ),
    .I1(_04446_),
    .S(_04554_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09414_ (.I0(\dp.rf.rf[13][5] ),
    .I1(_04455_),
    .S(_04554_),
    .Z(_00158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09415_ (.A1(\dp.rf.rf[13][6] ),
    .A2(_04557_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09416_ (.A1(_04466_),
    .A2(_04557_),
    .B(_04570_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09417_ (.I0(\dp.rf.rf[13][7] ),
    .I1(_04473_),
    .S(_04554_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09418_ (.A1(\dp.rf.rf[13][8] ),
    .A2(_04557_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09419_ (.A1(_04485_),
    .A2(_04557_),
    .B(_04571_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09420_ (.I0(\dp.rf.rf[13][9] ),
    .I1(_04497_),
    .S(_04554_),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09421_ (.A1(_04034_),
    .A2(_04529_),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_58_clk (.I(clknet_6_40__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place487 (.I(_04013_),
    .Z(net487));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09424_ (.I0(\dp.rf.rf[14][0] ),
    .I1(net478),
    .S(_04572_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09425_ (.I0(\dp.rf.rf[14][10] ),
    .I1(_04069_),
    .S(_04572_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09426_ (.I0(\dp.rf.rf[14][11] ),
    .I1(_04092_),
    .S(_04572_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09427_ (.I0(\dp.rf.rf[14][12] ),
    .I1(_04106_),
    .S(_04572_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09428_ (.I0(\dp.rf.rf[14][13] ),
    .I1(_04119_),
    .S(_04572_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09429_ (.I0(\dp.rf.rf[14][14] ),
    .I1(_04136_),
    .S(_04572_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09430_ (.I0(\dp.rf.rf[14][15] ),
    .I1(_04152_),
    .S(_04572_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09431_ (.A1(_04034_),
    .A2(_04529_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_60_clk (.I(clknet_6_40__leaf_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09433_ (.A1(\dp.rf.rf[14][16] ),
    .A2(_04575_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09434_ (.A1(_04178_),
    .A2(_04575_),
    .B(_04577_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09435_ (.I0(\dp.rf.rf[14][17] ),
    .I1(net483),
    .S(_04572_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09436_ (.I0(\dp.rf.rf[14][18] ),
    .I1(net482),
    .S(_04572_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09437_ (.I0(\dp.rf.rf[14][19] ),
    .I1(_04222_),
    .S(_04572_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_64_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09439_ (.I0(\dp.rf.rf[14][1] ),
    .I1(_04228_),
    .S(_04572_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09440_ (.A1(\dp.rf.rf[14][20] ),
    .A2(_04575_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09441_ (.A1(_04250_),
    .A2(_04575_),
    .B(_04579_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09442_ (.I0(\dp.rf.rf[14][21] ),
    .I1(_04267_),
    .S(_04572_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09443_ (.I0(\dp.rf.rf[14][22] ),
    .I1(net481),
    .S(_04572_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09444_ (.I(\dp.rf.rf[14][23] ),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09445_ (.A1(_04301_),
    .A2(_04572_),
    .Z(_04581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09446_ (.A1(_04580_),
    .A2(_04575_),
    .B1(_04581_),
    .B2(net485),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09447_ (.I0(\dp.rf.rf[14][24] ),
    .I1(_04314_),
    .S(_04572_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09448_ (.I(\dp.rf.rf[14][25] ),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09449_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04572_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09450_ (.A1(_04582_),
    .A2(_04575_),
    .B1(_04583_),
    .B2(_04325_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09451_ (.I0(\dp.rf.rf[14][26] ),
    .I1(_04343_),
    .S(_04572_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09452_ (.I0(\dp.rf.rf[14][27] ),
    .I1(_04355_),
    .S(_04572_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09453_ (.I0(\dp.rf.rf[14][28] ),
    .I1(_04370_),
    .S(_04572_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09454_ (.I(\dp.rf.rf[14][29] ),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09455_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04572_),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09456_ (.A1(_04584_),
    .A2(_04575_),
    .B1(_04585_),
    .B2(net480),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09457_ (.I0(\dp.rf.rf[14][2] ),
    .I1(_04396_),
    .S(_04572_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09458_ (.I0(\dp.rf.rf[14][30] ),
    .I1(net477),
    .S(_04572_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09459_ (.I(\dp.rf.rf[14][31] ),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09460_ (.A1(_04429_),
    .A2(_04572_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09461_ (.A1(_04586_),
    .A2(_04575_),
    .B1(_04587_),
    .B2(net479),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09462_ (.I0(\dp.rf.rf[14][3] ),
    .I1(_04436_),
    .S(_04572_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09463_ (.I0(\dp.rf.rf[14][4] ),
    .I1(_04446_),
    .S(_04572_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09464_ (.I0(\dp.rf.rf[14][5] ),
    .I1(_04455_),
    .S(_04572_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09465_ (.A1(\dp.rf.rf[14][6] ),
    .A2(_04575_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09466_ (.A1(_04466_),
    .A2(_04575_),
    .B(_04588_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09467_ (.I0(\dp.rf.rf[14][7] ),
    .I1(_04473_),
    .S(_04572_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09468_ (.A1(\dp.rf.rf[14][8] ),
    .A2(_04575_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09469_ (.A1(_04485_),
    .A2(_04575_),
    .B(_04589_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09470_ (.I0(\dp.rf.rf[14][9] ),
    .I1(_04497_),
    .S(_04572_),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09471_ (.A1(_04499_),
    .A2(_04529_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place485 (.I(_04297_),
    .Z(net485));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_65_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09474_ (.I0(\dp.rf.rf[15][0] ),
    .I1(net478),
    .S(_04590_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09475_ (.I0(\dp.rf.rf[15][10] ),
    .I1(_04069_),
    .S(_04590_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09476_ (.I0(\dp.rf.rf[15][11] ),
    .I1(_04092_),
    .S(_04590_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09477_ (.I0(\dp.rf.rf[15][12] ),
    .I1(_04106_),
    .S(_04590_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09478_ (.I0(\dp.rf.rf[15][13] ),
    .I1(_04119_),
    .S(_04590_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09479_ (.I0(\dp.rf.rf[15][14] ),
    .I1(_04136_),
    .S(_04590_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09480_ (.I0(\dp.rf.rf[15][15] ),
    .I1(_04152_),
    .S(_04590_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09481_ (.A1(_04499_),
    .A2(_04529_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_67_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09483_ (.A1(\dp.rf.rf[15][16] ),
    .A2(_04593_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09484_ (.A1(_04178_),
    .A2(_04593_),
    .B(_04595_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09485_ (.I0(\dp.rf.rf[15][17] ),
    .I1(net483),
    .S(_04590_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09486_ (.I0(\dp.rf.rf[15][18] ),
    .I1(net482),
    .S(_04590_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09487_ (.I0(\dp.rf.rf[15][19] ),
    .I1(_04222_),
    .S(_04590_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_68_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09489_ (.I0(\dp.rf.rf[15][1] ),
    .I1(_04228_),
    .S(_04590_),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09490_ (.A1(\dp.rf.rf[15][20] ),
    .A2(_04593_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09491_ (.A1(_04250_),
    .A2(_04593_),
    .B(_04597_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09492_ (.I0(\dp.rf.rf[15][21] ),
    .I1(_04267_),
    .S(_04590_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09493_ (.I0(\dp.rf.rf[15][22] ),
    .I1(net481),
    .S(_04590_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09494_ (.I(\dp.rf.rf[15][23] ),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09495_ (.A1(_04301_),
    .A2(_04590_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09496_ (.A1(_04598_),
    .A2(_04593_),
    .B1(_04599_),
    .B2(net485),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09497_ (.I0(\dp.rf.rf[15][24] ),
    .I1(_04314_),
    .S(_04590_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09498_ (.I(\dp.rf.rf[15][25] ),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09499_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04590_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09500_ (.A1(_04600_),
    .A2(_04593_),
    .B1(_04601_),
    .B2(_04325_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09501_ (.I0(\dp.rf.rf[15][26] ),
    .I1(_04343_),
    .S(_04590_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09502_ (.I0(\dp.rf.rf[15][27] ),
    .I1(_04355_),
    .S(_04590_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09503_ (.I0(\dp.rf.rf[15][28] ),
    .I1(_04370_),
    .S(_04590_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09504_ (.I(\dp.rf.rf[15][29] ),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09505_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04590_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09506_ (.A1(_04602_),
    .A2(_04593_),
    .B1(_04603_),
    .B2(net480),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09507_ (.I0(\dp.rf.rf[15][2] ),
    .I1(_04396_),
    .S(_04590_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09508_ (.I0(\dp.rf.rf[15][30] ),
    .I1(net477),
    .S(_04590_),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09509_ (.I(\dp.rf.rf[15][31] ),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09510_ (.A1(_04429_),
    .A2(_04590_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09511_ (.A1(_04604_),
    .A2(_04593_),
    .B1(_04605_),
    .B2(net479),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09512_ (.I0(\dp.rf.rf[15][3] ),
    .I1(_04436_),
    .S(_04590_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09513_ (.I0(\dp.rf.rf[15][4] ),
    .I1(_04446_),
    .S(_04590_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09514_ (.I0(\dp.rf.rf[15][5] ),
    .I1(_04455_),
    .S(_04590_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09515_ (.A1(\dp.rf.rf[15][6] ),
    .A2(_04593_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09516_ (.A1(_04466_),
    .A2(_04593_),
    .B(_04606_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09517_ (.I0(\dp.rf.rf[15][7] ),
    .I1(_04473_),
    .S(_04590_),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09518_ (.A1(\dp.rf.rf[15][8] ),
    .A2(_04593_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09519_ (.A1(_04485_),
    .A2(_04593_),
    .B(_04607_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09520_ (.I0(\dp.rf.rf[15][9] ),
    .I1(_04497_),
    .S(_04590_),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09521_ (.A1(net30),
    .A2(_04530_),
    .A3(_04532_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _09522_ (.A1(_02684_),
    .A2(net2),
    .A3(net32),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_73_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09524_ (.A1(_04608_),
    .A2(_04609_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_74_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09526_ (.I0(\dp.rf.rf[16][0] ),
    .I1(net478),
    .S(net495),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09527_ (.I0(\dp.rf.rf[16][10] ),
    .I1(_04069_),
    .S(net495),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09528_ (.I0(\dp.rf.rf[16][11] ),
    .I1(_04092_),
    .S(net495),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09529_ (.I0(\dp.rf.rf[16][12] ),
    .I1(_04106_),
    .S(net495),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09530_ (.I0(\dp.rf.rf[16][13] ),
    .I1(_04119_),
    .S(net495),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09531_ (.I0(\dp.rf.rf[16][14] ),
    .I1(_04136_),
    .S(net495),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09532_ (.I0(\dp.rf.rf[16][15] ),
    .I1(_04152_),
    .S(net495),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09533_ (.A1(_04608_),
    .A2(_04609_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_75_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09535_ (.A1(\dp.rf.rf[16][16] ),
    .A2(_04613_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09536_ (.A1(_04178_),
    .A2(_04613_),
    .B(_04615_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09537_ (.I0(\dp.rf.rf[16][17] ),
    .I1(net483),
    .S(net495),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09538_ (.I0(\dp.rf.rf[16][18] ),
    .I1(net482),
    .S(net495),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09539_ (.I0(\dp.rf.rf[16][19] ),
    .I1(_04222_),
    .S(net495),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_76_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09541_ (.I0(\dp.rf.rf[16][1] ),
    .I1(_04228_),
    .S(_04611_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09542_ (.A1(\dp.rf.rf[16][20] ),
    .A2(_04613_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09543_ (.A1(_04250_),
    .A2(_04613_),
    .B(_04617_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09544_ (.I0(\dp.rf.rf[16][21] ),
    .I1(_04267_),
    .S(_04611_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09545_ (.I0(\dp.rf.rf[16][22] ),
    .I1(net481),
    .S(_04611_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09546_ (.A1(_04301_),
    .A2(_04611_),
    .Z(_04618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09547_ (.A1(_01795_),
    .A2(_04613_),
    .B1(_04618_),
    .B2(net485),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09548_ (.I0(\dp.rf.rf[16][24] ),
    .I1(_04314_),
    .S(_04611_),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09549_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04611_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09550_ (.A1(_01674_),
    .A2(_04613_),
    .B1(_04619_),
    .B2(_04325_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09551_ (.I0(\dp.rf.rf[16][26] ),
    .I1(_04343_),
    .S(_04611_),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09552_ (.I0(\dp.rf.rf[16][27] ),
    .I1(_04355_),
    .S(_04611_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09553_ (.I0(\dp.rf.rf[16][28] ),
    .I1(_04370_),
    .S(_04611_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09554_ (.I(\dp.rf.rf[16][29] ),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09555_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04611_),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09556_ (.A1(_04620_),
    .A2(_04613_),
    .B1(_04621_),
    .B2(net480),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09557_ (.I0(\dp.rf.rf[16][2] ),
    .I1(_04396_),
    .S(_04611_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09558_ (.I0(\dp.rf.rf[16][30] ),
    .I1(net477),
    .S(_04611_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09559_ (.A1(_04429_),
    .A2(net495),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09560_ (.A1(_01258_),
    .A2(_04613_),
    .B1(_04622_),
    .B2(net479),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09561_ (.I0(\dp.rf.rf[16][3] ),
    .I1(_04436_),
    .S(net495),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09562_ (.I0(\dp.rf.rf[16][4] ),
    .I1(_04446_),
    .S(_04611_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09563_ (.I0(\dp.rf.rf[16][5] ),
    .I1(_04455_),
    .S(net495),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09564_ (.A1(\dp.rf.rf[16][6] ),
    .A2(_04613_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09565_ (.A1(_04466_),
    .A2(_04613_),
    .B(_04623_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09566_ (.I0(\dp.rf.rf[16][7] ),
    .I1(_04473_),
    .S(net495),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09567_ (.A1(\dp.rf.rf[16][8] ),
    .A2(_04613_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09568_ (.A1(_04485_),
    .A2(_04613_),
    .B(_04624_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09569_ (.I0(\dp.rf.rf[16][9] ),
    .I1(_04497_),
    .S(_04611_),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09570_ (.A1(_01131_),
    .A2(_04530_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09571_ (.A1(_04625_),
    .A2(_04609_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09573_ (.I0(\dp.rf.rf[17][0] ),
    .I1(net478),
    .S(net494),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09574_ (.I0(\dp.rf.rf[17][10] ),
    .I1(_04069_),
    .S(net494),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09575_ (.I0(\dp.rf.rf[17][11] ),
    .I1(_04092_),
    .S(net494),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09576_ (.I0(\dp.rf.rf[17][12] ),
    .I1(_04106_),
    .S(net494),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09577_ (.I0(\dp.rf.rf[17][13] ),
    .I1(_04119_),
    .S(net494),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09578_ (.I0(\dp.rf.rf[17][14] ),
    .I1(_04136_),
    .S(net494),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09579_ (.I0(\dp.rf.rf[17][15] ),
    .I1(_04152_),
    .S(net494),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09580_ (.A1(_04625_),
    .A2(_04609_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place481 (.I(_04284_),
    .Z(net481));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09582_ (.A1(\dp.rf.rf[17][16] ),
    .A2(_04628_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09583_ (.A1(_04178_),
    .A2(_04628_),
    .B(_04630_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09584_ (.I0(\dp.rf.rf[17][17] ),
    .I1(net483),
    .S(net494),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09585_ (.I0(\dp.rf.rf[17][18] ),
    .I1(net482),
    .S(net494),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09586_ (.I0(\dp.rf.rf[17][19] ),
    .I1(_04222_),
    .S(net494),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_78_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09588_ (.I0(\dp.rf.rf[17][1] ),
    .I1(_04228_),
    .S(_04626_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09589_ (.A1(\dp.rf.rf[17][20] ),
    .A2(_04628_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09590_ (.A1(_04250_),
    .A2(_04628_),
    .B(_04632_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09591_ (.I0(\dp.rf.rf[17][21] ),
    .I1(_04267_),
    .S(_04626_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09592_ (.I0(\dp.rf.rf[17][22] ),
    .I1(net481),
    .S(_04626_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09593_ (.A1(_04301_),
    .A2(_04626_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09594_ (.A1(_01796_),
    .A2(_04628_),
    .B1(_04633_),
    .B2(net485),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09595_ (.I0(\dp.rf.rf[17][24] ),
    .I1(_04314_),
    .S(_04626_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09596_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04626_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09597_ (.A1(_01675_),
    .A2(_04628_),
    .B1(_04634_),
    .B2(_04325_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09598_ (.I0(\dp.rf.rf[17][26] ),
    .I1(_04343_),
    .S(_04626_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09599_ (.I0(\dp.rf.rf[17][27] ),
    .I1(_04355_),
    .S(_04626_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09600_ (.I0(\dp.rf.rf[17][28] ),
    .I1(_04370_),
    .S(_04626_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09601_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04626_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09602_ (.A1(_01470_),
    .A2(_04628_),
    .B1(_04635_),
    .B2(net480),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09603_ (.I0(\dp.rf.rf[17][2] ),
    .I1(_04396_),
    .S(_04626_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09604_ (.I0(\dp.rf.rf[17][30] ),
    .I1(net477),
    .S(_04626_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09605_ (.I(\dp.rf.rf[17][31] ),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09606_ (.A1(_04429_),
    .A2(net494),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09607_ (.A1(_04636_),
    .A2(_04628_),
    .B1(_04637_),
    .B2(net479),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09608_ (.I0(\dp.rf.rf[17][3] ),
    .I1(_04436_),
    .S(net494),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09609_ (.I0(\dp.rf.rf[17][4] ),
    .I1(_04446_),
    .S(_04626_),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09610_ (.I0(\dp.rf.rf[17][5] ),
    .I1(_04455_),
    .S(net494),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09611_ (.A1(\dp.rf.rf[17][6] ),
    .A2(_04628_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09612_ (.A1(_04466_),
    .A2(_04628_),
    .B(_04638_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09613_ (.I0(\dp.rf.rf[17][7] ),
    .I1(_04473_),
    .S(net494),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09614_ (.A1(\dp.rf.rf[17][8] ),
    .A2(_04628_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09615_ (.A1(_04485_),
    .A2(_04628_),
    .B(_04639_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09616_ (.I0(\dp.rf.rf[17][9] ),
    .I1(_04497_),
    .S(_04626_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09617_ (.A1(net30),
    .A2(_04033_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09618_ (.A1(_04640_),
    .A2(_04609_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_25_clk (.I(clknet_6_10__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09620_ (.I0(\dp.rf.rf[18][0] ),
    .I1(net478),
    .S(net493),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09621_ (.I0(\dp.rf.rf[18][10] ),
    .I1(_04069_),
    .S(net493),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09622_ (.I0(\dp.rf.rf[18][11] ),
    .I1(_04092_),
    .S(net493),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09623_ (.I0(\dp.rf.rf[18][12] ),
    .I1(_04106_),
    .S(net493),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09624_ (.I0(\dp.rf.rf[18][13] ),
    .I1(_04119_),
    .S(net493),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09625_ (.I0(\dp.rf.rf[18][14] ),
    .I1(_04136_),
    .S(net493),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09626_ (.I0(\dp.rf.rf[18][15] ),
    .I1(_04152_),
    .S(net493),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09627_ (.A1(_04640_),
    .A2(_04609_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output164 (.I(net164),
    .Z(writedata[9]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09629_ (.A1(\dp.rf.rf[18][16] ),
    .A2(_04643_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09630_ (.A1(_04178_),
    .A2(_04643_),
    .B(_04645_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09631_ (.I0(\dp.rf.rf[18][17] ),
    .I1(net483),
    .S(net493),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09632_ (.I0(\dp.rf.rf[18][18] ),
    .I1(net482),
    .S(net493),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09633_ (.I0(\dp.rf.rf[18][19] ),
    .I1(_04222_),
    .S(net493),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output163 (.I(net163),
    .Z(writedata[8]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09635_ (.I0(\dp.rf.rf[18][1] ),
    .I1(_04228_),
    .S(_04641_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09636_ (.A1(\dp.rf.rf[18][20] ),
    .A2(_04643_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09637_ (.A1(_04250_),
    .A2(_04643_),
    .B(_04647_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09638_ (.I0(\dp.rf.rf[18][21] ),
    .I1(_04267_),
    .S(_04641_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09639_ (.I0(\dp.rf.rf[18][22] ),
    .I1(net481),
    .S(_04641_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09640_ (.A1(_04301_),
    .A2(_04641_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09641_ (.A1(_01797_),
    .A2(_04643_),
    .B1(_04648_),
    .B2(net485),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09642_ (.I0(\dp.rf.rf[18][24] ),
    .I1(_04314_),
    .S(_04641_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09643_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04641_),
    .Z(_04649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09644_ (.A1(_01676_),
    .A2(_04643_),
    .B1(_04649_),
    .B2(_04325_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09645_ (.I0(\dp.rf.rf[18][26] ),
    .I1(_04343_),
    .S(_04641_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09646_ (.I0(\dp.rf.rf[18][27] ),
    .I1(_04355_),
    .S(_04641_),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09647_ (.I0(\dp.rf.rf[18][28] ),
    .I1(_04370_),
    .S(_04641_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09648_ (.I(\dp.rf.rf[18][29] ),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09649_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04641_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09650_ (.A1(_04650_),
    .A2(_04643_),
    .B1(_04651_),
    .B2(net480),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09651_ (.I0(\dp.rf.rf[18][2] ),
    .I1(_04396_),
    .S(_04641_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09652_ (.I0(\dp.rf.rf[18][30] ),
    .I1(net477),
    .S(_04641_),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09653_ (.A1(_04429_),
    .A2(net493),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09654_ (.A1(_01255_),
    .A2(_04643_),
    .B1(_04652_),
    .B2(net479),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09655_ (.I0(\dp.rf.rf[18][3] ),
    .I1(_04436_),
    .S(net493),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09656_ (.I0(\dp.rf.rf[18][4] ),
    .I1(_04446_),
    .S(_04641_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09657_ (.I0(\dp.rf.rf[18][5] ),
    .I1(_04455_),
    .S(net493),
    .Z(_00318_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09658_ (.A1(\dp.rf.rf[18][6] ),
    .A2(_04643_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09659_ (.A1(_04466_),
    .A2(_04643_),
    .B(_04653_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09660_ (.I0(\dp.rf.rf[18][7] ),
    .I1(_04473_),
    .S(net493),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09661_ (.A1(\dp.rf.rf[18][8] ),
    .A2(_04643_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09662_ (.A1(_04485_),
    .A2(_04643_),
    .B(_04654_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09663_ (.I0(\dp.rf.rf[18][9] ),
    .I1(_04497_),
    .S(_04641_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09664_ (.A1(_01131_),
    .A2(_04033_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _09665_ (.A1(_04655_),
    .A2(_04609_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output162 (.I(net162),
    .Z(writedata[7]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09667_ (.I0(\dp.rf.rf[19][0] ),
    .I1(net478),
    .S(net492),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09668_ (.I0(\dp.rf.rf[19][10] ),
    .I1(_04069_),
    .S(net492),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09669_ (.I0(\dp.rf.rf[19][11] ),
    .I1(_04092_),
    .S(net492),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09670_ (.I0(\dp.rf.rf[19][12] ),
    .I1(_04106_),
    .S(net492),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09671_ (.I0(\dp.rf.rf[19][13] ),
    .I1(_04119_),
    .S(net492),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09672_ (.I0(\dp.rf.rf[19][14] ),
    .I1(_04136_),
    .S(net492),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09673_ (.I0(\dp.rf.rf[19][15] ),
    .I1(_04152_),
    .S(net492),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _09674_ (.A1(_04655_),
    .A2(_04609_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output161 (.I(net161),
    .Z(writedata[6]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09676_ (.A1(\dp.rf.rf[19][16] ),
    .A2(_04658_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09677_ (.A1(_04178_),
    .A2(_04658_),
    .B(_04660_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09678_ (.I0(\dp.rf.rf[19][17] ),
    .I1(net483),
    .S(net492),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09679_ (.I0(\dp.rf.rf[19][18] ),
    .I1(net482),
    .S(net492),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09680_ (.I0(\dp.rf.rf[19][19] ),
    .I1(_04222_),
    .S(net492),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output160 (.I(net160),
    .Z(writedata[5]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09682_ (.I0(\dp.rf.rf[19][1] ),
    .I1(_04228_),
    .S(_04656_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09683_ (.A1(\dp.rf.rf[19][20] ),
    .A2(_04658_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09684_ (.A1(_04250_),
    .A2(_04658_),
    .B(_04662_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09685_ (.I0(\dp.rf.rf[19][21] ),
    .I1(_04267_),
    .S(_04656_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09686_ (.I0(\dp.rf.rf[19][22] ),
    .I1(net481),
    .S(_04656_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09687_ (.A1(_04301_),
    .A2(_04656_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09688_ (.A1(_01798_),
    .A2(_04658_),
    .B1(_04663_),
    .B2(net485),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09689_ (.I0(\dp.rf.rf[19][24] ),
    .I1(_04314_),
    .S(_04656_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09690_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04656_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09691_ (.A1(_01677_),
    .A2(_04658_),
    .B1(_04664_),
    .B2(_04325_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09692_ (.I0(\dp.rf.rf[19][26] ),
    .I1(_04343_),
    .S(_04656_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09693_ (.I0(\dp.rf.rf[19][27] ),
    .I1(_04355_),
    .S(_04656_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09694_ (.I0(\dp.rf.rf[19][28] ),
    .I1(_04370_),
    .S(_04656_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09695_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04656_),
    .Z(_04665_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09696_ (.A1(_01464_),
    .A2(_04658_),
    .B1(_04665_),
    .B2(net480),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09697_ (.I0(\dp.rf.rf[19][2] ),
    .I1(_04396_),
    .S(_04656_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09698_ (.I0(\dp.rf.rf[19][30] ),
    .I1(net477),
    .S(_04656_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09699_ (.I(\dp.rf.rf[19][31] ),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09700_ (.A1(_04429_),
    .A2(net492),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09701_ (.A1(_04666_),
    .A2(_04658_),
    .B1(_04667_),
    .B2(net479),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09702_ (.I0(\dp.rf.rf[19][3] ),
    .I1(_04436_),
    .S(net492),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09703_ (.I0(\dp.rf.rf[19][4] ),
    .I1(_04446_),
    .S(_04656_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09704_ (.I0(\dp.rf.rf[19][5] ),
    .I1(_04455_),
    .S(net492),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09705_ (.A1(\dp.rf.rf[19][6] ),
    .A2(_04658_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09706_ (.A1(_04466_),
    .A2(_04658_),
    .B(_04668_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09707_ (.I0(\dp.rf.rf[19][7] ),
    .I1(_04473_),
    .S(net492),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09708_ (.A1(\dp.rf.rf[19][8] ),
    .A2(_04658_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09709_ (.A1(_04485_),
    .A2(_04658_),
    .B(_04669_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09710_ (.I0(\dp.rf.rf[19][9] ),
    .I1(_04497_),
    .S(_04656_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output159 (.I(net159),
    .Z(writedata[4]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09712_ (.A1(_04532_),
    .A2(_04552_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output158 (.I(net158),
    .Z(writedata[3]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output157 (.I(net157),
    .Z(writedata[31]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09715_ (.I0(\dp.rf.rf[1][0] ),
    .I1(net478),
    .S(_04671_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output156 (.I(net156),
    .Z(writedata[30]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09717_ (.I0(\dp.rf.rf[1][10] ),
    .I1(_04069_),
    .S(_04671_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output155 (.I(net155),
    .Z(writedata[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09719_ (.I0(\dp.rf.rf[1][11] ),
    .I1(_04092_),
    .S(_04671_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output154 (.I(net154),
    .Z(writedata[29]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09721_ (.I0(\dp.rf.rf[1][12] ),
    .I1(_04106_),
    .S(_04671_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output153 (.I(net153),
    .Z(writedata[28]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09723_ (.I0(\dp.rf.rf[1][13] ),
    .I1(_04119_),
    .S(_04671_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output152 (.I(net152),
    .Z(writedata[27]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09725_ (.I0(\dp.rf.rf[1][14] ),
    .I1(_04136_),
    .S(_04671_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output151 (.I(net151),
    .Z(writedata[26]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09727_ (.I0(\dp.rf.rf[1][15] ),
    .I1(_04152_),
    .S(_04671_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09728_ (.A1(_04532_),
    .A2(_04552_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output150 (.I(net150),
    .Z(writedata[25]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09730_ (.A1(\dp.rf.rf[1][16] ),
    .A2(_04680_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09731_ (.A1(_04178_),
    .A2(_04680_),
    .B(_04682_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output149 (.I(net149),
    .Z(writedata[24]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09733_ (.I0(\dp.rf.rf[1][17] ),
    .I1(net483),
    .S(_04671_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output148 (.I(net148),
    .Z(writedata[23]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09735_ (.I0(\dp.rf.rf[1][18] ),
    .I1(net482),
    .S(_04671_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output147 (.I(net147),
    .Z(writedata[22]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09737_ (.I0(\dp.rf.rf[1][19] ),
    .I1(_04222_),
    .S(_04671_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output146 (.I(net146),
    .Z(writedata[21]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output145 (.I(net145),
    .Z(writedata[20]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09740_ (.I0(\dp.rf.rf[1][1] ),
    .I1(_04228_),
    .S(_04671_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09741_ (.A1(\dp.rf.rf[1][20] ),
    .A2(_04680_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09742_ (.A1(_04250_),
    .A2(_04680_),
    .B(_04688_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output144 (.I(net144),
    .Z(writedata[1]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09744_ (.I0(\dp.rf.rf[1][21] ),
    .I1(_04267_),
    .S(_04671_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output143 (.I(net143),
    .Z(writedata[19]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09746_ (.I0(\dp.rf.rf[1][22] ),
    .I1(net481),
    .S(_04671_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09747_ (.I(\dp.rf.rf[1][23] ),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09748_ (.A1(_04301_),
    .A2(_04671_),
    .Z(_04692_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output142 (.I(net142),
    .Z(writedata[18]));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09750_ (.A1(_04691_),
    .A2(_04680_),
    .B1(_04692_),
    .B2(net485),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output141 (.I(net141),
    .Z(writedata[17]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09752_ (.I0(\dp.rf.rf[1][24] ),
    .I1(_04314_),
    .S(_04671_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09753_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04671_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output140 (.I(net140),
    .Z(writedata[16]));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09755_ (.A1(_01708_),
    .A2(_04680_),
    .B1(_04695_),
    .B2(_04325_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output139 (.I(net139),
    .Z(writedata[15]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09757_ (.I0(\dp.rf.rf[1][26] ),
    .I1(_04343_),
    .S(_04671_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output138 (.I(net138),
    .Z(writedata[14]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09759_ (.I0(\dp.rf.rf[1][27] ),
    .I1(_04355_),
    .S(_04671_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output137 (.I(net137),
    .Z(writedata[13]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09761_ (.I0(\dp.rf.rf[1][28] ),
    .I1(_04370_),
    .S(_04671_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09762_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04671_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output136 (.I(net136),
    .Z(writedata[12]));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09764_ (.A1(_01452_),
    .A2(_04680_),
    .B1(_04700_),
    .B2(net480),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output135 (.I(net135),
    .Z(writedata[11]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09766_ (.I0(\dp.rf.rf[1][2] ),
    .I1(_04396_),
    .S(_04671_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output134 (.I(net134),
    .Z(writedata[10]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09768_ (.I0(\dp.rf.rf[1][30] ),
    .I1(net477),
    .S(_04671_),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09769_ (.A1(_04429_),
    .A2(_04671_),
    .Z(_04704_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output133 (.I(net133),
    .Z(writedata[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09771_ (.A1(_01246_),
    .A2(_04680_),
    .B1(_04704_),
    .B2(net479),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output132 (.I(net132),
    .Z(suspend));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09773_ (.I0(\dp.rf.rf[1][3] ),
    .I1(_04436_),
    .S(_04671_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output131 (.I(net131),
    .Z(pc[9]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09775_ (.I0(\dp.rf.rf[1][4] ),
    .I1(_04446_),
    .S(_04671_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output130 (.I(net130),
    .Z(pc[8]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09777_ (.I0(\dp.rf.rf[1][5] ),
    .I1(_04455_),
    .S(_04671_),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09778_ (.A1(\dp.rf.rf[1][6] ),
    .A2(_04680_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09779_ (.A1(_04466_),
    .A2(_04680_),
    .B(_04709_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output129 (.I(net129),
    .Z(pc[7]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09781_ (.I0(\dp.rf.rf[1][7] ),
    .I1(_04473_),
    .S(_04671_),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09782_ (.A1(\dp.rf.rf[1][8] ),
    .A2(_04680_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09783_ (.A1(_04485_),
    .A2(_04680_),
    .B(_04711_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output128 (.I(net128),
    .Z(pc[6]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09785_ (.I0(\dp.rf.rf[1][9] ),
    .I1(_04497_),
    .S(_04671_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _09786_ (.A1(net3),
    .A2(_04531_),
    .A3(net32),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09787_ (.A1(_04533_),
    .A2(_04713_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output127 (.I(net127),
    .Z(pc[5]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output126 (.I(net126),
    .Z(pc[4]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09790_ (.I0(\dp.rf.rf[20][0] ),
    .I1(net478),
    .S(_04714_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09791_ (.I0(\dp.rf.rf[20][10] ),
    .I1(_04069_),
    .S(_04714_),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09792_ (.I0(\dp.rf.rf[20][11] ),
    .I1(_04092_),
    .S(_04714_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09793_ (.I0(\dp.rf.rf[20][12] ),
    .I1(_04106_),
    .S(_04714_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09794_ (.I0(\dp.rf.rf[20][13] ),
    .I1(_04119_),
    .S(_04714_),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09795_ (.I0(\dp.rf.rf[20][14] ),
    .I1(_04136_),
    .S(_04714_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09796_ (.I0(\dp.rf.rf[20][15] ),
    .I1(_04152_),
    .S(_04714_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output125 (.I(net125),
    .Z(pc[3]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09798_ (.A1(_04533_),
    .A2(_04713_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output124 (.I(net124),
    .Z(pc[31]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09800_ (.A1(\dp.rf.rf[20][16] ),
    .A2(_04718_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09801_ (.A1(_04178_),
    .A2(_04718_),
    .B(_04720_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09802_ (.I0(\dp.rf.rf[20][17] ),
    .I1(net483),
    .S(_04714_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09803_ (.I0(\dp.rf.rf[20][18] ),
    .I1(net482),
    .S(_04714_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09804_ (.I0(\dp.rf.rf[20][19] ),
    .I1(_04222_),
    .S(_04714_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output123 (.I(net123),
    .Z(pc[30]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09806_ (.I0(\dp.rf.rf[20][1] ),
    .I1(_04228_),
    .S(_04714_),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output122 (.I(net122),
    .Z(pc[2]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09808_ (.A1(\dp.rf.rf[20][20] ),
    .A2(_04718_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09809_ (.A1(_04250_),
    .A2(_04718_),
    .B(_04723_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09810_ (.I0(\dp.rf.rf[20][21] ),
    .I1(_04267_),
    .S(_04714_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09811_ (.I0(\dp.rf.rf[20][22] ),
    .I1(net481),
    .S(_04714_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output121 (.I(net121),
    .Z(pc[29]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09813_ (.A1(_04301_),
    .A2(_04714_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09814_ (.A1(_01805_),
    .A2(_04718_),
    .B1(_04725_),
    .B2(net485),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09815_ (.I0(\dp.rf.rf[20][24] ),
    .I1(_04314_),
    .S(_04714_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output120 (.I(net120),
    .Z(pc[28]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output119 (.I(net119),
    .Z(pc[27]));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09818_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04714_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09819_ (.A1(_01664_),
    .A2(_04718_),
    .B1(_04728_),
    .B2(_04325_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09820_ (.I0(\dp.rf.rf[20][26] ),
    .I1(_04343_),
    .S(_04714_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09821_ (.I0(\dp.rf.rf[20][27] ),
    .I1(_04355_),
    .S(_04714_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09822_ (.I0(\dp.rf.rf[20][28] ),
    .I1(_04370_),
    .S(_04714_),
    .Z(_00407_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output118 (.I(net118),
    .Z(pc[26]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output117 (.I(net117),
    .Z(pc[25]));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09825_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04714_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09826_ (.A1(_01469_),
    .A2(_04718_),
    .B1(_04731_),
    .B2(net480),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09827_ (.I0(\dp.rf.rf[20][2] ),
    .I1(_04396_),
    .S(_04714_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09828_ (.I0(\dp.rf.rf[20][30] ),
    .I1(net477),
    .S(_04714_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output116 (.I(net116),
    .Z(pc[24]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09830_ (.A1(_04429_),
    .A2(_04714_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09831_ (.A1(_01260_),
    .A2(_04718_),
    .B1(_04733_),
    .B2(net479),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09832_ (.I0(\dp.rf.rf[20][3] ),
    .I1(_04436_),
    .S(_04714_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09833_ (.I0(\dp.rf.rf[20][4] ),
    .I1(_04446_),
    .S(_04714_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09834_ (.I0(\dp.rf.rf[20][5] ),
    .I1(_04455_),
    .S(_04714_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output115 (.I(net115),
    .Z(pc[23]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09836_ (.A1(\dp.rf.rf[20][6] ),
    .A2(_04718_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09837_ (.A1(_04466_),
    .A2(_04718_),
    .B(_04735_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09838_ (.I0(\dp.rf.rf[20][7] ),
    .I1(_04473_),
    .S(_04714_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output114 (.I(net114),
    .Z(pc[22]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09840_ (.A1(\dp.rf.rf[20][8] ),
    .A2(_04718_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09841_ (.A1(_04485_),
    .A2(_04718_),
    .B(_04737_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09842_ (.I0(\dp.rf.rf[20][9] ),
    .I1(_04497_),
    .S(_04714_),
    .Z(_00418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09843_ (.A1(_04552_),
    .A2(_04713_),
    .Z(_04738_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output113 (.I(net113),
    .Z(pc[21]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output112 (.I(net112),
    .Z(pc[20]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09846_ (.I0(\dp.rf.rf[21][0] ),
    .I1(net478),
    .S(_04738_),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09847_ (.I0(\dp.rf.rf[21][10] ),
    .I1(_04069_),
    .S(_04738_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09848_ (.I0(\dp.rf.rf[21][11] ),
    .I1(_04092_),
    .S(_04738_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09849_ (.I0(\dp.rf.rf[21][12] ),
    .I1(_04106_),
    .S(_04738_),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09850_ (.I0(\dp.rf.rf[21][13] ),
    .I1(_04119_),
    .S(_04738_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09851_ (.I0(\dp.rf.rf[21][14] ),
    .I1(_04136_),
    .S(_04738_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09852_ (.I0(\dp.rf.rf[21][15] ),
    .I1(_04152_),
    .S(_04738_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09853_ (.A1(_04552_),
    .A2(_04713_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output111 (.I(net111),
    .Z(pc[1]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09855_ (.A1(\dp.rf.rf[21][16] ),
    .A2(_04741_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09856_ (.A1(_04178_),
    .A2(_04741_),
    .B(_04743_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09857_ (.I0(\dp.rf.rf[21][17] ),
    .I1(net483),
    .S(_04738_),
    .Z(_00427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09858_ (.I0(\dp.rf.rf[21][18] ),
    .I1(net482),
    .S(_04738_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09859_ (.I0(\dp.rf.rf[21][19] ),
    .I1(_04222_),
    .S(_04738_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output110 (.I(net110),
    .Z(pc[19]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09861_ (.I0(\dp.rf.rf[21][1] ),
    .I1(_04228_),
    .S(_04738_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09862_ (.A1(\dp.rf.rf[21][20] ),
    .A2(_04741_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09863_ (.A1(_04250_),
    .A2(_04741_),
    .B(_04745_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09864_ (.I0(\dp.rf.rf[21][21] ),
    .I1(_04267_),
    .S(_04738_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09865_ (.I0(\dp.rf.rf[21][22] ),
    .I1(net481),
    .S(_04738_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09866_ (.A1(_04301_),
    .A2(_04738_),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09867_ (.A1(_01806_),
    .A2(_04741_),
    .B1(_04746_),
    .B2(net485),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09868_ (.I0(\dp.rf.rf[21][24] ),
    .I1(_04314_),
    .S(_04738_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09869_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04738_),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09870_ (.A1(_01665_),
    .A2(_04741_),
    .B1(_04747_),
    .B2(_04325_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09871_ (.I0(\dp.rf.rf[21][26] ),
    .I1(_04343_),
    .S(_04738_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09872_ (.I0(\dp.rf.rf[21][27] ),
    .I1(_04355_),
    .S(_04738_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09873_ (.I0(\dp.rf.rf[21][28] ),
    .I1(_04370_),
    .S(_04738_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09874_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04738_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09875_ (.A1(_01471_),
    .A2(_04741_),
    .B1(_04748_),
    .B2(net480),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09876_ (.I0(\dp.rf.rf[21][2] ),
    .I1(_04396_),
    .S(_04738_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09877_ (.I0(\dp.rf.rf[21][30] ),
    .I1(net477),
    .S(_04738_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09878_ (.A1(_04429_),
    .A2(_04738_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09879_ (.A1(_01261_),
    .A2(_04741_),
    .B1(_04749_),
    .B2(net479),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09880_ (.I0(\dp.rf.rf[21][3] ),
    .I1(_04436_),
    .S(_04738_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09881_ (.I0(\dp.rf.rf[21][4] ),
    .I1(_04446_),
    .S(_04738_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09882_ (.I0(\dp.rf.rf[21][5] ),
    .I1(_04455_),
    .S(_04738_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09883_ (.A1(\dp.rf.rf[21][6] ),
    .A2(_04741_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09884_ (.A1(_04466_),
    .A2(_04741_),
    .B(_04750_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09885_ (.I0(\dp.rf.rf[21][7] ),
    .I1(_04473_),
    .S(_04738_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09886_ (.A1(\dp.rf.rf[21][8] ),
    .A2(_04741_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09887_ (.A1(_04485_),
    .A2(_04741_),
    .B(_04751_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09888_ (.I0(\dp.rf.rf[21][9] ),
    .I1(_04497_),
    .S(_04738_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09889_ (.A1(_04034_),
    .A2(_04713_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output109 (.I(net109),
    .Z(pc[18]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output108 (.I(net108),
    .Z(pc[17]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09892_ (.I0(\dp.rf.rf[22][0] ),
    .I1(net478),
    .S(_04752_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09893_ (.I0(\dp.rf.rf[22][10] ),
    .I1(_04069_),
    .S(_04752_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09894_ (.I0(\dp.rf.rf[22][11] ),
    .I1(_04092_),
    .S(_04752_),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09895_ (.I0(\dp.rf.rf[22][12] ),
    .I1(_04106_),
    .S(_04752_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09896_ (.I0(\dp.rf.rf[22][13] ),
    .I1(_04119_),
    .S(_04752_),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09897_ (.I0(\dp.rf.rf[22][14] ),
    .I1(_04136_),
    .S(_04752_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09898_ (.I0(\dp.rf.rf[22][15] ),
    .I1(_04152_),
    .S(_04752_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09899_ (.A1(_04034_),
    .A2(_04713_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output107 (.I(net107),
    .Z(pc[16]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09901_ (.A1(\dp.rf.rf[22][16] ),
    .A2(_04755_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09902_ (.A1(_04178_),
    .A2(_04755_),
    .B(_04757_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09903_ (.I0(\dp.rf.rf[22][17] ),
    .I1(net483),
    .S(_04752_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09904_ (.I0(\dp.rf.rf[22][18] ),
    .I1(net482),
    .S(_04752_),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09905_ (.I0(\dp.rf.rf[22][19] ),
    .I1(_04222_),
    .S(_04752_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output106 (.I(net106),
    .Z(pc[15]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09907_ (.I0(\dp.rf.rf[22][1] ),
    .I1(_04228_),
    .S(_04752_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09908_ (.A1(\dp.rf.rf[22][20] ),
    .A2(_04755_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09909_ (.A1(_04250_),
    .A2(_04755_),
    .B(_04759_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09910_ (.I0(\dp.rf.rf[22][21] ),
    .I1(_04267_),
    .S(_04752_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09911_ (.I0(\dp.rf.rf[22][22] ),
    .I1(net481),
    .S(_04752_),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09912_ (.A1(_04301_),
    .A2(_04752_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09913_ (.A1(_01807_),
    .A2(_04755_),
    .B1(_04760_),
    .B2(net485),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09914_ (.I0(\dp.rf.rf[22][24] ),
    .I1(_04314_),
    .S(_04752_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09915_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04752_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09916_ (.A1(_01666_),
    .A2(_04755_),
    .B1(_04761_),
    .B2(_04325_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09917_ (.I0(\dp.rf.rf[22][26] ),
    .I1(_04343_),
    .S(_04752_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09918_ (.I0(\dp.rf.rf[22][27] ),
    .I1(_04355_),
    .S(_04752_),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09919_ (.I0(\dp.rf.rf[22][28] ),
    .I1(_04370_),
    .S(_04752_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09920_ (.I(\dp.rf.rf[22][29] ),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09921_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04752_),
    .Z(_04763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09922_ (.A1(_04762_),
    .A2(_04755_),
    .B1(_04763_),
    .B2(net480),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09923_ (.I0(\dp.rf.rf[22][2] ),
    .I1(_04396_),
    .S(_04752_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09924_ (.I0(\dp.rf.rf[22][30] ),
    .I1(net477),
    .S(_04752_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09925_ (.A1(_04429_),
    .A2(_04752_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09926_ (.A1(_01262_),
    .A2(_04755_),
    .B1(_04764_),
    .B2(net479),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09927_ (.I0(\dp.rf.rf[22][3] ),
    .I1(_04436_),
    .S(_04752_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09928_ (.I0(\dp.rf.rf[22][4] ),
    .I1(_04446_),
    .S(_04752_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09929_ (.I0(\dp.rf.rf[22][5] ),
    .I1(_04455_),
    .S(_04752_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09930_ (.A1(\dp.rf.rf[22][6] ),
    .A2(_04755_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09931_ (.A1(_04466_),
    .A2(_04755_),
    .B(_04765_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09932_ (.I0(\dp.rf.rf[22][7] ),
    .I1(_04473_),
    .S(_04752_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09933_ (.A1(\dp.rf.rf[22][8] ),
    .A2(_04755_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09934_ (.A1(_04485_),
    .A2(_04755_),
    .B(_04766_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09935_ (.I0(\dp.rf.rf[22][9] ),
    .I1(_04497_),
    .S(_04752_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09936_ (.A1(_04499_),
    .A2(_04713_),
    .Z(_04767_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output105 (.I(net105),
    .Z(pc[14]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output104 (.I(net104),
    .Z(pc[13]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09939_ (.I0(\dp.rf.rf[23][0] ),
    .I1(net478),
    .S(_04767_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09940_ (.I0(\dp.rf.rf[23][10] ),
    .I1(_04069_),
    .S(_04767_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09941_ (.I0(\dp.rf.rf[23][11] ),
    .I1(_04092_),
    .S(_04767_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09942_ (.I0(\dp.rf.rf[23][12] ),
    .I1(_04106_),
    .S(_04767_),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09943_ (.I0(\dp.rf.rf[23][13] ),
    .I1(_04119_),
    .S(_04767_),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09944_ (.I0(\dp.rf.rf[23][14] ),
    .I1(_04136_),
    .S(_04767_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09945_ (.I0(\dp.rf.rf[23][15] ),
    .I1(_04152_),
    .S(_04767_),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09946_ (.A1(_04499_),
    .A2(_04713_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output103 (.I(net103),
    .Z(pc[12]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09948_ (.A1(\dp.rf.rf[23][16] ),
    .A2(_04770_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09949_ (.A1(_04178_),
    .A2(_04770_),
    .B(_04772_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09950_ (.I0(\dp.rf.rf[23][17] ),
    .I1(net483),
    .S(_04767_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09951_ (.I0(\dp.rf.rf[23][18] ),
    .I1(net482),
    .S(_04767_),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09952_ (.I0(\dp.rf.rf[23][19] ),
    .I1(_04222_),
    .S(_04767_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output102 (.I(net102),
    .Z(pc[11]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09954_ (.I0(\dp.rf.rf[23][1] ),
    .I1(_04228_),
    .S(_04767_),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09955_ (.A1(\dp.rf.rf[23][20] ),
    .A2(_04770_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09956_ (.A1(_04250_),
    .A2(_04770_),
    .B(_04774_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09957_ (.I0(\dp.rf.rf[23][21] ),
    .I1(_04267_),
    .S(_04767_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09958_ (.I0(\dp.rf.rf[23][22] ),
    .I1(net481),
    .S(_04767_),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09959_ (.A1(_04301_),
    .A2(_04767_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09960_ (.A1(_01808_),
    .A2(_04770_),
    .B1(_04775_),
    .B2(net485),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09961_ (.I0(\dp.rf.rf[23][24] ),
    .I1(_04314_),
    .S(_04767_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09962_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04767_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09963_ (.A1(_01667_),
    .A2(_04770_),
    .B1(_04776_),
    .B2(_04325_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09964_ (.I0(\dp.rf.rf[23][26] ),
    .I1(_04343_),
    .S(_04767_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09965_ (.I0(\dp.rf.rf[23][27] ),
    .I1(_04355_),
    .S(_04767_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09966_ (.I0(\dp.rf.rf[23][28] ),
    .I1(_04370_),
    .S(_04767_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09967_ (.I(\dp.rf.rf[23][29] ),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _09968_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04767_),
    .Z(_04778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09969_ (.A1(_04777_),
    .A2(_04770_),
    .B1(_04778_),
    .B2(net480),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09970_ (.I0(\dp.rf.rf[23][2] ),
    .I1(_04396_),
    .S(_04767_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09971_ (.I0(\dp.rf.rf[23][30] ),
    .I1(net477),
    .S(_04767_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _09972_ (.A1(_04429_),
    .A2(_04767_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _09973_ (.A1(_01263_),
    .A2(_04770_),
    .B1(_04779_),
    .B2(net479),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09974_ (.I0(\dp.rf.rf[23][3] ),
    .I1(_04436_),
    .S(_04767_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09975_ (.I0(\dp.rf.rf[23][4] ),
    .I1(_04446_),
    .S(_04767_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09976_ (.I0(\dp.rf.rf[23][5] ),
    .I1(_04455_),
    .S(_04767_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09977_ (.A1(\dp.rf.rf[23][6] ),
    .A2(_04770_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09978_ (.A1(_04466_),
    .A2(_04770_),
    .B(_04780_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09979_ (.I0(\dp.rf.rf[23][7] ),
    .I1(_04473_),
    .S(_04767_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09980_ (.A1(\dp.rf.rf[23][8] ),
    .A2(_04770_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09981_ (.A1(_04485_),
    .A2(_04770_),
    .B(_04781_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09982_ (.I0(\dp.rf.rf[23][9] ),
    .I1(_04497_),
    .S(_04767_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _09983_ (.A1(net3),
    .A2(net2),
    .A3(_04027_),
    .Z(_04782_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _09984_ (.A1(_04533_),
    .A2(_04782_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output101 (.I(net101),
    .Z(pc[10]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output100 (.I(net100),
    .Z(pc[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09987_ (.I0(\dp.rf.rf[24][0] ),
    .I1(net478),
    .S(_04783_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09988_ (.I0(\dp.rf.rf[24][10] ),
    .I1(_04069_),
    .S(_04783_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09989_ (.I0(\dp.rf.rf[24][11] ),
    .I1(_04092_),
    .S(_04783_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09990_ (.I0(\dp.rf.rf[24][12] ),
    .I1(_04106_),
    .S(_04783_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09991_ (.I0(\dp.rf.rf[24][13] ),
    .I1(_04119_),
    .S(_04783_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09992_ (.I0(\dp.rf.rf[24][14] ),
    .I1(_04136_),
    .S(_04783_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09993_ (.I0(\dp.rf.rf[24][15] ),
    .I1(_04152_),
    .S(_04783_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _09994_ (.A1(_04533_),
    .A2(_04782_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output99 (.I(net99),
    .Z(memwrite));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _09996_ (.A1(\dp.rf.rf[24][16] ),
    .A2(_04786_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _09997_ (.A1(_04178_),
    .A2(_04786_),
    .B(_04788_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09998_ (.I0(\dp.rf.rf[24][17] ),
    .I1(net483),
    .S(_04783_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _09999_ (.I0(\dp.rf.rf[24][18] ),
    .I1(net482),
    .S(_04783_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10000_ (.I0(\dp.rf.rf[24][19] ),
    .I1(_04222_),
    .S(_04783_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output98 (.I(net98),
    .Z(memread));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10002_ (.I0(\dp.rf.rf[24][1] ),
    .I1(_04228_),
    .S(_04783_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10003_ (.A1(\dp.rf.rf[24][20] ),
    .A2(_04786_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10004_ (.A1(_04250_),
    .A2(_04786_),
    .B(_04790_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10005_ (.I0(\dp.rf.rf[24][21] ),
    .I1(_04267_),
    .S(_04783_),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10006_ (.I0(\dp.rf.rf[24][22] ),
    .I1(net481),
    .S(_04783_),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10007_ (.A1(_04301_),
    .A2(_04783_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10008_ (.A1(_01788_),
    .A2(_04786_),
    .B1(_04791_),
    .B2(net485),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10009_ (.I0(\dp.rf.rf[24][24] ),
    .I1(_04314_),
    .S(_04783_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10010_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04783_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10011_ (.A1(_01669_),
    .A2(_04786_),
    .B1(_04792_),
    .B2(net484),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10012_ (.I0(\dp.rf.rf[24][26] ),
    .I1(_04343_),
    .S(_04783_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10013_ (.I0(\dp.rf.rf[24][27] ),
    .I1(_04355_),
    .S(_04783_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10014_ (.I0(\dp.rf.rf[24][28] ),
    .I1(_04370_),
    .S(_04783_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10015_ (.I(\dp.rf.rf[24][29] ),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10016_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04783_),
    .Z(_04794_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10017_ (.A1(_04793_),
    .A2(_04786_),
    .B1(_04794_),
    .B2(net480),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10018_ (.I0(\dp.rf.rf[24][2] ),
    .I1(_04396_),
    .S(_04783_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10019_ (.I0(\dp.rf.rf[24][30] ),
    .I1(net477),
    .S(_04783_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10020_ (.I(\dp.rf.rf[24][31] ),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10021_ (.A1(_04429_),
    .A2(_04783_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10022_ (.A1(_04795_),
    .A2(_04786_),
    .B1(_04796_),
    .B2(net479),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10023_ (.I0(\dp.rf.rf[24][3] ),
    .I1(_04436_),
    .S(_04783_),
    .Z(_00540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10024_ (.I0(\dp.rf.rf[24][4] ),
    .I1(_04446_),
    .S(_04783_),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10025_ (.I0(\dp.rf.rf[24][5] ),
    .I1(_04455_),
    .S(_04783_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10026_ (.A1(\dp.rf.rf[24][6] ),
    .A2(_04786_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10027_ (.A1(_04466_),
    .A2(_04786_),
    .B(_04797_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10028_ (.I0(\dp.rf.rf[24][7] ),
    .I1(_04473_),
    .S(_04783_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10029_ (.A1(\dp.rf.rf[24][8] ),
    .A2(_04786_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10030_ (.A1(_04485_),
    .A2(_04786_),
    .B(_04798_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10031_ (.I0(\dp.rf.rf[24][9] ),
    .I1(_04497_),
    .S(_04783_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10032_ (.A1(_04552_),
    .A2(_04782_),
    .Z(_04799_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output97 (.I(net97),
    .Z(aluout[9]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output96 (.I(net96),
    .Z(aluout[8]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10035_ (.I0(\dp.rf.rf[25][0] ),
    .I1(net478),
    .S(_04799_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10036_ (.I0(\dp.rf.rf[25][10] ),
    .I1(_04069_),
    .S(_04799_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10037_ (.I0(\dp.rf.rf[25][11] ),
    .I1(_04092_),
    .S(_04799_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10038_ (.I0(\dp.rf.rf[25][12] ),
    .I1(_04106_),
    .S(_04799_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10039_ (.I0(\dp.rf.rf[25][13] ),
    .I1(_04119_),
    .S(_04799_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10040_ (.I0(\dp.rf.rf[25][14] ),
    .I1(_04136_),
    .S(_04799_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10041_ (.I0(\dp.rf.rf[25][15] ),
    .I1(_04152_),
    .S(_04799_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10042_ (.A1(_04552_),
    .A2(_04782_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output95 (.I(net95),
    .Z(aluout[7]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10044_ (.A1(\dp.rf.rf[25][16] ),
    .A2(_04802_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10045_ (.A1(_04178_),
    .A2(_04802_),
    .B(_04804_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10046_ (.I0(\dp.rf.rf[25][17] ),
    .I1(net483),
    .S(_04799_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10047_ (.I0(\dp.rf.rf[25][18] ),
    .I1(net482),
    .S(_04799_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10048_ (.I0(\dp.rf.rf[25][19] ),
    .I1(_04222_),
    .S(_04799_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output94 (.I(net94),
    .Z(aluout[6]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10050_ (.I0(\dp.rf.rf[25][1] ),
    .I1(_04228_),
    .S(_04799_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10051_ (.A1(\dp.rf.rf[25][20] ),
    .A2(_04802_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10052_ (.A1(_04250_),
    .A2(_04802_),
    .B(_04806_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10053_ (.I0(\dp.rf.rf[25][21] ),
    .I1(_04267_),
    .S(_04799_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10054_ (.I0(\dp.rf.rf[25][22] ),
    .I1(net481),
    .S(_04799_),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10055_ (.A1(_04301_),
    .A2(_04799_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10056_ (.A1(_01789_),
    .A2(_04802_),
    .B1(_04807_),
    .B2(net485),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10057_ (.I0(\dp.rf.rf[25][24] ),
    .I1(_04314_),
    .S(_04799_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10058_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04799_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10059_ (.A1(_01670_),
    .A2(_04802_),
    .B1(_04808_),
    .B2(net484),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10060_ (.I0(\dp.rf.rf[25][26] ),
    .I1(_04343_),
    .S(_04799_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10061_ (.I0(\dp.rf.rf[25][27] ),
    .I1(_04355_),
    .S(_04799_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10062_ (.I0(\dp.rf.rf[25][28] ),
    .I1(_04370_),
    .S(_04799_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10063_ (.I(\dp.rf.rf[25][29] ),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10064_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04799_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10065_ (.A1(_04809_),
    .A2(_04802_),
    .B1(_04810_),
    .B2(net480),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10066_ (.I0(\dp.rf.rf[25][2] ),
    .I1(_04396_),
    .S(_04799_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10067_ (.I0(\dp.rf.rf[25][30] ),
    .I1(net477),
    .S(_04799_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10068_ (.A1(_04429_),
    .A2(_04799_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10069_ (.A1(_01267_),
    .A2(_04802_),
    .B1(_04811_),
    .B2(net479),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10070_ (.I0(\dp.rf.rf[25][3] ),
    .I1(_04436_),
    .S(_04799_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10071_ (.I0(\dp.rf.rf[25][4] ),
    .I1(_04446_),
    .S(_04799_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10072_ (.I0(\dp.rf.rf[25][5] ),
    .I1(_04455_),
    .S(_04799_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10073_ (.A1(\dp.rf.rf[25][6] ),
    .A2(_04802_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10074_ (.A1(_04466_),
    .A2(_04802_),
    .B(_04812_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10075_ (.I0(\dp.rf.rf[25][7] ),
    .I1(_04473_),
    .S(_04799_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10076_ (.A1(\dp.rf.rf[25][8] ),
    .A2(_04802_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10077_ (.A1(_04485_),
    .A2(_04802_),
    .B(_04813_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10078_ (.I0(\dp.rf.rf[25][9] ),
    .I1(_04497_),
    .S(_04799_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10079_ (.A1(_04034_),
    .A2(_04782_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output93 (.I(net93),
    .Z(aluout[5]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output92 (.I(net92),
    .Z(aluout[4]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10082_ (.I0(\dp.rf.rf[26][0] ),
    .I1(net478),
    .S(_04814_),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10083_ (.I0(\dp.rf.rf[26][10] ),
    .I1(_04069_),
    .S(_04814_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10084_ (.I0(\dp.rf.rf[26][11] ),
    .I1(_04092_),
    .S(_04814_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10085_ (.I0(\dp.rf.rf[26][12] ),
    .I1(_04106_),
    .S(_04814_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10086_ (.I0(\dp.rf.rf[26][13] ),
    .I1(_04119_),
    .S(_04814_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10087_ (.I0(\dp.rf.rf[26][14] ),
    .I1(_04136_),
    .S(_04814_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10088_ (.I0(\dp.rf.rf[26][15] ),
    .I1(_04152_),
    .S(_04814_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10089_ (.A1(_04034_),
    .A2(_04782_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output91 (.I(net91),
    .Z(aluout[3]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10091_ (.A1(\dp.rf.rf[26][16] ),
    .A2(_04817_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10092_ (.A1(_04178_),
    .A2(_04817_),
    .B(_04819_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10093_ (.I0(\dp.rf.rf[26][17] ),
    .I1(net483),
    .S(_04814_),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10094_ (.I0(\dp.rf.rf[26][18] ),
    .I1(net482),
    .S(_04814_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10095_ (.I0(\dp.rf.rf[26][19] ),
    .I1(_04222_),
    .S(_04814_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output90 (.I(net90),
    .Z(aluout[31]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10097_ (.I0(\dp.rf.rf[26][1] ),
    .I1(_04228_),
    .S(_04814_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10098_ (.A1(\dp.rf.rf[26][20] ),
    .A2(_04817_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10099_ (.A1(_04250_),
    .A2(_04817_),
    .B(_04821_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10100_ (.I0(\dp.rf.rf[26][21] ),
    .I1(_04267_),
    .S(_04814_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10101_ (.I0(\dp.rf.rf[26][22] ),
    .I1(net481),
    .S(_04814_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10102_ (.A1(_04301_),
    .A2(_04814_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10103_ (.A1(_01790_),
    .A2(_04817_),
    .B1(_04822_),
    .B2(net485),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10104_ (.I0(\dp.rf.rf[26][24] ),
    .I1(_04314_),
    .S(_04814_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10105_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04814_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10106_ (.A1(_01671_),
    .A2(_04817_),
    .B1(_04823_),
    .B2(net484),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10107_ (.I0(\dp.rf.rf[26][26] ),
    .I1(_04343_),
    .S(_04814_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10108_ (.I0(\dp.rf.rf[26][27] ),
    .I1(_04355_),
    .S(_04814_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10109_ (.I0(\dp.rf.rf[26][28] ),
    .I1(_04370_),
    .S(_04814_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10110_ (.I(\dp.rf.rf[26][29] ),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10111_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04814_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10112_ (.A1(_04824_),
    .A2(_04817_),
    .B1(_04825_),
    .B2(net480),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10113_ (.I0(\dp.rf.rf[26][2] ),
    .I1(_04396_),
    .S(_04814_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10114_ (.I0(\dp.rf.rf[26][30] ),
    .I1(net477),
    .S(_04814_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10115_ (.I(\dp.rf.rf[26][31] ),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10116_ (.A1(_04429_),
    .A2(_04814_),
    .Z(_04827_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10117_ (.A1(_04826_),
    .A2(_04817_),
    .B1(_04827_),
    .B2(net479),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10118_ (.I0(\dp.rf.rf[26][3] ),
    .I1(_04436_),
    .S(_04814_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10119_ (.I0(\dp.rf.rf[26][4] ),
    .I1(_04446_),
    .S(_04814_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10120_ (.I0(\dp.rf.rf[26][5] ),
    .I1(_04455_),
    .S(_04814_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10121_ (.A1(\dp.rf.rf[26][6] ),
    .A2(_04817_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10122_ (.A1(_04466_),
    .A2(_04817_),
    .B(_04828_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10123_ (.I0(\dp.rf.rf[26][7] ),
    .I1(_04473_),
    .S(_04814_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10124_ (.A1(\dp.rf.rf[26][8] ),
    .A2(_04817_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10125_ (.A1(_04485_),
    .A2(_04817_),
    .B(_04829_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10126_ (.I0(\dp.rf.rf[26][9] ),
    .I1(_04497_),
    .S(_04814_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10127_ (.A1(_04499_),
    .A2(_04782_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output89 (.I(net89),
    .Z(aluout[30]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output88 (.I(net88),
    .Z(aluout[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10130_ (.I0(\dp.rf.rf[27][0] ),
    .I1(net478),
    .S(_04830_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10131_ (.I0(\dp.rf.rf[27][10] ),
    .I1(_04069_),
    .S(_04830_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10132_ (.I0(\dp.rf.rf[27][11] ),
    .I1(_04092_),
    .S(_04830_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10133_ (.I0(\dp.rf.rf[27][12] ),
    .I1(_04106_),
    .S(_04830_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10134_ (.I0(\dp.rf.rf[27][13] ),
    .I1(_04119_),
    .S(_04830_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10135_ (.I0(\dp.rf.rf[27][14] ),
    .I1(_04136_),
    .S(_04830_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10136_ (.I0(\dp.rf.rf[27][15] ),
    .I1(_04152_),
    .S(_04830_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10137_ (.A1(_04499_),
    .A2(_04782_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output87 (.I(net87),
    .Z(aluout[29]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10139_ (.A1(\dp.rf.rf[27][16] ),
    .A2(_04833_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10140_ (.A1(_04178_),
    .A2(_04833_),
    .B(_04835_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10141_ (.I0(\dp.rf.rf[27][17] ),
    .I1(net483),
    .S(_04830_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10142_ (.I0(\dp.rf.rf[27][18] ),
    .I1(net482),
    .S(_04830_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10143_ (.I0(\dp.rf.rf[27][19] ),
    .I1(_04222_),
    .S(_04830_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output86 (.I(net86),
    .Z(aluout[28]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10145_ (.I0(\dp.rf.rf[27][1] ),
    .I1(_04228_),
    .S(_04830_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10146_ (.A1(\dp.rf.rf[27][20] ),
    .A2(_04833_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10147_ (.A1(_04250_),
    .A2(_04833_),
    .B(_04837_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10148_ (.I0(\dp.rf.rf[27][21] ),
    .I1(_04267_),
    .S(_04830_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10149_ (.I0(\dp.rf.rf[27][22] ),
    .I1(net481),
    .S(_04830_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10150_ (.A1(_04301_),
    .A2(_04830_),
    .Z(_04838_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10151_ (.A1(_01791_),
    .A2(_04833_),
    .B1(_04838_),
    .B2(net485),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10152_ (.I0(\dp.rf.rf[27][24] ),
    .I1(_04314_),
    .S(_04830_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10153_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04830_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10154_ (.A1(_01672_),
    .A2(_04833_),
    .B1(_04839_),
    .B2(net484),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10155_ (.I0(\dp.rf.rf[27][26] ),
    .I1(_04343_),
    .S(_04830_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10156_ (.I0(\dp.rf.rf[27][27] ),
    .I1(_04355_),
    .S(_04830_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10157_ (.I0(\dp.rf.rf[27][28] ),
    .I1(_04370_),
    .S(_04830_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10158_ (.I(\dp.rf.rf[27][29] ),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10159_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04830_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10160_ (.A1(_04840_),
    .A2(_04833_),
    .B1(_04841_),
    .B2(net480),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10161_ (.I0(\dp.rf.rf[27][2] ),
    .I1(_04396_),
    .S(_04830_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10162_ (.I0(\dp.rf.rf[27][30] ),
    .I1(net477),
    .S(_04830_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10163_ (.I(\dp.rf.rf[27][31] ),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10164_ (.A1(_04429_),
    .A2(_04830_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10165_ (.A1(_04842_),
    .A2(_04833_),
    .B1(_04843_),
    .B2(net479),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10166_ (.I0(\dp.rf.rf[27][3] ),
    .I1(_04436_),
    .S(_04830_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10167_ (.I0(\dp.rf.rf[27][4] ),
    .I1(_04446_),
    .S(_04830_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10168_ (.I0(\dp.rf.rf[27][5] ),
    .I1(_04455_),
    .S(_04830_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10169_ (.A1(\dp.rf.rf[27][6] ),
    .A2(_04833_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10170_ (.A1(_04466_),
    .A2(_04833_),
    .B(_04844_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10171_ (.I0(\dp.rf.rf[27][7] ),
    .I1(_04473_),
    .S(_04830_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10172_ (.A1(\dp.rf.rf[27][8] ),
    .A2(_04833_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10173_ (.A1(_04485_),
    .A2(_04833_),
    .B(_04845_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10174_ (.I0(\dp.rf.rf[27][9] ),
    .I1(_04497_),
    .S(_04830_),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _10175_ (.A1(net3),
    .A2(net2),
    .A3(net32),
    .Z(_04846_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10176_ (.A1(_04533_),
    .A2(_04846_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output85 (.I(net85),
    .Z(aluout[27]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output84 (.I(net84),
    .Z(aluout[26]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10179_ (.I0(\dp.rf.rf[28][0] ),
    .I1(net478),
    .S(_04847_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10180_ (.I0(\dp.rf.rf[28][10] ),
    .I1(_04069_),
    .S(_04847_),
    .Z(_00644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10181_ (.I0(\dp.rf.rf[28][11] ),
    .I1(_04092_),
    .S(_04847_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10182_ (.I0(\dp.rf.rf[28][12] ),
    .I1(_04106_),
    .S(_04847_),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10183_ (.I0(\dp.rf.rf[28][13] ),
    .I1(_04119_),
    .S(_04847_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10184_ (.I0(\dp.rf.rf[28][14] ),
    .I1(_04136_),
    .S(_04847_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10185_ (.I0(\dp.rf.rf[28][15] ),
    .I1(_04152_),
    .S(_04847_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10186_ (.A1(_04533_),
    .A2(_04846_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output83 (.I(net83),
    .Z(aluout[25]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10188_ (.A1(\dp.rf.rf[28][16] ),
    .A2(_04850_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10189_ (.A1(_04178_),
    .A2(_04850_),
    .B(_04852_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10190_ (.I0(\dp.rf.rf[28][17] ),
    .I1(net483),
    .S(_04847_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10191_ (.I0(\dp.rf.rf[28][18] ),
    .I1(net482),
    .S(_04847_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10192_ (.I0(\dp.rf.rf[28][19] ),
    .I1(_04222_),
    .S(_04847_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output82 (.I(net82),
    .Z(aluout[24]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10194_ (.I0(\dp.rf.rf[28][1] ),
    .I1(_04228_),
    .S(_04847_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10195_ (.A1(\dp.rf.rf[28][20] ),
    .A2(_04850_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10196_ (.A1(_04250_),
    .A2(_04850_),
    .B(_04854_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10197_ (.I0(\dp.rf.rf[28][21] ),
    .I1(_04267_),
    .S(_04847_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10198_ (.I0(\dp.rf.rf[28][22] ),
    .I1(net481),
    .S(_04847_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10199_ (.A1(_04301_),
    .A2(_04847_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10200_ (.A1(_01800_),
    .A2(_04850_),
    .B1(_04855_),
    .B2(net485),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10201_ (.I0(\dp.rf.rf[28][24] ),
    .I1(_04314_),
    .S(_04847_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10202_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04847_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10203_ (.A1(_01659_),
    .A2(_04850_),
    .B1(_04856_),
    .B2(net484),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10204_ (.I0(\dp.rf.rf[28][26] ),
    .I1(_04343_),
    .S(_04847_),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10205_ (.I0(\dp.rf.rf[28][27] ),
    .I1(_04355_),
    .S(_04847_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10206_ (.I0(\dp.rf.rf[28][28] ),
    .I1(_04370_),
    .S(_04847_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10207_ (.I(\dp.rf.rf[28][29] ),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10208_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04847_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10209_ (.A1(_04857_),
    .A2(_04850_),
    .B1(_04858_),
    .B2(net480),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10210_ (.I0(\dp.rf.rf[28][2] ),
    .I1(_04396_),
    .S(_04847_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10211_ (.I0(\dp.rf.rf[28][30] ),
    .I1(net477),
    .S(_04847_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10212_ (.I(\dp.rf.rf[28][31] ),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10213_ (.A1(_04429_),
    .A2(_04847_),
    .Z(_04860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10214_ (.A1(_04859_),
    .A2(_04850_),
    .B1(_04860_),
    .B2(net479),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10215_ (.I0(\dp.rf.rf[28][3] ),
    .I1(_04436_),
    .S(_04847_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10216_ (.I0(\dp.rf.rf[28][4] ),
    .I1(_04446_),
    .S(_04847_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10217_ (.I0(\dp.rf.rf[28][5] ),
    .I1(_04455_),
    .S(_04847_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10218_ (.A1(\dp.rf.rf[28][6] ),
    .A2(_04850_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10219_ (.A1(_04466_),
    .A2(_04850_),
    .B(_04861_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10220_ (.I0(\dp.rf.rf[28][7] ),
    .I1(_04473_),
    .S(_04847_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10221_ (.A1(\dp.rf.rf[28][8] ),
    .A2(_04850_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10222_ (.A1(_04485_),
    .A2(_04850_),
    .B(_04862_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10223_ (.I0(\dp.rf.rf[28][9] ),
    .I1(_04497_),
    .S(_04847_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output81 (.I(net81),
    .Z(aluout[23]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10225_ (.A1(_04552_),
    .A2(_04846_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output80 (.I(net80),
    .Z(aluout[22]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output79 (.I(net79),
    .Z(aluout[21]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10228_ (.I0(\dp.rf.rf[29][0] ),
    .I1(net478),
    .S(_04864_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output78 (.I(net78),
    .Z(aluout[20]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10230_ (.I0(\dp.rf.rf[29][10] ),
    .I1(_04069_),
    .S(_04864_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output77 (.I(net77),
    .Z(aluout[1]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10232_ (.I0(\dp.rf.rf[29][11] ),
    .I1(_04092_),
    .S(_04864_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output76 (.I(net76),
    .Z(aluout[19]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10234_ (.I0(\dp.rf.rf[29][12] ),
    .I1(_04106_),
    .S(_04864_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output75 (.I(net75),
    .Z(aluout[18]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10236_ (.I0(\dp.rf.rf[29][13] ),
    .I1(_04119_),
    .S(_04864_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output74 (.I(net74),
    .Z(aluout[17]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10238_ (.I0(\dp.rf.rf[29][14] ),
    .I1(_04136_),
    .S(_04864_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output73 (.I(net73),
    .Z(aluout[16]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10240_ (.I0(\dp.rf.rf[29][15] ),
    .I1(_04152_),
    .S(_04864_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10241_ (.A1(_04552_),
    .A2(_04846_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output72 (.I(net72),
    .Z(aluout[15]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10243_ (.A1(\dp.rf.rf[29][16] ),
    .A2(_04873_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10244_ (.A1(_04178_),
    .A2(_04873_),
    .B(_04875_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output71 (.I(net71),
    .Z(aluout[14]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10246_ (.I0(\dp.rf.rf[29][17] ),
    .I1(net483),
    .S(_04864_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output70 (.I(net70),
    .Z(aluout[13]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10248_ (.I0(\dp.rf.rf[29][18] ),
    .I1(net482),
    .S(_04864_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output69 (.I(net69),
    .Z(aluout[12]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10250_ (.I0(\dp.rf.rf[29][19] ),
    .I1(_04222_),
    .S(_04864_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output68 (.I(net68),
    .Z(aluout[11]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output67 (.I(net67),
    .Z(aluout[10]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10253_ (.I0(\dp.rf.rf[29][1] ),
    .I1(_04228_),
    .S(_04864_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10254_ (.A1(\dp.rf.rf[29][20] ),
    .A2(_04873_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10255_ (.A1(_04250_),
    .A2(_04873_),
    .B(_04881_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output66 (.I(net66),
    .Z(aluout[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10257_ (.I0(\dp.rf.rf[29][21] ),
    .I1(_04267_),
    .S(_04864_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input65 (.I(reset),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10259_ (.I0(\dp.rf.rf[29][22] ),
    .I1(net481),
    .S(_04864_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10260_ (.A1(_04301_),
    .A2(_04864_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input64 (.I(readdata[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10262_ (.A1(_01801_),
    .A2(_04873_),
    .B1(_04884_),
    .B2(net485),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input63 (.I(readdata[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10264_ (.I0(\dp.rf.rf[29][24] ),
    .I1(_04314_),
    .S(_04864_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10265_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04864_),
    .Z(_04887_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input62 (.I(readdata[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10267_ (.A1(_01660_),
    .A2(_04873_),
    .B1(_04887_),
    .B2(net484),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input61 (.I(readdata[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10269_ (.I0(\dp.rf.rf[29][26] ),
    .I1(_04343_),
    .S(_04864_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input60 (.I(readdata[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10271_ (.I0(\dp.rf.rf[29][27] ),
    .I1(_04355_),
    .S(_04864_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input59 (.I(readdata[4]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10273_ (.I0(\dp.rf.rf[29][28] ),
    .I1(_04370_),
    .S(_04864_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10274_ (.I(\dp.rf.rf[29][29] ),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10275_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04864_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input58 (.I(readdata[3]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10277_ (.A1(_04892_),
    .A2(_04873_),
    .B1(_04893_),
    .B2(net480),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input57 (.I(readdata[31]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10279_ (.I0(\dp.rf.rf[29][2] ),
    .I1(_04396_),
    .S(_04864_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input56 (.I(readdata[30]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10281_ (.I0(\dp.rf.rf[29][30] ),
    .I1(net477),
    .S(_04864_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10282_ (.I(\dp.rf.rf[29][31] ),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10283_ (.A1(_04429_),
    .A2(_04864_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input55 (.I(readdata[2]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10285_ (.A1(_04897_),
    .A2(_04873_),
    .B1(_04898_),
    .B2(net479),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input54 (.I(readdata[29]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10287_ (.I0(\dp.rf.rf[29][3] ),
    .I1(_04436_),
    .S(_04864_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input53 (.I(readdata[28]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10289_ (.I0(\dp.rf.rf[29][4] ),
    .I1(_04446_),
    .S(_04864_),
    .Z(_00701_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input52 (.I(readdata[27]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10291_ (.I0(\dp.rf.rf[29][5] ),
    .I1(_04455_),
    .S(_04864_),
    .Z(_00702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10292_ (.A1(\dp.rf.rf[29][6] ),
    .A2(_04873_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10293_ (.A1(_04466_),
    .A2(_04873_),
    .B(_04903_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input51 (.I(readdata[26]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10295_ (.I0(\dp.rf.rf[29][7] ),
    .I1(_04473_),
    .S(_04864_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10296_ (.A1(\dp.rf.rf[29][8] ),
    .A2(_04873_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10297_ (.A1(_04485_),
    .A2(_04873_),
    .B(_04905_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input50 (.I(readdata[25]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10299_ (.I0(\dp.rf.rf[29][9] ),
    .I1(_04497_),
    .S(_04864_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10300_ (.A1(_04034_),
    .A2(_04532_),
    .Z(_04907_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input49 (.I(readdata[24]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input48 (.I(readdata[23]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10303_ (.I0(\dp.rf.rf[2][0] ),
    .I1(net478),
    .S(_04907_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10304_ (.I0(\dp.rf.rf[2][10] ),
    .I1(_04069_),
    .S(_04907_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10305_ (.I0(\dp.rf.rf[2][11] ),
    .I1(_04092_),
    .S(_04907_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10306_ (.I0(\dp.rf.rf[2][12] ),
    .I1(_04106_),
    .S(_04907_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10307_ (.I0(\dp.rf.rf[2][13] ),
    .I1(_04119_),
    .S(_04907_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10308_ (.I0(\dp.rf.rf[2][14] ),
    .I1(_04136_),
    .S(_04907_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10309_ (.I0(\dp.rf.rf[2][15] ),
    .I1(_04152_),
    .S(_04907_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input47 (.I(readdata[22]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10311_ (.A1(_04034_),
    .A2(_04532_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input46 (.I(readdata[21]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10313_ (.A1(\dp.rf.rf[2][16] ),
    .A2(_04911_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10314_ (.A1(_04178_),
    .A2(_04911_),
    .B(_04913_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10315_ (.I0(\dp.rf.rf[2][17] ),
    .I1(net483),
    .S(_04907_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10316_ (.I0(\dp.rf.rf[2][18] ),
    .I1(net482),
    .S(_04907_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10317_ (.I0(\dp.rf.rf[2][19] ),
    .I1(_04222_),
    .S(_04907_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input45 (.I(readdata[20]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10319_ (.I0(\dp.rf.rf[2][1] ),
    .I1(_04228_),
    .S(_04907_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input44 (.I(readdata[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10321_ (.A1(\dp.rf.rf[2][20] ),
    .A2(_04911_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10322_ (.A1(_04250_),
    .A2(_04911_),
    .B(_04916_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10323_ (.I0(\dp.rf.rf[2][21] ),
    .I1(_04267_),
    .S(_04907_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10324_ (.I0(\dp.rf.rf[2][22] ),
    .I1(net481),
    .S(_04907_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input43 (.I(readdata[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10326_ (.A1(_04301_),
    .A2(_04907_),
    .Z(_04918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10327_ (.A1(_01834_),
    .A2(_04911_),
    .B1(_04918_),
    .B2(net485),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10328_ (.I0(\dp.rf.rf[2][24] ),
    .I1(_04314_),
    .S(_04907_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10329_ (.I(\dp.rf.rf[2][25] ),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input42 (.I(readdata[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input41 (.I(readdata[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10332_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04907_),
    .Z(_04922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10333_ (.A1(_04919_),
    .A2(_04911_),
    .B1(_04922_),
    .B2(_04325_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10334_ (.I0(\dp.rf.rf[2][26] ),
    .I1(_04343_),
    .S(_04907_),
    .Z(_00725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10335_ (.I0(\dp.rf.rf[2][27] ),
    .I1(_04355_),
    .S(_04907_),
    .Z(_00726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10336_ (.I0(\dp.rf.rf[2][28] ),
    .I1(_04370_),
    .S(_04907_),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10337_ (.I(\dp.rf.rf[2][29] ),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input40 (.I(readdata[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input39 (.I(readdata[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10340_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04907_),
    .Z(_04926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10341_ (.A1(_04923_),
    .A2(_04911_),
    .B1(_04926_),
    .B2(net480),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10342_ (.I0(\dp.rf.rf[2][2] ),
    .I1(_04396_),
    .S(_04907_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10343_ (.I0(\dp.rf.rf[2][30] ),
    .I1(net477),
    .S(_04907_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10344_ (.I(\dp.rf.rf[2][31] ),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input38 (.I(readdata[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10346_ (.A1(_04429_),
    .A2(_04907_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10347_ (.A1(_04927_),
    .A2(_04911_),
    .B1(_04929_),
    .B2(net479),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10348_ (.I0(\dp.rf.rf[2][3] ),
    .I1(_04436_),
    .S(_04907_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10349_ (.I0(\dp.rf.rf[2][4] ),
    .I1(_04446_),
    .S(_04907_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10350_ (.I0(\dp.rf.rf[2][5] ),
    .I1(_04455_),
    .S(_04907_),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input37 (.I(readdata[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10352_ (.A1(\dp.rf.rf[2][6] ),
    .A2(_04911_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10353_ (.A1(_04466_),
    .A2(_04911_),
    .B(_04931_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10354_ (.I0(\dp.rf.rf[2][7] ),
    .I1(_04473_),
    .S(_04907_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input36 (.I(readdata[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10356_ (.A1(\dp.rf.rf[2][8] ),
    .A2(_04911_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10357_ (.A1(_04485_),
    .A2(_04911_),
    .B(_04933_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10358_ (.I0(\dp.rf.rf[2][9] ),
    .I1(_04497_),
    .S(_04907_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10359_ (.A1(_04034_),
    .A2(_04846_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input35 (.I(readdata[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input34 (.I(readdata[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10362_ (.I0(\dp.rf.rf[30][0] ),
    .I1(net478),
    .S(_04934_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10363_ (.I0(\dp.rf.rf[30][10] ),
    .I1(_04069_),
    .S(_04934_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10364_ (.I0(\dp.rf.rf[30][11] ),
    .I1(_04092_),
    .S(_04934_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10365_ (.I0(\dp.rf.rf[30][12] ),
    .I1(_04106_),
    .S(_04934_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10366_ (.I0(\dp.rf.rf[30][13] ),
    .I1(_04119_),
    .S(_04934_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10367_ (.I0(\dp.rf.rf[30][14] ),
    .I1(_04136_),
    .S(_04934_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10368_ (.I0(\dp.rf.rf[30][15] ),
    .I1(_04152_),
    .S(_04934_),
    .Z(_00745_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10369_ (.A1(_04034_),
    .A2(_04846_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input33 (.I(readdata[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10371_ (.A1(\dp.rf.rf[30][16] ),
    .A2(_04937_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10372_ (.A1(_04178_),
    .A2(_04937_),
    .B(_04939_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10373_ (.I0(\dp.rf.rf[30][17] ),
    .I1(net483),
    .S(_04934_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10374_ (.I0(\dp.rf.rf[30][18] ),
    .I1(net482),
    .S(_04934_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10375_ (.I0(\dp.rf.rf[30][19] ),
    .I1(_04222_),
    .S(_04934_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input32 (.I(instr[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10377_ (.I0(\dp.rf.rf[30][1] ),
    .I1(_04228_),
    .S(_04934_),
    .Z(_00750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10378_ (.A1(\dp.rf.rf[30][20] ),
    .A2(_04937_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10379_ (.A1(_04250_),
    .A2(_04937_),
    .B(_04941_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10380_ (.I0(\dp.rf.rf[30][21] ),
    .I1(_04267_),
    .S(_04934_),
    .Z(_00752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10381_ (.I0(\dp.rf.rf[30][22] ),
    .I1(net481),
    .S(_04934_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10382_ (.A1(_04301_),
    .A2(_04934_),
    .Z(_04942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10383_ (.A1(_01802_),
    .A2(_04937_),
    .B1(_04942_),
    .B2(net485),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10384_ (.I0(\dp.rf.rf[30][24] ),
    .I1(_04314_),
    .S(_04934_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10385_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04934_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10386_ (.A1(_01661_),
    .A2(_04937_),
    .B1(_04943_),
    .B2(_04325_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10387_ (.I0(\dp.rf.rf[30][26] ),
    .I1(_04343_),
    .S(_04934_),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10388_ (.I0(\dp.rf.rf[30][27] ),
    .I1(_04355_),
    .S(_04934_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10389_ (.I0(\dp.rf.rf[30][28] ),
    .I1(_04370_),
    .S(_04934_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10390_ (.I(\dp.rf.rf[30][29] ),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10391_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04934_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10392_ (.A1(_04944_),
    .A2(_04937_),
    .B1(_04945_),
    .B2(net480),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10393_ (.I0(\dp.rf.rf[30][2] ),
    .I1(_04396_),
    .S(_04934_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10394_ (.I0(\dp.rf.rf[30][30] ),
    .I1(net477),
    .S(_04934_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10395_ (.I(\dp.rf.rf[30][31] ),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10396_ (.A1(_04429_),
    .A2(_04934_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10397_ (.A1(_04946_),
    .A2(_04937_),
    .B1(_04947_),
    .B2(net479),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10398_ (.I0(\dp.rf.rf[30][3] ),
    .I1(_04436_),
    .S(_04934_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10399_ (.I0(\dp.rf.rf[30][4] ),
    .I1(_04446_),
    .S(_04934_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10400_ (.I0(\dp.rf.rf[30][5] ),
    .I1(_04455_),
    .S(_04934_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10401_ (.A1(\dp.rf.rf[30][6] ),
    .A2(_04937_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10402_ (.A1(_04466_),
    .A2(_04937_),
    .B(_04948_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10403_ (.I0(\dp.rf.rf[30][7] ),
    .I1(_04473_),
    .S(_04934_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10404_ (.A1(\dp.rf.rf[30][8] ),
    .A2(_04937_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10405_ (.A1(_04485_),
    .A2(_04937_),
    .B(_04949_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10406_ (.I0(\dp.rf.rf[30][9] ),
    .I1(_04497_),
    .S(_04934_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10407_ (.A1(_04499_),
    .A2(_04846_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input31 (.I(instr[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input30 (.I(instr[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10410_ (.I0(\dp.rf.rf[31][0] ),
    .I1(net478),
    .S(_04950_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10411_ (.I0(\dp.rf.rf[31][10] ),
    .I1(_04069_),
    .S(_04950_),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10412_ (.I0(\dp.rf.rf[31][11] ),
    .I1(_04092_),
    .S(_04950_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10413_ (.I0(\dp.rf.rf[31][12] ),
    .I1(_04106_),
    .S(_04950_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10414_ (.I0(\dp.rf.rf[31][13] ),
    .I1(_04119_),
    .S(_04950_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10415_ (.I0(\dp.rf.rf[31][14] ),
    .I1(_04136_),
    .S(_04950_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10416_ (.I0(\dp.rf.rf[31][15] ),
    .I1(_04152_),
    .S(_04950_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10417_ (.A1(_04499_),
    .A2(_04846_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input29 (.I(instr[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10419_ (.A1(\dp.rf.rf[31][16] ),
    .A2(_04953_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10420_ (.A1(_04178_),
    .A2(_04953_),
    .B(_04955_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10421_ (.I0(\dp.rf.rf[31][17] ),
    .I1(net483),
    .S(_04950_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10422_ (.I0(\dp.rf.rf[31][18] ),
    .I1(net482),
    .S(_04950_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10423_ (.I0(\dp.rf.rf[31][19] ),
    .I1(_04222_),
    .S(_04950_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input28 (.I(instr[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10425_ (.I0(\dp.rf.rf[31][1] ),
    .I1(_04228_),
    .S(_04950_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10426_ (.A1(\dp.rf.rf[31][20] ),
    .A2(_04953_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10427_ (.A1(_04250_),
    .A2(_04953_),
    .B(_04957_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10428_ (.I0(\dp.rf.rf[31][21] ),
    .I1(_04267_),
    .S(_04950_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10429_ (.I0(\dp.rf.rf[31][22] ),
    .I1(net481),
    .S(_04950_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10430_ (.A1(_04301_),
    .A2(_04950_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10431_ (.A1(_01803_),
    .A2(_04953_),
    .B1(_04958_),
    .B2(net485),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10432_ (.I0(\dp.rf.rf[31][24] ),
    .I1(_04314_),
    .S(_04950_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10433_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04950_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10434_ (.A1(_01662_),
    .A2(_04953_),
    .B1(_04959_),
    .B2(net484),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10435_ (.I0(\dp.rf.rf[31][26] ),
    .I1(_04343_),
    .S(_04950_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10436_ (.I0(\dp.rf.rf[31][27] ),
    .I1(_04355_),
    .S(_04950_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10437_ (.I0(\dp.rf.rf[31][28] ),
    .I1(_04370_),
    .S(_04950_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10438_ (.I(\dp.rf.rf[31][29] ),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10439_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04950_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10440_ (.A1(_04960_),
    .A2(_04953_),
    .B1(_04961_),
    .B2(net480),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10441_ (.I0(\dp.rf.rf[31][2] ),
    .I1(_04396_),
    .S(_04950_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10442_ (.I0(\dp.rf.rf[31][30] ),
    .I1(net477),
    .S(_04950_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10443_ (.I(\dp.rf.rf[31][31] ),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10444_ (.A1(_04429_),
    .A2(_04950_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10445_ (.A1(_04962_),
    .A2(_04953_),
    .B1(_04963_),
    .B2(net479),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10446_ (.I0(\dp.rf.rf[31][3] ),
    .I1(_04436_),
    .S(_04950_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10447_ (.I0(\dp.rf.rf[31][4] ),
    .I1(_04446_),
    .S(_04950_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10448_ (.I0(\dp.rf.rf[31][5] ),
    .I1(_04455_),
    .S(_04950_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10449_ (.A1(\dp.rf.rf[31][6] ),
    .A2(_04953_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10450_ (.A1(_04466_),
    .A2(_04953_),
    .B(_04964_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10451_ (.I0(\dp.rf.rf[31][7] ),
    .I1(_04473_),
    .S(_04950_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10452_ (.A1(\dp.rf.rf[31][8] ),
    .A2(_04953_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10453_ (.A1(_04485_),
    .A2(_04953_),
    .B(_04965_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10454_ (.I0(\dp.rf.rf[31][9] ),
    .I1(_04497_),
    .S(_04950_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10455_ (.A1(_04499_),
    .A2(_04532_),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input27 (.I(instr[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input26 (.I(instr[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10458_ (.I0(\dp.rf.rf[3][0] ),
    .I1(net478),
    .S(_04966_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10459_ (.I0(\dp.rf.rf[3][10] ),
    .I1(_04069_),
    .S(_04966_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10460_ (.I0(\dp.rf.rf[3][11] ),
    .I1(_04092_),
    .S(_04966_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10461_ (.I0(\dp.rf.rf[3][12] ),
    .I1(_04106_),
    .S(_04966_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10462_ (.I0(\dp.rf.rf[3][13] ),
    .I1(_04119_),
    .S(_04966_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10463_ (.I0(\dp.rf.rf[3][14] ),
    .I1(_04136_),
    .S(_04966_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10464_ (.I0(\dp.rf.rf[3][15] ),
    .I1(_04152_),
    .S(_04966_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10465_ (.A1(_04499_),
    .A2(_04532_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input25 (.I(instr[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10467_ (.A1(\dp.rf.rf[3][16] ),
    .A2(_04969_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10468_ (.A1(_04178_),
    .A2(_04969_),
    .B(_04971_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10469_ (.I0(\dp.rf.rf[3][17] ),
    .I1(net483),
    .S(_04966_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10470_ (.I0(\dp.rf.rf[3][18] ),
    .I1(net482),
    .S(_04966_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10471_ (.I0(\dp.rf.rf[3][19] ),
    .I1(_04222_),
    .S(_04966_),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 input24 (.I(instr[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10473_ (.I0(\dp.rf.rf[3][1] ),
    .I1(_04228_),
    .S(_04966_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10474_ (.A1(\dp.rf.rf[3][20] ),
    .A2(_04969_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10475_ (.A1(_04250_),
    .A2(_04969_),
    .B(_04973_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10476_ (.I0(\dp.rf.rf[3][21] ),
    .I1(_04267_),
    .S(_04966_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10477_ (.I0(\dp.rf.rf[3][22] ),
    .I1(net481),
    .S(_04966_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10478_ (.A1(_04301_),
    .A2(_04966_),
    .Z(_04974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10479_ (.A1(_01835_),
    .A2(_04969_),
    .B1(_04974_),
    .B2(net485),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10480_ (.I0(\dp.rf.rf[3][24] ),
    .I1(_04314_),
    .S(_04966_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10481_ (.I(\dp.rf.rf[3][25] ),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10482_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04966_),
    .Z(_04976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10483_ (.A1(_04975_),
    .A2(_04969_),
    .B1(_04976_),
    .B2(_04325_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10484_ (.I0(\dp.rf.rf[3][26] ),
    .I1(_04343_),
    .S(_04966_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10485_ (.I0(\dp.rf.rf[3][27] ),
    .I1(_04355_),
    .S(_04966_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10486_ (.I0(\dp.rf.rf[3][28] ),
    .I1(_04370_),
    .S(_04966_),
    .Z(_00823_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10487_ (.I(\dp.rf.rf[3][29] ),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10488_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04966_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10489_ (.A1(_04977_),
    .A2(_04969_),
    .B1(_04978_),
    .B2(net480),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10490_ (.I0(\dp.rf.rf[3][2] ),
    .I1(_04396_),
    .S(_04966_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10491_ (.I0(\dp.rf.rf[3][30] ),
    .I1(net477),
    .S(_04966_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10492_ (.A1(_04429_),
    .A2(_04966_),
    .Z(_04979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10493_ (.A1(_01234_),
    .A2(_04969_),
    .B1(_04979_),
    .B2(net479),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10494_ (.I0(\dp.rf.rf[3][3] ),
    .I1(_04436_),
    .S(_04966_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10495_ (.I0(\dp.rf.rf[3][4] ),
    .I1(_04446_),
    .S(_04966_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10496_ (.I0(\dp.rf.rf[3][5] ),
    .I1(_04455_),
    .S(_04966_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10497_ (.A1(\dp.rf.rf[3][6] ),
    .A2(_04969_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10498_ (.A1(_04466_),
    .A2(_04969_),
    .B(_04980_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10499_ (.I0(\dp.rf.rf[3][7] ),
    .I1(_04473_),
    .S(_04966_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10500_ (.A1(\dp.rf.rf[3][8] ),
    .A2(_04969_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10501_ (.A1(_04485_),
    .A2(_04969_),
    .B(_04981_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10502_ (.I0(\dp.rf.rf[3][9] ),
    .I1(_04497_),
    .S(_04966_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _10503_ (.A1(net3),
    .A2(net2),
    .A3(_04027_),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input23 (.I(instr[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10505_ (.A1(_04608_),
    .A2(_04982_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input22 (.I(instr[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10507_ (.I0(\dp.rf.rf[4][0] ),
    .I1(net478),
    .S(net491),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10508_ (.I0(\dp.rf.rf[4][10] ),
    .I1(_04069_),
    .S(net491),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10509_ (.I0(\dp.rf.rf[4][11] ),
    .I1(_04092_),
    .S(net491),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10510_ (.I0(\dp.rf.rf[4][12] ),
    .I1(_04106_),
    .S(net491),
    .Z(_00838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10511_ (.I0(\dp.rf.rf[4][13] ),
    .I1(_04119_),
    .S(net491),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10512_ (.I0(\dp.rf.rf[4][14] ),
    .I1(_04136_),
    .S(net491),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10513_ (.I0(\dp.rf.rf[4][15] ),
    .I1(_04152_),
    .S(net491),
    .Z(_00841_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10514_ (.A1(_04608_),
    .A2(_04982_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input21 (.I(instr[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10516_ (.A1(\dp.rf.rf[4][16] ),
    .A2(_04986_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10517_ (.A1(_04178_),
    .A2(_04986_),
    .B(_04988_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10518_ (.I0(\dp.rf.rf[4][17] ),
    .I1(net483),
    .S(net491),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10519_ (.I0(\dp.rf.rf[4][18] ),
    .I1(net482),
    .S(net491),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10520_ (.I0(\dp.rf.rf[4][19] ),
    .I1(_04222_),
    .S(net491),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input20 (.I(instr[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10522_ (.I0(\dp.rf.rf[4][1] ),
    .I1(_04228_),
    .S(_04984_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10523_ (.A1(\dp.rf.rf[4][20] ),
    .A2(_04986_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10524_ (.A1(_04250_),
    .A2(_04986_),
    .B(_04990_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10525_ (.I0(\dp.rf.rf[4][21] ),
    .I1(_04267_),
    .S(_04984_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10526_ (.I0(\dp.rf.rf[4][22] ),
    .I1(net481),
    .S(_04984_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10527_ (.I(\dp.rf.rf[4][23] ),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10528_ (.A1(_04301_),
    .A2(_04984_),
    .Z(_04992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10529_ (.A1(_04991_),
    .A2(_04986_),
    .B1(_04992_),
    .B2(net485),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10530_ (.I0(\dp.rf.rf[4][24] ),
    .I1(_04314_),
    .S(_04984_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10531_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04984_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10532_ (.A1(_01707_),
    .A2(_04986_),
    .B1(_04993_),
    .B2(_04325_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10533_ (.I0(\dp.rf.rf[4][26] ),
    .I1(_04343_),
    .S(_04984_),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10534_ (.I0(\dp.rf.rf[4][27] ),
    .I1(_04355_),
    .S(_04984_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10535_ (.I0(\dp.rf.rf[4][28] ),
    .I1(_04370_),
    .S(_04984_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10536_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04984_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10537_ (.A1(_01450_),
    .A2(_04986_),
    .B1(_04994_),
    .B2(net480),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10538_ (.I0(\dp.rf.rf[4][2] ),
    .I1(_04396_),
    .S(_04984_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10539_ (.I0(\dp.rf.rf[4][30] ),
    .I1(net477),
    .S(_04984_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10540_ (.A1(_04429_),
    .A2(_04984_),
    .Z(_04995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10541_ (.A1(_01244_),
    .A2(_04986_),
    .B1(_04995_),
    .B2(net479),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10542_ (.I0(\dp.rf.rf[4][3] ),
    .I1(_04436_),
    .S(net491),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10543_ (.I0(\dp.rf.rf[4][4] ),
    .I1(_04446_),
    .S(_04984_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10544_ (.I0(\dp.rf.rf[4][5] ),
    .I1(_04455_),
    .S(net491),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10545_ (.A1(\dp.rf.rf[4][6] ),
    .A2(_04986_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10546_ (.A1(_04466_),
    .A2(_04986_),
    .B(_04996_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10547_ (.I0(\dp.rf.rf[4][7] ),
    .I1(_04473_),
    .S(net491),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10548_ (.A1(\dp.rf.rf[4][8] ),
    .A2(_04986_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10549_ (.A1(_04485_),
    .A2(_04986_),
    .B(_04997_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10550_ (.I0(\dp.rf.rf[4][9] ),
    .I1(_04497_),
    .S(_04984_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10551_ (.A1(_04625_),
    .A2(_04982_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input19 (.I(instr[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10553_ (.I0(\dp.rf.rf[5][0] ),
    .I1(net478),
    .S(net490),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10554_ (.I0(\dp.rf.rf[5][10] ),
    .I1(_04069_),
    .S(net490),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10555_ (.I0(\dp.rf.rf[5][11] ),
    .I1(_04092_),
    .S(net490),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10556_ (.I0(\dp.rf.rf[5][12] ),
    .I1(_04106_),
    .S(net490),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10557_ (.I0(\dp.rf.rf[5][13] ),
    .I1(_04119_),
    .S(net490),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10558_ (.I0(\dp.rf.rf[5][14] ),
    .I1(_04136_),
    .S(net490),
    .Z(_00872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10559_ (.I0(\dp.rf.rf[5][15] ),
    .I1(_04152_),
    .S(net490),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10560_ (.A1(_04625_),
    .A2(_04982_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input18 (.I(instr[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10562_ (.A1(\dp.rf.rf[5][16] ),
    .A2(_05000_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10563_ (.A1(_04178_),
    .A2(_05000_),
    .B(_05002_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10564_ (.I0(\dp.rf.rf[5][17] ),
    .I1(net483),
    .S(net490),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10565_ (.I0(\dp.rf.rf[5][18] ),
    .I1(net482),
    .S(net490),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10566_ (.I0(\dp.rf.rf[5][19] ),
    .I1(_04222_),
    .S(net490),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input17 (.I(instr[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10568_ (.I0(\dp.rf.rf[5][1] ),
    .I1(_04228_),
    .S(_04998_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10569_ (.A1(\dp.rf.rf[5][20] ),
    .A2(_05000_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10570_ (.A1(_04250_),
    .A2(_05000_),
    .B(_05004_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10571_ (.I0(\dp.rf.rf[5][21] ),
    .I1(_04267_),
    .S(_04998_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10572_ (.I0(\dp.rf.rf[5][22] ),
    .I1(net481),
    .S(_04998_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10573_ (.I(\dp.rf.rf[5][23] ),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10574_ (.A1(_04301_),
    .A2(_04998_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10575_ (.A1(_05005_),
    .A2(_05000_),
    .B1(_05006_),
    .B2(net485),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10576_ (.I0(\dp.rf.rf[5][24] ),
    .I1(_04314_),
    .S(_04998_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10577_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_04998_),
    .Z(_05007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10578_ (.A1(_01709_),
    .A2(_05000_),
    .B1(_05007_),
    .B2(_04325_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10579_ (.I0(\dp.rf.rf[5][26] ),
    .I1(_04343_),
    .S(_04998_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10580_ (.I0(\dp.rf.rf[5][27] ),
    .I1(_04355_),
    .S(_04998_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10581_ (.I0(\dp.rf.rf[5][28] ),
    .I1(_04370_),
    .S(_04998_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10582_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_04998_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10583_ (.A1(_01453_),
    .A2(_05000_),
    .B1(_05008_),
    .B2(net480),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10584_ (.I0(\dp.rf.rf[5][2] ),
    .I1(_04396_),
    .S(_04998_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10585_ (.I0(\dp.rf.rf[5][30] ),
    .I1(net477),
    .S(_04998_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10586_ (.A1(_04429_),
    .A2(_04998_),
    .Z(_05009_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10587_ (.A1(_01247_),
    .A2(_05000_),
    .B1(_05009_),
    .B2(net479),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10588_ (.I0(\dp.rf.rf[5][3] ),
    .I1(_04436_),
    .S(net490),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10589_ (.I0(\dp.rf.rf[5][4] ),
    .I1(_04446_),
    .S(_04998_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10590_ (.I0(\dp.rf.rf[5][5] ),
    .I1(_04455_),
    .S(net490),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10591_ (.A1(\dp.rf.rf[5][6] ),
    .A2(_05000_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10592_ (.A1(_04466_),
    .A2(_05000_),
    .B(_05010_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10593_ (.I0(\dp.rf.rf[5][7] ),
    .I1(_04473_),
    .S(net490),
    .Z(_00896_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10594_ (.A1(\dp.rf.rf[5][8] ),
    .A2(_05000_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10595_ (.A1(_04485_),
    .A2(_05000_),
    .B(_05011_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10596_ (.I0(\dp.rf.rf[5][9] ),
    .I1(_04497_),
    .S(_04998_),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10597_ (.A1(_04640_),
    .A2(_04982_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input16 (.I(instr[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10599_ (.I0(\dp.rf.rf[6][0] ),
    .I1(net478),
    .S(net489),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10600_ (.I0(\dp.rf.rf[6][10] ),
    .I1(_04069_),
    .S(net489),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10601_ (.I0(\dp.rf.rf[6][11] ),
    .I1(_04092_),
    .S(net489),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10602_ (.I0(\dp.rf.rf[6][12] ),
    .I1(_04106_),
    .S(net489),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10603_ (.I0(\dp.rf.rf[6][13] ),
    .I1(_04119_),
    .S(net489),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10604_ (.I0(\dp.rf.rf[6][14] ),
    .I1(_04136_),
    .S(net489),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10605_ (.I0(\dp.rf.rf[6][15] ),
    .I1(_04152_),
    .S(net489),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10606_ (.A1(_04640_),
    .A2(_04982_),
    .Z(_05014_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input15 (.I(instr[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10608_ (.A1(\dp.rf.rf[6][16] ),
    .A2(_05014_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10609_ (.A1(_04178_),
    .A2(_05014_),
    .B(_05016_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10610_ (.I0(\dp.rf.rf[6][17] ),
    .I1(net483),
    .S(net489),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10611_ (.I0(\dp.rf.rf[6][18] ),
    .I1(net482),
    .S(net489),
    .Z(_00908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10612_ (.I0(\dp.rf.rf[6][19] ),
    .I1(_04222_),
    .S(net489),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input14 (.I(instr[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10614_ (.I0(\dp.rf.rf[6][1] ),
    .I1(_04228_),
    .S(_05012_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10615_ (.A1(\dp.rf.rf[6][20] ),
    .A2(_05014_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10616_ (.A1(_04250_),
    .A2(_05014_),
    .B(_05018_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10617_ (.I0(\dp.rf.rf[6][21] ),
    .I1(_04267_),
    .S(_05012_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10618_ (.I0(\dp.rf.rf[6][22] ),
    .I1(net481),
    .S(_05012_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10619_ (.A1(_04301_),
    .A2(_05012_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10620_ (.A1(_01836_),
    .A2(_05014_),
    .B1(_05019_),
    .B2(net485),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10621_ (.I0(\dp.rf.rf[6][24] ),
    .I1(_04314_),
    .S(_05012_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10622_ (.I(\dp.rf.rf[6][25] ),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10623_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_05012_),
    .Z(_05021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10624_ (.A1(_05020_),
    .A2(_05014_),
    .B1(_05021_),
    .B2(_04325_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10625_ (.I0(\dp.rf.rf[6][26] ),
    .I1(_04343_),
    .S(_05012_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10626_ (.I0(\dp.rf.rf[6][27] ),
    .I1(_04355_),
    .S(_05012_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10627_ (.I0(\dp.rf.rf[6][28] ),
    .I1(_04370_),
    .S(_05012_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10628_ (.I(\dp.rf.rf[6][29] ),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10629_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_05012_),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10630_ (.A1(_05022_),
    .A2(_05014_),
    .B1(_05023_),
    .B2(net480),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10631_ (.I0(\dp.rf.rf[6][2] ),
    .I1(_04396_),
    .S(_05012_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10632_ (.I0(\dp.rf.rf[6][30] ),
    .I1(net477),
    .S(_05012_),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10633_ (.A1(_04429_),
    .A2(_05012_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10634_ (.A1(_01238_),
    .A2(_05014_),
    .B1(_05024_),
    .B2(net479),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10635_ (.I0(\dp.rf.rf[6][3] ),
    .I1(_04436_),
    .S(net489),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10636_ (.I0(\dp.rf.rf[6][4] ),
    .I1(_04446_),
    .S(_05012_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10637_ (.I0(\dp.rf.rf[6][5] ),
    .I1(_04455_),
    .S(net489),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10638_ (.A1(\dp.rf.rf[6][6] ),
    .A2(_05014_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10639_ (.A1(_04466_),
    .A2(_05014_),
    .B(_05025_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10640_ (.I0(\dp.rf.rf[6][7] ),
    .I1(_04473_),
    .S(net489),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10641_ (.A1(\dp.rf.rf[6][8] ),
    .A2(_05014_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10642_ (.A1(_04485_),
    .A2(_05014_),
    .B(_05026_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10643_ (.I0(\dp.rf.rf[6][9] ),
    .I1(_04497_),
    .S(_05012_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _10644_ (.A1(_04655_),
    .A2(_04982_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input13 (.I(instr[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10646_ (.I0(\dp.rf.rf[7][0] ),
    .I1(net478),
    .S(net488),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10647_ (.I0(\dp.rf.rf[7][10] ),
    .I1(_04069_),
    .S(net488),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10648_ (.I0(\dp.rf.rf[7][11] ),
    .I1(_04092_),
    .S(net488),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10649_ (.I0(\dp.rf.rf[7][12] ),
    .I1(_04106_),
    .S(net488),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10650_ (.I0(\dp.rf.rf[7][13] ),
    .I1(_04119_),
    .S(net488),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10651_ (.I0(\dp.rf.rf[7][14] ),
    .I1(_04136_),
    .S(net488),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10652_ (.I0(\dp.rf.rf[7][15] ),
    .I1(_04152_),
    .S(net488),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _10653_ (.A1(_04655_),
    .A2(_04982_),
    .Z(_05029_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(instr[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10655_ (.A1(\dp.rf.rf[7][16] ),
    .A2(_05029_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10656_ (.A1(_04178_),
    .A2(_05029_),
    .B(_05031_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10657_ (.I0(\dp.rf.rf[7][17] ),
    .I1(net483),
    .S(net488),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10658_ (.I0(\dp.rf.rf[7][18] ),
    .I1(net482),
    .S(net488),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10659_ (.I0(\dp.rf.rf[7][19] ),
    .I1(_04222_),
    .S(net488),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 input11 (.I(instr[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10661_ (.I0(\dp.rf.rf[7][1] ),
    .I1(_04228_),
    .S(_05027_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10662_ (.A1(\dp.rf.rf[7][20] ),
    .A2(_05029_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10663_ (.A1(_04250_),
    .A2(_05029_),
    .B(_05033_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10664_ (.I0(\dp.rf.rf[7][21] ),
    .I1(_04267_),
    .S(_05027_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10665_ (.I0(\dp.rf.rf[7][22] ),
    .I1(net481),
    .S(_05027_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10666_ (.A1(_04301_),
    .A2(_05027_),
    .Z(_05034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10667_ (.A1(_01837_),
    .A2(_05029_),
    .B1(_05034_),
    .B2(net485),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10668_ (.I0(\dp.rf.rf[7][24] ),
    .I1(_04314_),
    .S(_05027_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10669_ (.I(\dp.rf.rf[7][25] ),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10670_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_05027_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10671_ (.A1(_05035_),
    .A2(_05029_),
    .B1(_05036_),
    .B2(_04325_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10672_ (.I0(\dp.rf.rf[7][26] ),
    .I1(_04343_),
    .S(_05027_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10673_ (.I0(\dp.rf.rf[7][27] ),
    .I1(_04355_),
    .S(_05027_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10674_ (.I0(\dp.rf.rf[7][28] ),
    .I1(_04370_),
    .S(_05027_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10675_ (.I(\dp.rf.rf[7][29] ),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10676_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_05027_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10677_ (.A1(_05037_),
    .A2(_05029_),
    .B1(_05038_),
    .B2(net480),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10678_ (.I0(\dp.rf.rf[7][2] ),
    .I1(_04396_),
    .S(_05027_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10679_ (.I0(\dp.rf.rf[7][30] ),
    .I1(net477),
    .S(_05027_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10680_ (.A1(_04429_),
    .A2(_05027_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10681_ (.A1(_01236_),
    .A2(_05029_),
    .B1(_05039_),
    .B2(net479),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10682_ (.I0(\dp.rf.rf[7][3] ),
    .I1(_04436_),
    .S(net488),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10683_ (.I0(\dp.rf.rf[7][4] ),
    .I1(_04446_),
    .S(_05027_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10684_ (.I0(\dp.rf.rf[7][5] ),
    .I1(_04455_),
    .S(net488),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10685_ (.A1(\dp.rf.rf[7][6] ),
    .A2(_05029_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10686_ (.A1(_04466_),
    .A2(_05029_),
    .B(_05040_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10687_ (.I0(\dp.rf.rf[7][7] ),
    .I1(_04473_),
    .S(net488),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10688_ (.A1(\dp.rf.rf[7][8] ),
    .A2(_05029_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10689_ (.A1(_04485_),
    .A2(_05029_),
    .B(_05041_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10690_ (.I0(\dp.rf.rf[7][9] ),
    .I1(_04497_),
    .S(_05027_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10691_ (.A1(_04029_),
    .A2(_04533_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 input10 (.I(instr[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input9 (.I(instr[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10694_ (.I0(\dp.rf.rf[8][0] ),
    .I1(net478),
    .S(_05042_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10695_ (.I0(\dp.rf.rf[8][10] ),
    .I1(_04069_),
    .S(_05042_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10696_ (.I0(\dp.rf.rf[8][11] ),
    .I1(_04092_),
    .S(_05042_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10697_ (.I0(\dp.rf.rf[8][12] ),
    .I1(_04106_),
    .S(_05042_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10698_ (.I0(\dp.rf.rf[8][13] ),
    .I1(_04119_),
    .S(_05042_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10699_ (.I0(\dp.rf.rf[8][14] ),
    .I1(_04136_),
    .S(_05042_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10700_ (.I0(\dp.rf.rf[8][15] ),
    .I1(_04152_),
    .S(_05042_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10701_ (.A1(_04029_),
    .A2(_04533_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input8 (.I(instr[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10703_ (.A1(\dp.rf.rf[8][16] ),
    .A2(_05045_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10704_ (.A1(_04178_),
    .A2(_05045_),
    .B(_05047_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10705_ (.I0(\dp.rf.rf[8][17] ),
    .I1(net483),
    .S(_05042_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10706_ (.I0(\dp.rf.rf[8][18] ),
    .I1(net482),
    .S(_05042_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10707_ (.I0(\dp.rf.rf[8][19] ),
    .I1(_04222_),
    .S(_05042_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input7 (.I(instr[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10709_ (.I0(\dp.rf.rf[8][1] ),
    .I1(_04228_),
    .S(_05042_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10710_ (.A1(\dp.rf.rf[8][20] ),
    .A2(_05045_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10711_ (.A1(_04250_),
    .A2(_05045_),
    .B(_05049_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10712_ (.I0(\dp.rf.rf[8][21] ),
    .I1(_04267_),
    .S(_05042_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10713_ (.I0(\dp.rf.rf[8][22] ),
    .I1(net481),
    .S(_05042_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10714_ (.I(\dp.rf.rf[8][23] ),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10715_ (.A1(_04301_),
    .A2(_05042_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10716_ (.A1(_05050_),
    .A2(_05045_),
    .B1(_05051_),
    .B2(net485),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10717_ (.I0(\dp.rf.rf[8][24] ),
    .I1(_04314_),
    .S(_05042_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10718_ (.I(\dp.rf.rf[8][25] ),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10719_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_05042_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10720_ (.A1(_05052_),
    .A2(_05045_),
    .B1(_05053_),
    .B2(_04325_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10721_ (.I0(\dp.rf.rf[8][26] ),
    .I1(_04343_),
    .S(_05042_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10722_ (.I0(\dp.rf.rf[8][27] ),
    .I1(_04355_),
    .S(_05042_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10723_ (.I0(\dp.rf.rf[8][28] ),
    .I1(_04370_),
    .S(_05042_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10724_ (.I(\dp.rf.rf[8][29] ),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10725_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_05042_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10726_ (.A1(_05054_),
    .A2(_05045_),
    .B1(_05055_),
    .B2(net480),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10727_ (.I0(\dp.rf.rf[8][2] ),
    .I1(_04396_),
    .S(_05042_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10728_ (.I0(\dp.rf.rf[8][30] ),
    .I1(net477),
    .S(_05042_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10729_ (.I(\dp.rf.rf[8][31] ),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10730_ (.A1(_04429_),
    .A2(_05042_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10731_ (.A1(_05056_),
    .A2(_05045_),
    .B1(_05057_),
    .B2(net479),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10732_ (.I0(\dp.rf.rf[8][3] ),
    .I1(_04436_),
    .S(_05042_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10733_ (.I0(\dp.rf.rf[8][4] ),
    .I1(_04446_),
    .S(_05042_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10734_ (.I0(\dp.rf.rf[8][5] ),
    .I1(_04455_),
    .S(_05042_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10735_ (.A1(\dp.rf.rf[8][6] ),
    .A2(_05045_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10736_ (.A1(_04466_),
    .A2(_05045_),
    .B(_05058_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10737_ (.I0(\dp.rf.rf[8][7] ),
    .I1(_04473_),
    .S(_05042_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10738_ (.A1(\dp.rf.rf[8][8] ),
    .A2(_05045_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10739_ (.A1(_04485_),
    .A2(_05045_),
    .B(_05059_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10740_ (.I0(\dp.rf.rf[8][9] ),
    .I1(_04497_),
    .S(_05042_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10741_ (.A1(_04029_),
    .A2(_04552_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input6 (.I(instr[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input5 (.I(instr[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10744_ (.I0(\dp.rf.rf[9][0] ),
    .I1(net478),
    .S(_05060_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10745_ (.I0(\dp.rf.rf[9][10] ),
    .I1(_04069_),
    .S(_05060_),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10746_ (.I0(\dp.rf.rf[9][11] ),
    .I1(_04092_),
    .S(_05060_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10747_ (.I0(\dp.rf.rf[9][12] ),
    .I1(_04106_),
    .S(_05060_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10748_ (.I0(\dp.rf.rf[9][13] ),
    .I1(_04119_),
    .S(_05060_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10749_ (.I0(\dp.rf.rf[9][14] ),
    .I1(_04136_),
    .S(_05060_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10750_ (.I0(\dp.rf.rf[9][15] ),
    .I1(_04152_),
    .S(_05060_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10751_ (.A1(_04029_),
    .A2(_04552_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input4 (.I(instr[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10753_ (.A1(\dp.rf.rf[9][16] ),
    .A2(_05063_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10754_ (.A1(_04178_),
    .A2(_05063_),
    .B(_05065_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10755_ (.I0(\dp.rf.rf[9][17] ),
    .I1(net483),
    .S(_05060_),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10756_ (.I0(\dp.rf.rf[9][18] ),
    .I1(net482),
    .S(_05060_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10757_ (.I0(\dp.rf.rf[9][19] ),
    .I1(_04222_),
    .S(_05060_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input3 (.I(instr[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10759_ (.I0(\dp.rf.rf[9][1] ),
    .I1(_04228_),
    .S(_05060_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10760_ (.A1(\dp.rf.rf[9][20] ),
    .A2(_05063_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10761_ (.A1(_04250_),
    .A2(_05063_),
    .B(_05067_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10762_ (.I0(\dp.rf.rf[9][21] ),
    .I1(_04267_),
    .S(_05060_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10763_ (.I0(\dp.rf.rf[9][22] ),
    .I1(net481),
    .S(_05060_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10764_ (.I(\dp.rf.rf[9][23] ),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10765_ (.A1(_04301_),
    .A2(_05060_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10766_ (.A1(_05068_),
    .A2(_05063_),
    .B1(_05069_),
    .B2(net485),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10767_ (.I0(\dp.rf.rf[9][24] ),
    .I1(_04314_),
    .S(_05060_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10768_ (.I(\dp.rf.rf[9][25] ),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10769_ (.A1(_04327_),
    .A2(_04329_),
    .A3(_05060_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10770_ (.A1(_05070_),
    .A2(_05063_),
    .B1(_05071_),
    .B2(_04325_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10771_ (.I0(\dp.rf.rf[9][26] ),
    .I1(_04343_),
    .S(_05060_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10772_ (.I0(\dp.rf.rf[9][27] ),
    .I1(_04355_),
    .S(_05060_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10773_ (.I0(\dp.rf.rf[9][28] ),
    .I1(_04370_),
    .S(_05060_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10774_ (.I(\dp.rf.rf[9][29] ),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10775_ (.A1(_04388_),
    .A2(_04390_),
    .A3(_05060_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10776_ (.A1(_05072_),
    .A2(_05063_),
    .B1(_05073_),
    .B2(net480),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10777_ (.I0(\dp.rf.rf[9][2] ),
    .I1(_04396_),
    .S(_05060_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10778_ (.I0(\dp.rf.rf[9][30] ),
    .I1(net477),
    .S(_05060_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _10779_ (.I(\dp.rf.rf[9][31] ),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10780_ (.A1(_04429_),
    .A2(_05060_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _10781_ (.A1(_05074_),
    .A2(_05063_),
    .B1(_05075_),
    .B2(net479),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10782_ (.I0(\dp.rf.rf[9][3] ),
    .I1(_04436_),
    .S(_05060_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10783_ (.I0(\dp.rf.rf[9][4] ),
    .I1(_04446_),
    .S(_05060_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10784_ (.I0(\dp.rf.rf[9][5] ),
    .I1(_04455_),
    .S(_05060_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10785_ (.A1(\dp.rf.rf[9][6] ),
    .A2(_05063_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10786_ (.A1(_04466_),
    .A2(_05063_),
    .B(_05076_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10787_ (.I0(\dp.rf.rf[9][7] ),
    .I1(_04473_),
    .S(_05060_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10788_ (.A1(\dp.rf.rf[9][8] ),
    .A2(_05063_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10789_ (.A1(_04485_),
    .A2(_05063_),
    .B(_05077_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10790_ (.I0(\dp.rf.rf[9][9] ),
    .I1(_04497_),
    .S(_05060_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input2 (.I(instr[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10792_ (.A1(_04269_),
    .A2(net487),
    .A3(_04068_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10793_ (.A1(net486),
    .A2(_04063_),
    .B(_05079_),
    .ZN(\dp.ISRmux.d0[10] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10794_ (.I0(_04090_),
    .I1(_04079_),
    .S(net486),
    .Z(\dp.ISRmux.d0[11] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10795_ (.I0(_04101_),
    .I1(_04103_),
    .S(net486),
    .Z(\dp.ISRmux.d0[12] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10796_ (.I0(_04115_),
    .I1(_04117_),
    .S(net486),
    .Z(\dp.ISRmux.d0[13] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10797_ (.I0(_04131_),
    .I1(_04134_),
    .S(net486),
    .Z(\dp.ISRmux.d0[14] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10798_ (.I0(_04148_),
    .I1(_04150_),
    .S(net486),
    .Z(\dp.ISRmux.d0[15] ));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10799_ (.A1(_04269_),
    .A2(net487),
    .B(_04176_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _10800_ (.A1(_04269_),
    .A2(net487),
    .A3(_04168_),
    .B(_05080_),
    .ZN(\dp.ISRmux.d0[16] ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10801_ (.A1(net486),
    .A2(_04197_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10802_ (.A1(net486),
    .A2(_04193_),
    .B(_05081_),
    .ZN(\dp.ISRmux.d0[17] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10803_ (.I0(_04209_),
    .I1(_04204_),
    .S(net486),
    .Z(\dp.ISRmux.d0[18] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10804_ (.I0(_04218_),
    .I1(_04220_),
    .S(net486),
    .Z(\dp.ISRmux.d0[19] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10805_ (.A1(_04269_),
    .A2(_04013_),
    .A3(_04236_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10806_ (.A1(net486),
    .A2(_04248_),
    .B(_05082_),
    .ZN(\dp.ISRmux.d0[20] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10807_ (.I0(_04265_),
    .I1(_04256_),
    .S(net486),
    .Z(\dp.ISRmux.d0[21] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(instr[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10809_ (.I0(_04278_),
    .I1(_04271_),
    .S(net486),
    .Z(\dp.ISRmux.d0[22] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10810_ (.I0(_04295_),
    .I1(_04288_),
    .S(net486),
    .Z(\dp.ISRmux.d0[23] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10811_ (.A1(_04269_),
    .A2(_04013_),
    .A3(_04305_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10812_ (.A1(net486),
    .A2(_04309_),
    .B(_05084_),
    .ZN(\dp.ISRmux.d0[24] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10813_ (.I0(_04323_),
    .I1(_04318_),
    .S(net486),
    .Z(\dp.ISRmux.d0[25] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10814_ (.I0(_04334_),
    .I1(_04339_),
    .S(net486),
    .Z(\dp.ISRmux.d0[26] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10815_ (.I0(_04353_),
    .I1(_04349_),
    .S(net486),
    .Z(\dp.ISRmux.d0[27] ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _10816_ (.A1(net486),
    .A2(_04364_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10817_ (.A1(net486),
    .A2(_04360_),
    .B(_05085_),
    .ZN(\dp.ISRmux.d0[28] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10818_ (.I0(_04382_),
    .I1(_04375_),
    .S(net486),
    .Z(\dp.ISRmux.d0[29] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10819_ (.I0(_04392_),
    .I1(_04393_),
    .S(net486),
    .Z(\dp.ISRmux.d0[2] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10820_ (.A1(_04269_),
    .A2(net487),
    .A3(_04400_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10821_ (.A1(net486),
    .A2(_04406_),
    .B(_05086_),
    .ZN(\dp.ISRmux.d0[30] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10822_ (.I0(_04423_),
    .I1(_04416_),
    .S(net486),
    .Z(\dp.ISRmux.d0[31] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10823_ (.I0(_04433_),
    .I1(_05371_[0]),
    .S(net486),
    .Z(\dp.ISRmux.d0[3] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10824_ (.A1(_04269_),
    .A2(net487),
    .A3(_04440_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10825_ (.A1(net486),
    .A2(_04444_),
    .B(_05087_),
    .ZN(\dp.ISRmux.d0[4] ));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _10826_ (.A1(_04269_),
    .A2(net487),
    .A3(_04451_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _10827_ (.A1(net486),
    .A2(_04453_),
    .B(_05088_),
    .ZN(\dp.ISRmux.d0[5] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10828_ (.I0(_04462_),
    .I1(_04457_),
    .S(net486),
    .Z(\dp.ISRmux.d0[6] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10829_ (.I0(_04469_),
    .I1(_04471_),
    .S(net486),
    .Z(\dp.ISRmux.d0[7] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10830_ (.I0(_04483_),
    .I1(_04480_),
    .S(net486),
    .Z(\dp.ISRmux.d0[8] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10831_ (.I0(_04495_),
    .I1(_04490_),
    .S(net486),
    .Z(\dp.ISRmux.d0[9] ));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _10832_ (.A1(net27),
    .A2(_02383_),
    .A3(_01115_),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _10833_ (.A1(_01098_),
    .A2(_01089_),
    .A3(net99),
    .A4(_01092_),
    .Z(_05089_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _10834_ (.A1(_01095_),
    .A2(_05089_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10835_ (.A1(_02443_),
    .A2(_05090_),
    .ZN(net134));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10836_ (.A1(_02402_),
    .A2(_05090_),
    .ZN(net135));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _10837_ (.A1(_01095_),
    .A2(_05089_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10838_ (.A1(_02343_),
    .A2(_05091_),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10839_ (.A1(_02297_),
    .A2(_05091_),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10840_ (.A1(_02255_),
    .A2(_05091_),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10841_ (.A1(_03938_),
    .A2(_05091_),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10842_ (.A1(_02164_),
    .A2(_05089_),
    .ZN(net140));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10843_ (.A1(_02112_),
    .A2(_05089_),
    .ZN(net141));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _10844_ (.A1(net29),
    .A2(net5),
    .A3(_01033_),
    .A4(_02902_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10845_ (.A1(_03876_),
    .A2(_05092_),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10846_ (.A1(_03878_),
    .A2(_05092_),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10847_ (.A1(_01965_),
    .A2(_05092_),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10848_ (.A1(_01916_),
    .A2(_05089_),
    .ZN(net146));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10849_ (.A1(_01868_),
    .A2(_05089_),
    .ZN(net147));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10850_ (.A1(_01820_),
    .A2(_05092_),
    .Z(net148));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10851_ (.A1(_01743_),
    .A2(_05092_),
    .Z(net149));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10852_ (.A1(_01693_),
    .A2(_05092_),
    .Z(net150));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10853_ (.A1(_01626_),
    .A2(_05092_),
    .Z(net151));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10854_ (.A1(_01566_),
    .A2(_05089_),
    .ZN(net152));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10855_ (.A1(_01500_),
    .A2(_05092_),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10856_ (.A1(_01437_),
    .A2(_05092_),
    .Z(net154));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10857_ (.A1(_01350_),
    .A2(_05092_),
    .Z(net156));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _10858_ (.A1(_01310_),
    .A2(_05089_),
    .ZN(net157));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10859_ (.A1(_02533_),
    .A2(_05091_),
    .Z(net163));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _10860_ (.A1(_02486_),
    .A2(_05091_),
    .Z(net164));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _10861_ (.A(_05093_[0]),
    .B(_02892_),
    .CI(_05095_[0]),
    .CO(_05096_[0]),
    .S(_05097_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _10862_ (.A(_05098_[0]),
    .B(_05099_[0]),
    .CI(_05100_[0]),
    .CO(_05101_[0]),
    .S(_05102_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10863_ (.A(_01230_),
    .B(_05104_[0]),
    .CO(_05105_[0]),
    .S(_05106_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10864_ (.A(_05107_[0]),
    .B(_05108_[0]),
    .CO(_05109_[0]),
    .S(_05110_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10865_ (.A(_05111_[0]),
    .B(_01287_),
    .CO(_05113_[0]),
    .S(_05114_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10866_ (.A(_05115_[0]),
    .B(_01288_),
    .CO(_05117_[0]),
    .S(_05118_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10867_ (.A(_01414_),
    .B(_05120_[0]),
    .CO(_05121_[0]),
    .S(_05122_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10868_ (.A(_05123_[0]),
    .B(_05124_[0]),
    .CO(_05125_[0]),
    .S(_05126_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10869_ (.A(_05127_[0]),
    .B(_05128_[0]),
    .CO(_05129_[0]),
    .S(_05130_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10870_ (.A(_05131_[0]),
    .B(_05132_[0]),
    .CO(_05133_[0]),
    .S(_05134_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10871_ (.A(_05135_[0]),
    .B(_05136_[0]),
    .CO(_05137_[0]),
    .S(_05138_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10872_ (.A(_05139_[0]),
    .B(_05140_[0]),
    .CO(_05141_[0]),
    .S(_05142_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10873_ (.A(_01602_),
    .B(_05144_[0]),
    .CO(_05145_[0]),
    .S(_05146_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10874_ (.A(_05147_[0]),
    .B(_05148_[0]),
    .CO(_05149_[0]),
    .S(_05150_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10875_ (.A(_01657_),
    .B(_05152_[0]),
    .CO(_05153_[0]),
    .S(_05154_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10876_ (.A(_05155_[0]),
    .B(_05156_[0]),
    .CO(_05157_[0]),
    .S(_05158_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10877_ (.A(_05159_[0]),
    .B(_05160_[0]),
    .CO(_05161_[0]),
    .S(_05162_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10878_ (.A(_05163_[0]),
    .B(_05164_[0]),
    .CO(_05165_[0]),
    .S(_05166_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10879_ (.A(_01786_),
    .B(_05168_[0]),
    .CO(_05169_[0]),
    .S(_05170_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10880_ (.A(_05171_[0]),
    .B(_05172_[0]),
    .CO(_05173_[0]),
    .S(_05174_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10881_ (.A(_01852_),
    .B(_05176_[0]),
    .CO(_05177_[0]),
    .S(_05178_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10882_ (.A(_05179_[0]),
    .B(_05180_[0]),
    .CO(_05181_[0]),
    .S(_05182_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10883_ (.A(_01899_),
    .B(_05184_[0]),
    .CO(_05185_[0]),
    .S(_05186_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10884_ (.A(_05187_[0]),
    .B(_05188_[0]),
    .CO(_05189_[0]),
    .S(_05190_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10885_ (.A(_01947_),
    .B(_05192_[0]),
    .CO(_05193_[0]),
    .S(_05194_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10886_ (.A(_05195_[0]),
    .B(_05196_[0]),
    .CO(_05197_[0]),
    .S(_05198_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10887_ (.A(_01997_),
    .B(_05200_[0]),
    .CO(_05201_[0]),
    .S(_05202_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10888_ (.A(_05203_[0]),
    .B(_05204_[0]),
    .CO(_05205_[0]),
    .S(_05206_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10889_ (.A(_02044_),
    .B(_05208_[0]),
    .CO(_05209_[0]),
    .S(_05210_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10890_ (.A(_05211_[0]),
    .B(_05212_[0]),
    .CO(_05213_[0]),
    .S(_05214_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10891_ (.A(_02086_),
    .B(_05216_[0]),
    .CO(_05217_[0]),
    .S(_05218_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10892_ (.A(_05219_[0]),
    .B(_05220_[0]),
    .CO(_05221_[0]),
    .S(_05222_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10893_ (.A(_02142_),
    .B(_05224_[0]),
    .CO(_05225_[0]),
    .S(_05226_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10894_ (.A(_05227_[0]),
    .B(_05228_[0]),
    .CO(_05229_[0]),
    .S(_05230_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10895_ (.A(net508),
    .B(_05232_[0]),
    .CO(_05233_[0]),
    .S(_05234_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10896_ (.A(_05235_[0]),
    .B(_05236_[0]),
    .CO(_05237_[0]),
    .S(_05238_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10897_ (.A(_02236_),
    .B(_05240_[0]),
    .CO(_05241_[0]),
    .S(_05242_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10898_ (.A(_05243_[0]),
    .B(_05244_[0]),
    .CO(_05245_[0]),
    .S(_05246_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10899_ (.A(_02284_),
    .B(_05248_[0]),
    .CO(_05249_[0]),
    .S(_05250_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10900_ (.A(_05251_[0]),
    .B(_05252_[0]),
    .CO(_05253_[0]),
    .S(_05254_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10901_ (.A(_02327_),
    .B(_05256_[0]),
    .CO(_05257_[0]),
    .S(_05258_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10902_ (.A(_05259_[0]),
    .B(_05260_[0]),
    .CO(_05261_[0]),
    .S(_05262_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10903_ (.A(_02382_),
    .B(_05264_[0]),
    .CO(_05265_[0]),
    .S(_05266_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10904_ (.A(_05267_[0]),
    .B(_05268_[0]),
    .CO(_05269_[0]),
    .S(_05270_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10905_ (.A(_02428_),
    .B(_05272_[0]),
    .CO(_05273_[0]),
    .S(_05274_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10906_ (.A(_05275_[0]),
    .B(_05276_[0]),
    .CO(_05277_[0]),
    .S(_05278_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10907_ (.A(_02470_),
    .B(_05280_[0]),
    .CO(_05281_[0]),
    .S(_05282_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10908_ (.A(_05283_[0]),
    .B(_05284_[0]),
    .CO(_05285_[0]),
    .S(_05286_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10909_ (.A(_02518_),
    .B(_05288_[0]),
    .CO(_05289_[0]),
    .S(_05290_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10910_ (.A(_05291_[0]),
    .B(_05292_[0]),
    .CO(_05293_[0]),
    .S(_05294_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10911_ (.A(_02560_),
    .B(_05296_[0]),
    .CO(_05297_[0]),
    .S(_05298_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10912_ (.A(_05299_[0]),
    .B(_05300_[0]),
    .CO(_05301_[0]),
    .S(_05302_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10913_ (.A(_05303_[0]),
    .B(_05304_[0]),
    .CO(_05305_[0]),
    .S(_05306_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10914_ (.A(_05307_[0]),
    .B(_05308_[0]),
    .CO(_05309_[0]),
    .S(_05310_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10915_ (.A(_02645_),
    .B(_05312_[0]),
    .CO(_05313_[0]),
    .S(_05314_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10916_ (.A(_05315_[0]),
    .B(_05316_[0]),
    .CO(_05317_[0]),
    .S(_05318_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10917_ (.A(_02683_),
    .B(_05320_[0]),
    .CO(_05321_[0]),
    .S(_05322_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10918_ (.A(_05323_[0]),
    .B(_05324_[0]),
    .CO(_05325_[0]),
    .S(_05326_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10919_ (.A(net506),
    .B(_05328_[0]),
    .CO(_05329_[0]),
    .S(_05330_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10920_ (.A(_05331_[0]),
    .B(_05332_[0]),
    .CO(_05333_[0]),
    .S(_05334_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10921_ (.A(net501),
    .B(_05336_[0]),
    .CO(_05337_[0]),
    .S(_05338_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10922_ (.A(_05339_[0]),
    .B(_05340_[0]),
    .CO(_05341_[0]),
    .S(_05342_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10923_ (.A(_02828_),
    .B(_05344_[0]),
    .CO(_05345_[0]),
    .S(_05346_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10924_ (.A(_05347_[0]),
    .B(_05348_[0]),
    .CO(_05349_[0]),
    .S(_05350_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10925_ (.A(_02892_),
    .B(_05095_[0]),
    .CO(_05351_[0]),
    .S(_05352_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10926_ (.A(_05353_[0]),
    .B(_05354_[0]),
    .CO(_05355_[0]),
    .S(_05356_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10927_ (.A(_05357_[0]),
    .B(_05358_[0]),
    .CO(_05098_[0]),
    .S(_05359_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10928_ (.A(_05099_[0]),
    .B(_05100_[0]),
    .CO(_05360_[0]),
    .S(_05361_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10929_ (.A(_05362_[0]),
    .B(_05363_[0]),
    .CO(_05364_[0]),
    .S(_05365_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10930_ (.A(_05366_[0]),
    .B(_05367_[0]),
    .CO(_05368_[0]),
    .S(_05369_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10931_ (.A(net122),
    .B(net125),
    .CO(_05370_[0]),
    .S(_05371_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10932_ (.A(_05372_[0]),
    .B(_05373_[0]),
    .CO(_05374_[0]),
    .S(_05375_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10933_ (.A(_05376_[0]),
    .B(_05377_[0]),
    .CO(_05378_[0]),
    .S(_05379_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10934_ (.A(_05380_[0]),
    .B(_05381_[0]),
    .CO(_05382_[0]),
    .S(_05383_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10935_ (.A(_05384_[0]),
    .B(_05385_[0]),
    .CO(_05386_[0]),
    .S(_05387_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10936_ (.A(_05388_[0]),
    .B(_05389_[0]),
    .CO(_05390_[0]),
    .S(_05391_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10937_ (.A(_05392_[0]),
    .B(_05393_[0]),
    .CO(_05394_[0]),
    .S(_05395_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10938_ (.A(_05396_[0]),
    .B(_05397_[0]),
    .CO(_05398_[0]),
    .S(_05399_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10939_ (.A(_05400_[0]),
    .B(_05401_[0]),
    .CO(_05402_[0]),
    .S(_05403_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10940_ (.A(_05404_[0]),
    .B(_05405_[0]),
    .CO(_05406_[0]),
    .S(_05407_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10941_ (.A(_05408_[0]),
    .B(_05409_[0]),
    .CO(_05410_[0]),
    .S(_05411_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10942_ (.A(_05412_[0]),
    .B(_05413_[0]),
    .CO(_05414_[0]),
    .S(_05415_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10943_ (.A(_05416_[0]),
    .B(_05417_[0]),
    .CO(_05418_[0]),
    .S(_05419_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10944_ (.A(_05420_[0]),
    .B(_05421_[0]),
    .CO(_05422_[0]),
    .S(_05423_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10945_ (.A(_05424_[0]),
    .B(_05425_[0]),
    .CO(_05426_[0]),
    .S(_05427_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10946_ (.A(_05428_[0]),
    .B(_05429_[0]),
    .CO(_05430_[0]),
    .S(_05431_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _10947_ (.A(_05432_[0]),
    .B(_05433_[0]),
    .CO(_05434_[0]),
    .S(_05435_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10948_ (.A(_05436_[0]),
    .B(_05437_[0]),
    .CO(_05438_[0]),
    .S(_05439_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10949_ (.A(_05440_[0]),
    .B(_05441_[0]),
    .CO(_05442_[0]),
    .S(_05443_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10950_ (.A(_05444_[0]),
    .B(_05445_[0]),
    .CO(_05446_[0]),
    .S(_05447_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10951_ (.A(_05448_[0]),
    .B(_05449_[0]),
    .CO(_05450_[0]),
    .S(_05451_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10952_ (.A(_05452_[0]),
    .B(_05453_[0]),
    .CO(_05454_[0]),
    .S(_05455_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10953_ (.A(_05456_[0]),
    .B(_05457_[0]),
    .CO(_05458_[0]),
    .S(_05459_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10954_ (.A(_05460_[0]),
    .B(_05461_[0]),
    .CO(_05462_[0]),
    .S(_05463_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10955_ (.A(_05464_[0]),
    .B(_05465_[0]),
    .CO(_05466_[0]),
    .S(_05467_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10956_ (.A(_05468_[0]),
    .B(_05469_[0]),
    .CO(_05470_[0]),
    .S(_05471_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10957_ (.A(_05472_[0]),
    .B(_05473_[0]),
    .CO(_05474_[0]),
    .S(_05475_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _10958_ (.A(_05476_[0]),
    .B(_05477_[0]),
    .CO(_05478_[0]),
    .S(_05479_[0]));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[0]$_DFFE_PP0P_  (.D(_00001_),
    .RN(_00000_),
    .CLK(clknet_6_45__leaf_clk),
    .Q(net100));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[10]$_DFF_PP0_  (.D(\dp.ISRmux.d0[10] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net101));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[11]$_DFF_PP0_  (.D(\dp.ISRmux.d0[11] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net102));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[12]$_DFF_PP0_  (.D(\dp.ISRmux.d0[12] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net103));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[13]$_DFF_PP0_  (.D(\dp.ISRmux.d0[13] ),
    .RN(_00000_),
    .CLK(clknet_6_41__leaf_clk),
    .Q(net104));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[14]$_DFF_PP0_  (.D(\dp.ISRmux.d0[14] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net105));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[15]$_DFF_PP0_  (.D(\dp.ISRmux.d0[15] ),
    .RN(_00000_),
    .CLK(clknet_6_40__leaf_clk),
    .Q(net106));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[16]$_DFF_PP0_  (.D(\dp.ISRmux.d0[16] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net107));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[17]$_DFF_PP0_  (.D(\dp.ISRmux.d0[17] ),
    .RN(_00000_),
    .CLK(clknet_6_11__leaf_clk),
    .Q(net108));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[18]$_DFF_PP0_  (.D(\dp.ISRmux.d0[18] ),
    .RN(_00000_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(net109));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[19]$_DFF_PP0_  (.D(\dp.ISRmux.d0[19] ),
    .RN(_00000_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(net110));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[1]$_DFFE_PP0P_  (.D(_00002_),
    .RN(_00000_),
    .CLK(clknet_6_15__leaf_clk),
    .Q(net111));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[20]$_DFF_PP0_  (.D(\dp.ISRmux.d0[20] ),
    .RN(_00000_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(net112));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[21]$_DFF_PP0_  (.D(\dp.ISRmux.d0[21] ),
    .RN(_00000_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(net113));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[22]$_DFF_PP0_  (.D(\dp.ISRmux.d0[22] ),
    .RN(_00000_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(net114));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[23]$_DFF_PP0_  (.D(\dp.ISRmux.d0[23] ),
    .RN(_00000_),
    .CLK(clknet_6_11__leaf_clk),
    .Q(net115));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[24]$_DFF_PP0_  (.D(\dp.ISRmux.d0[24] ),
    .RN(_00000_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(net116));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[25]$_DFF_PP0_  (.D(\dp.ISRmux.d0[25] ),
    .RN(_00000_),
    .CLK(clknet_6_11__leaf_clk),
    .Q(net117));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[26]$_DFF_PP0_  (.D(\dp.ISRmux.d0[26] ),
    .RN(_00000_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(net118));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[27]$_DFF_PP0_  (.D(\dp.ISRmux.d0[27] ),
    .RN(_00000_),
    .CLK(clknet_6_11__leaf_clk),
    .Q(net119));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[28]$_DFF_PP0_  (.D(\dp.ISRmux.d0[28] ),
    .RN(_00000_),
    .CLK(clknet_leaf_20_clk),
    .Q(net120));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[29]$_DFF_PP0_  (.D(\dp.ISRmux.d0[29] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net121));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[2]$_DFF_PP0_  (.D(\dp.ISRmux.d0[2] ),
    .RN(_00000_),
    .CLK(clknet_6_15__leaf_clk),
    .Q(net122));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[30]$_DFF_PP0_  (.D(\dp.ISRmux.d0[30] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net123));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[31]$_DFF_PP0_  (.D(\dp.ISRmux.d0[31] ),
    .RN(_00000_),
    .CLK(clknet_6_15__leaf_clk),
    .Q(net124));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[3]$_DFF_PP0_  (.D(\dp.ISRmux.d0[3] ),
    .RN(_00000_),
    .CLK(clknet_6_15__leaf_clk),
    .Q(net125));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[4]$_DFF_PP0_  (.D(\dp.ISRmux.d0[4] ),
    .RN(_00000_),
    .CLK(clknet_6_15__leaf_clk),
    .Q(net126));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[5]$_DFF_PP0_  (.D(\dp.ISRmux.d0[5] ),
    .RN(_00000_),
    .CLK(clknet_6_15__leaf_clk),
    .Q(net127));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[6]$_DFF_PP0_  (.D(\dp.ISRmux.d0[6] ),
    .RN(_00000_),
    .CLK(clknet_6_15__leaf_clk),
    .Q(net128));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[7]$_DFF_PP0_  (.D(\dp.ISRmux.d0[7] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net129));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[8]$_DFF_PP0_  (.D(\dp.ISRmux.d0[8] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net130));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \dp.pcreg.q[9]$_DFF_PP0_  (.D(\dp.ISRmux.d0[9] ),
    .RN(_00000_),
    .CLK(clknet_6_14__leaf_clk),
    .Q(net131));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][0]$_DFFE_PP_  (.D(\dp.rf.rf[0][0] ),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\dp.rf.rf[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][10]$_DFFE_PP_  (.D(\dp.rf.rf[0][10] ),
    .CLK(clknet_leaf_270_clk),
    .Q(\dp.rf.rf[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][11]$_DFFE_PP_  (.D(\dp.rf.rf[0][11] ),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][12]$_DFFE_PP_  (.D(\dp.rf.rf[0][12] ),
    .CLK(clknet_6_32__leaf_clk),
    .Q(\dp.rf.rf[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][13]$_DFFE_PP_  (.D(\dp.rf.rf[0][13] ),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\dp.rf.rf[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][14]$_DFFE_PP_  (.D(\dp.rf.rf[0][14] ),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\dp.rf.rf[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][15]$_DFFE_PP_  (.D(\dp.rf.rf[0][15] ),
    .CLK(clknet_leaf_261_clk),
    .Q(\dp.rf.rf[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][16]$_DFFE_PP_  (.D(\dp.rf.rf[0][16] ),
    .CLK(clknet_leaf_411_clk),
    .Q(\dp.rf.rf[0][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][17]$_DFFE_PP_  (.D(\dp.rf.rf[0][17] ),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\dp.rf.rf[0][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][18]$_DFFE_PP_  (.D(\dp.rf.rf[0][18] ),
    .CLK(clknet_leaf_107_clk),
    .Q(\dp.rf.rf[0][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][19]$_DFFE_PP_  (.D(\dp.rf.rf[0][19] ),
    .CLK(clknet_leaf_116_clk),
    .Q(\dp.rf.rf[0][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][1]$_DFFE_PP_  (.D(\dp.rf.rf[0][1] ),
    .CLK(clknet_leaf_497_clk),
    .Q(\dp.rf.rf[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][20]$_DFFE_PP_  (.D(\dp.rf.rf[0][20] ),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\dp.rf.rf[0][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][21]$_DFFE_PP_  (.D(\dp.rf.rf[0][21] ),
    .CLK(clknet_leaf_670_clk),
    .Q(\dp.rf.rf[0][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][22]$_DFFE_PP_  (.D(\dp.rf.rf[0][22] ),
    .CLK(clknet_leaf_679_clk),
    .Q(\dp.rf.rf[0][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][23]$_DFFE_PP_  (.D(\dp.rf.rf[0][23] ),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\dp.rf.rf[0][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][24]$_DFFE_PP_  (.D(\dp.rf.rf[0][24] ),
    .CLK(clknet_leaf_647_clk),
    .Q(\dp.rf.rf[0][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][25]$_DFFE_PP_  (.D(\dp.rf.rf[0][25] ),
    .CLK(clknet_leaf_484_clk),
    .Q(\dp.rf.rf[0][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][26]$_DFFE_PP_  (.D(\dp.rf.rf[0][26] ),
    .CLK(clknet_leaf_668_clk),
    .Q(\dp.rf.rf[0][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][27]$_DFFE_PP_  (.D(\dp.rf.rf[0][27] ),
    .CLK(clknet_leaf_492_clk),
    .Q(\dp.rf.rf[0][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][28]$_DFFE_PP_  (.D(\dp.rf.rf[0][28] ),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[0][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][29]$_DFFE_PP_  (.D(\dp.rf.rf[0][29] ),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[0][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][2]$_DFFE_PP_  (.D(\dp.rf.rf[0][2] ),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\dp.rf.rf[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][30]$_DFFE_PP_  (.D(\dp.rf.rf[0][30] ),
    .CLK(clknet_leaf_569_clk),
    .Q(\dp.rf.rf[0][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][31]$_DFFE_PP_  (.D(\dp.rf.rf[0][31] ),
    .CLK(clknet_6_26__leaf_clk),
    .Q(\dp.rf.rf[0][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][3]$_DFFE_PP_  (.D(\dp.rf.rf[0][3] ),
    .CLK(clknet_leaf_173_clk),
    .Q(\dp.rf.rf[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][4]$_DFFE_PP_  (.D(\dp.rf.rf[0][4] ),
    .CLK(clknet_leaf_513_clk),
    .Q(\dp.rf.rf[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][5]$_DFFE_PP_  (.D(\dp.rf.rf[0][5] ),
    .CLK(clknet_leaf_221_clk),
    .Q(\dp.rf.rf[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][6]$_DFFE_PP_  (.D(\dp.rf.rf[0][6] ),
    .CLK(clknet_leaf_423_clk),
    .Q(\dp.rf.rf[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][7]$_DFFE_PP_  (.D(\dp.rf.rf[0][7] ),
    .CLK(clknet_leaf_113_clk),
    .Q(\dp.rf.rf[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][8]$_DFFE_PP_  (.D(\dp.rf.rf[0][8] ),
    .CLK(clknet_leaf_446_clk),
    .Q(\dp.rf.rf[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[0][9]$_DFFE_PP_  (.D(\dp.rf.rf[0][9] ),
    .CLK(clknet_leaf_640_clk),
    .Q(\dp.rf.rf[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][0]$_DFFE_PP_  (.D(_00035_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\dp.rf.rf[10][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][10]$_DFFE_PP_  (.D(_00036_),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[10][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][11]$_DFFE_PP_  (.D(_00037_),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[10][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][12]$_DFFE_PP_  (.D(_00038_),
    .CLK(clknet_leaf_116_clk),
    .Q(\dp.rf.rf[10][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][13]$_DFFE_PP_  (.D(_00039_),
    .CLK(clknet_leaf_223_clk),
    .Q(\dp.rf.rf[10][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][14]$_DFFE_PP_  (.D(_00040_),
    .CLK(clknet_leaf_237_clk),
    .Q(\dp.rf.rf[10][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][15]$_DFFE_PP_  (.D(_00041_),
    .CLK(clknet_leaf_277_clk),
    .Q(\dp.rf.rf[10][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][16]$_DFFE_PP_  (.D(_00042_),
    .CLK(clknet_leaf_419_clk),
    .Q(\dp.rf.rf[10][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][17]$_DFFE_PP_  (.D(_00043_),
    .CLK(clknet_leaf_313_clk),
    .Q(\dp.rf.rf[10][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][18]$_DFFE_PP_  (.D(_00044_),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\dp.rf.rf[10][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][19]$_DFFE_PP_  (.D(_00045_),
    .CLK(clknet_leaf_78_clk),
    .Q(\dp.rf.rf[10][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][1]$_DFFE_PP_  (.D(_00046_),
    .CLK(clknet_leaf_505_clk),
    .Q(\dp.rf.rf[10][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][20]$_DFFE_PP_  (.D(_00047_),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\dp.rf.rf[10][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][21]$_DFFE_PP_  (.D(_00048_),
    .CLK(clknet_leaf_689_clk),
    .Q(\dp.rf.rf[10][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][22]$_DFFE_PP_  (.D(_00049_),
    .CLK(clknet_leaf_682_clk),
    .Q(\dp.rf.rf[10][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][23]$_DFFE_PP_  (.D(_00050_),
    .CLK(clknet_leaf_469_clk),
    .Q(\dp.rf.rf[10][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][24]$_DFFE_PP_  (.D(_00051_),
    .CLK(clknet_leaf_693_clk),
    .Q(\dp.rf.rf[10][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][25]$_DFFE_PP_  (.D(_00052_),
    .CLK(clknet_leaf_491_clk),
    .Q(\dp.rf.rf[10][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][26]$_DFFE_PP_  (.D(_00053_),
    .CLK(clknet_leaf_704_clk),
    .Q(\dp.rf.rf[10][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][27]$_DFFE_PP_  (.D(_00054_),
    .CLK(clknet_6_20__leaf_clk),
    .Q(\dp.rf.rf[10][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][28]$_DFFE_PP_  (.D(_00055_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[10][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][29]$_DFFE_PP_  (.D(_00056_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[10][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][2]$_DFFE_PP_  (.D(_00057_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[10][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][30]$_DFFE_PP_  (.D(_00058_),
    .CLK(clknet_leaf_530_clk),
    .Q(\dp.rf.rf[10][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][31]$_DFFE_PP_  (.D(_00059_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[10][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][3]$_DFFE_PP_  (.D(_00060_),
    .CLK(clknet_6_58__leaf_clk),
    .Q(\dp.rf.rf[10][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][4]$_DFFE_PP_  (.D(_00061_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\dp.rf.rf[10][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][5]$_DFFE_PP_  (.D(_00062_),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\dp.rf.rf[10][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][6]$_DFFE_PP_  (.D(_00063_),
    .CLK(clknet_leaf_421_clk),
    .Q(\dp.rf.rf[10][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][7]$_DFFE_PP_  (.D(_00064_),
    .CLK(clknet_leaf_74_clk),
    .Q(\dp.rf.rf[10][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][8]$_DFFE_PP_  (.D(_00065_),
    .CLK(clknet_leaf_456_clk),
    .Q(\dp.rf.rf[10][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[10][9]$_DFFE_PP_  (.D(_00066_),
    .CLK(clknet_leaf_632_clk),
    .Q(\dp.rf.rf[10][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][0]$_DFFE_PP_  (.D(_00067_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\dp.rf.rf[11][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][10]$_DFFE_PP_  (.D(_00068_),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[11][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][11]$_DFFE_PP_  (.D(_00069_),
    .CLK(clknet_leaf_264_clk),
    .Q(\dp.rf.rf[11][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][12]$_DFFE_PP_  (.D(_00070_),
    .CLK(clknet_leaf_117_clk),
    .Q(\dp.rf.rf[11][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][13]$_DFFE_PP_  (.D(_00071_),
    .CLK(clknet_leaf_223_clk),
    .Q(\dp.rf.rf[11][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][14]$_DFFE_PP_  (.D(_00072_),
    .CLK(clknet_leaf_237_clk),
    .Q(\dp.rf.rf[11][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][15]$_DFFE_PP_  (.D(_00073_),
    .CLK(clknet_leaf_277_clk),
    .Q(\dp.rf.rf[11][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][16]$_DFFE_PP_  (.D(_00074_),
    .CLK(clknet_leaf_419_clk),
    .Q(\dp.rf.rf[11][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][17]$_DFFE_PP_  (.D(_00075_),
    .CLK(clknet_leaf_313_clk),
    .Q(\dp.rf.rf[11][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][18]$_DFFE_PP_  (.D(_00076_),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\dp.rf.rf[11][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][19]$_DFFE_PP_  (.D(_00077_),
    .CLK(clknet_leaf_78_clk),
    .Q(\dp.rf.rf[11][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][1]$_DFFE_PP_  (.D(_00078_),
    .CLK(clknet_leaf_505_clk),
    .Q(\dp.rf.rf[11][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][20]$_DFFE_PP_  (.D(_00079_),
    .CLK(clknet_leaf_459_clk),
    .Q(\dp.rf.rf[11][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][21]$_DFFE_PP_  (.D(_00080_),
    .CLK(clknet_leaf_689_clk),
    .Q(\dp.rf.rf[11][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][22]$_DFFE_PP_  (.D(_00081_),
    .CLK(clknet_leaf_682_clk),
    .Q(\dp.rf.rf[11][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][23]$_DFFE_PP_  (.D(_00082_),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\dp.rf.rf[11][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][24]$_DFFE_PP_  (.D(_00083_),
    .CLK(clknet_leaf_693_clk),
    .Q(\dp.rf.rf[11][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][25]$_DFFE_PP_  (.D(_00084_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[11][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][26]$_DFFE_PP_  (.D(_00085_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[11][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][27]$_DFFE_PP_  (.D(_00086_),
    .CLK(clknet_6_20__leaf_clk),
    .Q(\dp.rf.rf[11][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][28]$_DFFE_PP_  (.D(_00087_),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\dp.rf.rf[11][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][29]$_DFFE_PP_  (.D(_00088_),
    .CLK(clknet_leaf_441_clk),
    .Q(\dp.rf.rf[11][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][2]$_DFFE_PP_  (.D(_00089_),
    .CLK(clknet_leaf_2_clk),
    .Q(\dp.rf.rf[11][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][30]$_DFFE_PP_  (.D(_00090_),
    .CLK(clknet_leaf_530_clk),
    .Q(\dp.rf.rf[11][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][31]$_DFFE_PP_  (.D(_00091_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[11][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][3]$_DFFE_PP_  (.D(_00092_),
    .CLK(clknet_leaf_198_clk),
    .Q(\dp.rf.rf[11][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][4]$_DFFE_PP_  (.D(_00093_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\dp.rf.rf[11][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][5]$_DFFE_PP_  (.D(_00094_),
    .CLK(clknet_leaf_131_clk),
    .Q(\dp.rf.rf[11][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][6]$_DFFE_PP_  (.D(_00095_),
    .CLK(clknet_leaf_421_clk),
    .Q(\dp.rf.rf[11][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][7]$_DFFE_PP_  (.D(_00096_),
    .CLK(clknet_leaf_74_clk),
    .Q(\dp.rf.rf[11][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][8]$_DFFE_PP_  (.D(_00097_),
    .CLK(clknet_leaf_456_clk),
    .Q(\dp.rf.rf[11][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[11][9]$_DFFE_PP_  (.D(_00098_),
    .CLK(clknet_leaf_632_clk),
    .Q(\dp.rf.rf[11][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][0]$_DFFE_PP_  (.D(_00099_),
    .CLK(clknet_leaf_160_clk),
    .Q(\dp.rf.rf[12][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][10]$_DFFE_PP_  (.D(_00100_),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[12][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][11]$_DFFE_PP_  (.D(_00101_),
    .CLK(clknet_leaf_261_clk),
    .Q(\dp.rf.rf[12][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][12]$_DFFE_PP_  (.D(_00102_),
    .CLK(clknet_leaf_116_clk),
    .Q(\dp.rf.rf[12][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][13]$_DFFE_PP_  (.D(_00103_),
    .CLK(clknet_leaf_224_clk),
    .Q(\dp.rf.rf[12][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][14]$_DFFE_PP_  (.D(_00104_),
    .CLK(clknet_leaf_228_clk),
    .Q(\dp.rf.rf[12][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][15]$_DFFE_PP_  (.D(_00105_),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\dp.rf.rf[12][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][16]$_DFFE_PP_  (.D(_00106_),
    .CLK(clknet_leaf_411_clk),
    .Q(\dp.rf.rf[12][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][17]$_DFFE_PP_  (.D(_00107_),
    .CLK(clknet_leaf_294_clk),
    .Q(\dp.rf.rf[12][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][18]$_DFFE_PP_  (.D(_00108_),
    .CLK(clknet_leaf_68_clk),
    .Q(\dp.rf.rf[12][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][19]$_DFFE_PP_  (.D(_00109_),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\dp.rf.rf[12][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][1]$_DFFE_PP_  (.D(_00110_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[12][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][20]$_DFFE_PP_  (.D(_00111_),
    .CLK(clknet_6_21__leaf_clk),
    .Q(\dp.rf.rf[12][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][21]$_DFFE_PP_  (.D(_00112_),
    .CLK(clknet_leaf_702_clk),
    .Q(\dp.rf.rf[12][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][22]$_DFFE_PP_  (.D(_00113_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\dp.rf.rf[12][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][23]$_DFFE_PP_  (.D(_00114_),
    .CLK(clknet_leaf_469_clk),
    .Q(\dp.rf.rf[12][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][24]$_DFFE_PP_  (.D(_00115_),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\dp.rf.rf[12][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][25]$_DFFE_PP_  (.D(_00116_),
    .CLK(clknet_leaf_468_clk),
    .Q(\dp.rf.rf[12][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][26]$_DFFE_PP_  (.D(_00117_),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\dp.rf.rf[12][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][27]$_DFFE_PP_  (.D(_00118_),
    .CLK(clknet_leaf_493_clk),
    .Q(\dp.rf.rf[12][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][28]$_DFFE_PP_  (.D(_00119_),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\dp.rf.rf[12][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][29]$_DFFE_PP_  (.D(_00120_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[12][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][2]$_DFFE_PP_  (.D(_00121_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\dp.rf.rf[12][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][30]$_DFFE_PP_  (.D(_00122_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[12][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][31]$_DFFE_PP_  (.D(_00123_),
    .CLK(clknet_leaf_436_clk),
    .Q(\dp.rf.rf[12][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][3]$_DFFE_PP_  (.D(_00124_),
    .CLK(clknet_leaf_198_clk),
    .Q(\dp.rf.rf[12][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][4]$_DFFE_PP_  (.D(_00125_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\dp.rf.rf[12][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][5]$_DFFE_PP_  (.D(_00126_),
    .CLK(clknet_leaf_127_clk),
    .Q(\dp.rf.rf[12][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][6]$_DFFE_PP_  (.D(_00127_),
    .CLK(clknet_leaf_424_clk),
    .Q(\dp.rf.rf[12][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][7]$_DFFE_PP_  (.D(_00128_),
    .CLK(clknet_leaf_73_clk),
    .Q(\dp.rf.rf[12][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][8]$_DFFE_PP_  (.D(_00129_),
    .CLK(clknet_leaf_458_clk),
    .Q(\dp.rf.rf[12][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[12][9]$_DFFE_PP_  (.D(_00130_),
    .CLK(clknet_leaf_631_clk),
    .Q(\dp.rf.rf[12][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][0]$_DFFE_PP_  (.D(_00131_),
    .CLK(clknet_leaf_161_clk),
    .Q(\dp.rf.rf[13][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][10]$_DFFE_PP_  (.D(_00132_),
    .CLK(clknet_leaf_264_clk),
    .Q(\dp.rf.rf[13][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][11]$_DFFE_PP_  (.D(_00133_),
    .CLK(clknet_leaf_261_clk),
    .Q(\dp.rf.rf[13][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][12]$_DFFE_PP_  (.D(_00134_),
    .CLK(clknet_leaf_125_clk),
    .Q(\dp.rf.rf[13][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][13]$_DFFE_PP_  (.D(_00135_),
    .CLK(clknet_leaf_224_clk),
    .Q(\dp.rf.rf[13][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][14]$_DFFE_PP_  (.D(_00136_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\dp.rf.rf[13][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][15]$_DFFE_PP_  (.D(_00137_),
    .CLK(clknet_leaf_276_clk),
    .Q(\dp.rf.rf[13][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][16]$_DFFE_PP_  (.D(_00138_),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\dp.rf.rf[13][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][17]$_DFFE_PP_  (.D(_00139_),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\dp.rf.rf[13][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][18]$_DFFE_PP_  (.D(_00140_),
    .CLK(clknet_leaf_68_clk),
    .Q(\dp.rf.rf[13][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][19]$_DFFE_PP_  (.D(_00141_),
    .CLK(clknet_leaf_75_clk),
    .Q(\dp.rf.rf[13][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][1]$_DFFE_PP_  (.D(_00142_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[13][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][20]$_DFFE_PP_  (.D(_00143_),
    .CLK(clknet_6_21__leaf_clk),
    .Q(\dp.rf.rf[13][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][21]$_DFFE_PP_  (.D(_00144_),
    .CLK(clknet_leaf_702_clk),
    .Q(\dp.rf.rf[13][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][22]$_DFFE_PP_  (.D(_00145_),
    .CLK(clknet_leaf_684_clk),
    .Q(\dp.rf.rf[13][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][23]$_DFFE_PP_  (.D(_00146_),
    .CLK(clknet_6_21__leaf_clk),
    .Q(\dp.rf.rf[13][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][24]$_DFFE_PP_  (.D(_00147_),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\dp.rf.rf[13][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][25]$_DFFE_PP_  (.D(_00148_),
    .CLK(clknet_leaf_473_clk),
    .Q(\dp.rf.rf[13][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][26]$_DFFE_PP_  (.D(_00149_),
    .CLK(clknet_leaf_704_clk),
    .Q(\dp.rf.rf[13][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][27]$_DFFE_PP_  (.D(_00150_),
    .CLK(clknet_leaf_493_clk),
    .Q(\dp.rf.rf[13][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][28]$_DFFE_PP_  (.D(_00151_),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\dp.rf.rf[13][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][29]$_DFFE_PP_  (.D(_00152_),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\dp.rf.rf[13][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][2]$_DFFE_PP_  (.D(_00153_),
    .CLK(clknet_leaf_22_clk),
    .Q(\dp.rf.rf[13][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][30]$_DFFE_PP_  (.D(_00154_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[13][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][31]$_DFFE_PP_  (.D(_00155_),
    .CLK(clknet_leaf_436_clk),
    .Q(\dp.rf.rf[13][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][3]$_DFFE_PP_  (.D(_00156_),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\dp.rf.rf[13][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][4]$_DFFE_PP_  (.D(_00157_),
    .CLK(clknet_leaf_513_clk),
    .Q(\dp.rf.rf[13][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][5]$_DFFE_PP_  (.D(_00158_),
    .CLK(clknet_leaf_127_clk),
    .Q(\dp.rf.rf[13][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][6]$_DFFE_PP_  (.D(_00159_),
    .CLK(clknet_leaf_423_clk),
    .Q(\dp.rf.rf[13][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][7]$_DFFE_PP_  (.D(_00160_),
    .CLK(clknet_leaf_73_clk),
    .Q(\dp.rf.rf[13][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][8]$_DFFE_PP_  (.D(_00161_),
    .CLK(clknet_leaf_458_clk),
    .Q(\dp.rf.rf[13][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[13][9]$_DFFE_PP_  (.D(_00162_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\dp.rf.rf[13][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][0]$_DFFE_PP_  (.D(_00163_),
    .CLK(clknet_leaf_162_clk),
    .Q(\dp.rf.rf[14][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][10]$_DFFE_PP_  (.D(_00164_),
    .CLK(clknet_leaf_268_clk),
    .Q(\dp.rf.rf[14][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][11]$_DFFE_PP_  (.D(_00165_),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\dp.rf.rf[14][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][12]$_DFFE_PP_  (.D(_00166_),
    .CLK(clknet_leaf_117_clk),
    .Q(\dp.rf.rf[14][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][13]$_DFFE_PP_  (.D(_00167_),
    .CLK(clknet_leaf_222_clk),
    .Q(\dp.rf.rf[14][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][14]$_DFFE_PP_  (.D(_00168_),
    .CLK(clknet_leaf_228_clk),
    .Q(\dp.rf.rf[14][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][15]$_DFFE_PP_  (.D(_00169_),
    .CLK(clknet_leaf_254_clk),
    .Q(\dp.rf.rf[14][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][16]$_DFFE_PP_  (.D(_00170_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[14][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][17]$_DFFE_PP_  (.D(_00171_),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\dp.rf.rf[14][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][18]$_DFFE_PP_  (.D(_00172_),
    .CLK(clknet_leaf_65_clk),
    .Q(\dp.rf.rf[14][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][19]$_DFFE_PP_  (.D(_00173_),
    .CLK(clknet_leaf_75_clk),
    .Q(\dp.rf.rf[14][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][1]$_DFFE_PP_  (.D(_00174_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[14][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][20]$_DFFE_PP_  (.D(_00175_),
    .CLK(clknet_6_21__leaf_clk),
    .Q(\dp.rf.rf[14][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][21]$_DFFE_PP_  (.D(_00176_),
    .CLK(clknet_leaf_700_clk),
    .Q(\dp.rf.rf[14][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][22]$_DFFE_PP_  (.D(_00177_),
    .CLK(clknet_leaf_692_clk),
    .Q(\dp.rf.rf[14][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][23]$_DFFE_PP_  (.D(_00178_),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\dp.rf.rf[14][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][24]$_DFFE_PP_  (.D(_00179_),
    .CLK(clknet_leaf_694_clk),
    .Q(\dp.rf.rf[14][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][25]$_DFFE_PP_  (.D(_00180_),
    .CLK(clknet_leaf_484_clk),
    .Q(\dp.rf.rf[14][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][26]$_DFFE_PP_  (.D(_00181_),
    .CLK(clknet_leaf_705_clk),
    .Q(\dp.rf.rf[14][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][27]$_DFFE_PP_  (.D(_00182_),
    .CLK(clknet_6_20__leaf_clk),
    .Q(\dp.rf.rf[14][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][28]$_DFFE_PP_  (.D(_00183_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[14][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][29]$_DFFE_PP_  (.D(_00184_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[14][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][2]$_DFFE_PP_  (.D(_00185_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\dp.rf.rf[14][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][30]$_DFFE_PP_  (.D(_00186_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[14][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][31]$_DFFE_PP_  (.D(_00187_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[14][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][3]$_DFFE_PP_  (.D(_00188_),
    .CLK(clknet_leaf_200_clk),
    .Q(\dp.rf.rf[14][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][4]$_DFFE_PP_  (.D(_00189_),
    .CLK(clknet_leaf_628_clk),
    .Q(\dp.rf.rf[14][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][5]$_DFFE_PP_  (.D(_00190_),
    .CLK(clknet_leaf_126_clk),
    .Q(\dp.rf.rf[14][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][6]$_DFFE_PP_  (.D(_00191_),
    .CLK(clknet_leaf_425_clk),
    .Q(\dp.rf.rf[14][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][7]$_DFFE_PP_  (.D(_00192_),
    .CLK(clknet_leaf_67_clk),
    .Q(\dp.rf.rf[14][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][8]$_DFFE_PP_  (.D(_00193_),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\dp.rf.rf[14][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[14][9]$_DFFE_PP_  (.D(_00194_),
    .CLK(clknet_leaf_640_clk),
    .Q(\dp.rf.rf[14][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][0]$_DFFE_PP_  (.D(_00195_),
    .CLK(clknet_leaf_162_clk),
    .Q(\dp.rf.rf[15][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][10]$_DFFE_PP_  (.D(_00196_),
    .CLK(clknet_leaf_268_clk),
    .Q(\dp.rf.rf[15][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][11]$_DFFE_PP_  (.D(_00197_),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\dp.rf.rf[15][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][12]$_DFFE_PP_  (.D(_00198_),
    .CLK(clknet_leaf_118_clk),
    .Q(\dp.rf.rf[15][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][13]$_DFFE_PP_  (.D(_00199_),
    .CLK(clknet_leaf_223_clk),
    .Q(\dp.rf.rf[15][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][14]$_DFFE_PP_  (.D(_00200_),
    .CLK(clknet_leaf_230_clk),
    .Q(\dp.rf.rf[15][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][15]$_DFFE_PP_  (.D(_00201_),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\dp.rf.rf[15][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][16]$_DFFE_PP_  (.D(_00202_),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\dp.rf.rf[15][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][17]$_DFFE_PP_  (.D(_00203_),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\dp.rf.rf[15][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][18]$_DFFE_PP_  (.D(_00204_),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\dp.rf.rf[15][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][19]$_DFFE_PP_  (.D(_00205_),
    .CLK(clknet_leaf_76_clk),
    .Q(\dp.rf.rf[15][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][1]$_DFFE_PP_  (.D(_00206_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[15][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][20]$_DFFE_PP_  (.D(_00207_),
    .CLK(clknet_leaf_449_clk),
    .Q(\dp.rf.rf[15][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][21]$_DFFE_PP_  (.D(_00208_),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\dp.rf.rf[15][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][22]$_DFFE_PP_  (.D(_00209_),
    .CLK(clknet_leaf_692_clk),
    .Q(\dp.rf.rf[15][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][23]$_DFFE_PP_  (.D(_00210_),
    .CLK(clknet_leaf_473_clk),
    .Q(\dp.rf.rf[15][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][24]$_DFFE_PP_  (.D(_00211_),
    .CLK(clknet_leaf_694_clk),
    .Q(\dp.rf.rf[15][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][25]$_DFFE_PP_  (.D(_00212_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[15][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][26]$_DFFE_PP_  (.D(_00213_),
    .CLK(clknet_leaf_705_clk),
    .Q(\dp.rf.rf[15][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][27]$_DFFE_PP_  (.D(_00214_),
    .CLK(clknet_leaf_491_clk),
    .Q(\dp.rf.rf[15][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][28]$_DFFE_PP_  (.D(_00215_),
    .CLK(clknet_leaf_0_clk),
    .Q(\dp.rf.rf[15][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][29]$_DFFE_PP_  (.D(_00216_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[15][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][2]$_DFFE_PP_  (.D(_00217_),
    .CLK(clknet_leaf_25_clk),
    .Q(\dp.rf.rf[15][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][30]$_DFFE_PP_  (.D(_00218_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[15][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][31]$_DFFE_PP_  (.D(_00219_),
    .CLK(clknet_leaf_380_clk),
    .Q(\dp.rf.rf[15][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][3]$_DFFE_PP_  (.D(_00220_),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\dp.rf.rf[15][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][4]$_DFFE_PP_  (.D(_00221_),
    .CLK(clknet_leaf_628_clk),
    .Q(\dp.rf.rf[15][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][5]$_DFFE_PP_  (.D(_00222_),
    .CLK(clknet_leaf_126_clk),
    .Q(\dp.rf.rf[15][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][6]$_DFFE_PP_  (.D(_00223_),
    .CLK(clknet_leaf_425_clk),
    .Q(\dp.rf.rf[15][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][7]$_DFFE_PP_  (.D(_00224_),
    .CLK(clknet_leaf_67_clk),
    .Q(\dp.rf.rf[15][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][8]$_DFFE_PP_  (.D(_00225_),
    .CLK(clknet_leaf_452_clk),
    .Q(\dp.rf.rf[15][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[15][9]$_DFFE_PP_  (.D(_00226_),
    .CLK(clknet_leaf_642_clk),
    .Q(\dp.rf.rf[15][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][0]$_DFFE_PP_  (.D(_00227_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[16][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][10]$_DFFE_PP_  (.D(_00228_),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\dp.rf.rf[16][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][11]$_DFFE_PP_  (.D(_00229_),
    .CLK(clknet_leaf_280_clk),
    .Q(\dp.rf.rf[16][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][12]$_DFFE_PP_  (.D(_00230_),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\dp.rf.rf[16][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][13]$_DFFE_PP_  (.D(_00231_),
    .CLK(clknet_leaf_193_clk),
    .Q(\dp.rf.rf[16][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][14]$_DFFE_PP_  (.D(_00232_),
    .CLK(clknet_leaf_250_clk),
    .Q(\dp.rf.rf[16][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][15]$_DFFE_PP_  (.D(_00233_),
    .CLK(clknet_leaf_195_clk),
    .Q(\dp.rf.rf[16][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][16]$_DFFE_PP_  (.D(_00234_),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\dp.rf.rf[16][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][17]$_DFFE_PP_  (.D(_00235_),
    .CLK(clknet_leaf_330_clk),
    .Q(\dp.rf.rf[16][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][18]$_DFFE_PP_  (.D(_00236_),
    .CLK(clknet_leaf_99_clk),
    .Q(\dp.rf.rf[16][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][19]$_DFFE_PP_  (.D(_00237_),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\dp.rf.rf[16][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][1]$_DFFE_PP_  (.D(_00238_),
    .CLK(clknet_leaf_533_clk),
    .Q(\dp.rf.rf[16][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][20]$_DFFE_PP_  (.D(_00239_),
    .CLK(clknet_6_26__leaf_clk),
    .Q(\dp.rf.rf[16][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][21]$_DFFE_PP_  (.D(_00240_),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\dp.rf.rf[16][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][22]$_DFFE_PP_  (.D(_00241_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\dp.rf.rf[16][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][23]$_DFFE_PP_  (.D(_00242_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\dp.rf.rf[16][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][24]$_DFFE_PP_  (.D(_00243_),
    .CLK(clknet_leaf_656_clk),
    .Q(\dp.rf.rf[16][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][25]$_DFFE_PP_  (.D(_00244_),
    .CLK(clknet_leaf_572_clk),
    .Q(\dp.rf.rf[16][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][26]$_DFFE_PP_  (.D(_00245_),
    .CLK(clknet_leaf_592_clk),
    .Q(\dp.rf.rf[16][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][27]$_DFFE_PP_  (.D(_00246_),
    .CLK(clknet_leaf_534_clk),
    .Q(\dp.rf.rf[16][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][28]$_DFFE_PP_  (.D(_00247_),
    .CLK(clknet_leaf_597_clk),
    .Q(\dp.rf.rf[16][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][29]$_DFFE_PP_  (.D(_00248_),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\dp.rf.rf[16][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][2]$_DFFE_PP_  (.D(_00249_),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\dp.rf.rf[16][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][30]$_DFFE_PP_  (.D(_00250_),
    .CLK(clknet_leaf_578_clk),
    .Q(\dp.rf.rf[16][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][31]$_DFFE_PP_  (.D(_00251_),
    .CLK(clknet_leaf_349_clk),
    .Q(\dp.rf.rf[16][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][3]$_DFFE_PP_  (.D(_00252_),
    .CLK(clknet_leaf_173_clk),
    .Q(\dp.rf.rf[16][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][4]$_DFFE_PP_  (.D(_00253_),
    .CLK(clknet_leaf_614_clk),
    .Q(\dp.rf.rf[16][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][5]$_DFFE_PP_  (.D(_00254_),
    .CLK(clknet_leaf_205_clk),
    .Q(\dp.rf.rf[16][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][6]$_DFFE_PP_  (.D(_00255_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\dp.rf.rf[16][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][7]$_DFFE_PP_  (.D(_00256_),
    .CLK(clknet_leaf_98_clk),
    .Q(\dp.rf.rf[16][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][8]$_DFFE_PP_  (.D(_00257_),
    .CLK(clknet_leaf_390_clk),
    .Q(\dp.rf.rf[16][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[16][9]$_DFFE_PP_  (.D(_00258_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\dp.rf.rf[16][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][0]$_DFFE_PP_  (.D(_00259_),
    .CLK(clknet_leaf_328_clk),
    .Q(\dp.rf.rf[17][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][10]$_DFFE_PP_  (.D(_00260_),
    .CLK(clknet_leaf_316_clk),
    .Q(\dp.rf.rf[17][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][11]$_DFFE_PP_  (.D(_00261_),
    .CLK(clknet_leaf_253_clk),
    .Q(\dp.rf.rf[17][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][12]$_DFFE_PP_  (.D(_00262_),
    .CLK(clknet_leaf_143_clk),
    .Q(\dp.rf.rf[17][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][13]$_DFFE_PP_  (.D(_00263_),
    .CLK(clknet_leaf_193_clk),
    .Q(\dp.rf.rf[17][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][14]$_DFFE_PP_  (.D(_00264_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\dp.rf.rf[17][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][15]$_DFFE_PP_  (.D(_00265_),
    .CLK(clknet_leaf_194_clk),
    .Q(\dp.rf.rf[17][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][16]$_DFFE_PP_  (.D(_00266_),
    .CLK(clknet_leaf_334_clk),
    .Q(\dp.rf.rf[17][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][17]$_DFFE_PP_  (.D(_00267_),
    .CLK(clknet_leaf_330_clk),
    .Q(\dp.rf.rf[17][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][18]$_DFFE_PP_  (.D(_00268_),
    .CLK(clknet_leaf_102_clk),
    .Q(\dp.rf.rf[17][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][19]$_DFFE_PP_  (.D(_00269_),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\dp.rf.rf[17][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][1]$_DFFE_PP_  (.D(_00270_),
    .CLK(clknet_leaf_533_clk),
    .Q(\dp.rf.rf[17][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][20]$_DFFE_PP_  (.D(_00271_),
    .CLK(clknet_leaf_366_clk),
    .Q(\dp.rf.rf[17][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][21]$_DFFE_PP_  (.D(_00272_),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\dp.rf.rf[17][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][22]$_DFFE_PP_  (.D(_00273_),
    .CLK(clknet_leaf_655_clk),
    .Q(\dp.rf.rf[17][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][23]$_DFFE_PP_  (.D(_00274_),
    .CLK(clknet_leaf_372_clk),
    .Q(\dp.rf.rf[17][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][24]$_DFFE_PP_  (.D(_00275_),
    .CLK(clknet_leaf_656_clk),
    .Q(\dp.rf.rf[17][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][25]$_DFFE_PP_  (.D(_00276_),
    .CLK(clknet_leaf_572_clk),
    .Q(\dp.rf.rf[17][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][26]$_DFFE_PP_  (.D(_00277_),
    .CLK(clknet_leaf_592_clk),
    .Q(\dp.rf.rf[17][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][27]$_DFFE_PP_  (.D(_00278_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[17][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][28]$_DFFE_PP_  (.D(_00279_),
    .CLK(clknet_leaf_597_clk),
    .Q(\dp.rf.rf[17][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][29]$_DFFE_PP_  (.D(_00280_),
    .CLK(clknet_leaf_561_clk),
    .Q(\dp.rf.rf[17][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][2]$_DFFE_PP_  (.D(_00281_),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\dp.rf.rf[17][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][30]$_DFFE_PP_  (.D(_00282_),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\dp.rf.rf[17][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][31]$_DFFE_PP_  (.D(_00283_),
    .CLK(clknet_leaf_351_clk),
    .Q(\dp.rf.rf[17][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][3]$_DFFE_PP_  (.D(_00284_),
    .CLK(clknet_leaf_174_clk),
    .Q(\dp.rf.rf[17][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][4]$_DFFE_PP_  (.D(_00285_),
    .CLK(clknet_leaf_616_clk),
    .Q(\dp.rf.rf[17][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][5]$_DFFE_PP_  (.D(_00286_),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\dp.rf.rf[17][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][6]$_DFFE_PP_  (.D(_00287_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\dp.rf.rf[17][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][7]$_DFFE_PP_  (.D(_00288_),
    .CLK(clknet_leaf_94_clk),
    .Q(\dp.rf.rf[17][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][8]$_DFFE_PP_  (.D(_00289_),
    .CLK(clknet_leaf_365_clk),
    .Q(\dp.rf.rf[17][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[17][9]$_DFFE_PP_  (.D(_00290_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\dp.rf.rf[17][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][0]$_DFFE_PP_  (.D(_00291_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[18][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][10]$_DFFE_PP_  (.D(_00292_),
    .CLK(clknet_leaf_319_clk),
    .Q(\dp.rf.rf[18][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][11]$_DFFE_PP_  (.D(_00293_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\dp.rf.rf[18][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][12]$_DFFE_PP_  (.D(_00294_),
    .CLK(clknet_6_32__leaf_clk),
    .Q(\dp.rf.rf[18][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][13]$_DFFE_PP_  (.D(_00295_),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\dp.rf.rf[18][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][14]$_DFFE_PP_  (.D(_00296_),
    .CLK(clknet_leaf_246_clk),
    .Q(\dp.rf.rf[18][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][15]$_DFFE_PP_  (.D(_00297_),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\dp.rf.rf[18][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][16]$_DFFE_PP_  (.D(_00298_),
    .CLK(clknet_leaf_333_clk),
    .Q(\dp.rf.rf[18][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][17]$_DFFE_PP_  (.D(_00299_),
    .CLK(clknet_leaf_328_clk),
    .Q(\dp.rf.rf[18][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][18]$_DFFE_PP_  (.D(_00300_),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\dp.rf.rf[18][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][19]$_DFFE_PP_  (.D(_00301_),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\dp.rf.rf[18][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][1]$_DFFE_PP_  (.D(_00302_),
    .CLK(clknet_leaf_614_clk),
    .Q(\dp.rf.rf[18][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][20]$_DFFE_PP_  (.D(_00303_),
    .CLK(clknet_6_26__leaf_clk),
    .Q(\dp.rf.rf[18][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][21]$_DFFE_PP_  (.D(_00304_),
    .CLK(clknet_leaf_596_clk),
    .Q(\dp.rf.rf[18][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][22]$_DFFE_PP_  (.D(_00305_),
    .CLK(clknet_leaf_598_clk),
    .Q(\dp.rf.rf[18][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][23]$_DFFE_PP_  (.D(_00306_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\dp.rf.rf[18][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][24]$_DFFE_PP_  (.D(_00307_),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\dp.rf.rf[18][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][25]$_DFFE_PP_  (.D(_00308_),
    .CLK(clknet_leaf_570_clk),
    .Q(\dp.rf.rf[18][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][26]$_DFFE_PP_  (.D(_00309_),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\dp.rf.rf[18][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][27]$_DFFE_PP_  (.D(_00310_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[18][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][28]$_DFFE_PP_  (.D(_00311_),
    .CLK(clknet_leaf_598_clk),
    .Q(\dp.rf.rf[18][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][29]$_DFFE_PP_  (.D(_00312_),
    .CLK(clknet_leaf_569_clk),
    .Q(\dp.rf.rf[18][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][2]$_DFFE_PP_  (.D(_00313_),
    .CLK(clknet_leaf_591_clk),
    .Q(\dp.rf.rf[18][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][30]$_DFFE_PP_  (.D(_00314_),
    .CLK(clknet_leaf_588_clk),
    .Q(\dp.rf.rf[18][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][31]$_DFFE_PP_  (.D(_00315_),
    .CLK(clknet_leaf_351_clk),
    .Q(\dp.rf.rf[18][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][3]$_DFFE_PP_  (.D(_00316_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\dp.rf.rf[18][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][4]$_DFFE_PP_  (.D(_00317_),
    .CLK(clknet_leaf_614_clk),
    .Q(\dp.rf.rf[18][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][5]$_DFFE_PP_  (.D(_00318_),
    .CLK(clknet_leaf_136_clk),
    .Q(\dp.rf.rf[18][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][6]$_DFFE_PP_  (.D(_00319_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\dp.rf.rf[18][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][7]$_DFFE_PP_  (.D(_00320_),
    .CLK(clknet_leaf_94_clk),
    .Q(\dp.rf.rf[18][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][8]$_DFFE_PP_  (.D(_00321_),
    .CLK(clknet_leaf_365_clk),
    .Q(\dp.rf.rf[18][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[18][9]$_DFFE_PP_  (.D(_00322_),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\dp.rf.rf[18][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][0]$_DFFE_PP_  (.D(_00323_),
    .CLK(clknet_leaf_326_clk),
    .Q(\dp.rf.rf[19][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][10]$_DFFE_PP_  (.D(_00324_),
    .CLK(clknet_leaf_319_clk),
    .Q(\dp.rf.rf[19][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][11]$_DFFE_PP_  (.D(_00325_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\dp.rf.rf[19][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][12]$_DFFE_PP_  (.D(_00326_),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\dp.rf.rf[19][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][13]$_DFFE_PP_  (.D(_00327_),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\dp.rf.rf[19][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][14]$_DFFE_PP_  (.D(_00328_),
    .CLK(clknet_leaf_248_clk),
    .Q(\dp.rf.rf[19][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][15]$_DFFE_PP_  (.D(_00329_),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\dp.rf.rf[19][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][16]$_DFFE_PP_  (.D(_00330_),
    .CLK(clknet_leaf_333_clk),
    .Q(\dp.rf.rf[19][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][17]$_DFFE_PP_  (.D(_00331_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[19][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][18]$_DFFE_PP_  (.D(_00332_),
    .CLK(clknet_leaf_99_clk),
    .Q(\dp.rf.rf[19][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][19]$_DFFE_PP_  (.D(_00333_),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\dp.rf.rf[19][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][1]$_DFFE_PP_  (.D(_00334_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\dp.rf.rf[19][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][20]$_DFFE_PP_  (.D(_00335_),
    .CLK(clknet_leaf_358_clk),
    .Q(\dp.rf.rf[19][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][21]$_DFFE_PP_  (.D(_00336_),
    .CLK(clknet_leaf_596_clk),
    .Q(\dp.rf.rf[19][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][22]$_DFFE_PP_  (.D(_00337_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\dp.rf.rf[19][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][23]$_DFFE_PP_  (.D(_00338_),
    .CLK(clknet_6_26__leaf_clk),
    .Q(\dp.rf.rf[19][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][24]$_DFFE_PP_  (.D(_00339_),
    .CLK(clknet_leaf_596_clk),
    .Q(\dp.rf.rf[19][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][25]$_DFFE_PP_  (.D(_00340_),
    .CLK(clknet_leaf_570_clk),
    .Q(\dp.rf.rf[19][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][26]$_DFFE_PP_  (.D(_00341_),
    .CLK(clknet_leaf_595_clk),
    .Q(\dp.rf.rf[19][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][27]$_DFFE_PP_  (.D(_00342_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[19][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][28]$_DFFE_PP_  (.D(_00343_),
    .CLK(clknet_leaf_598_clk),
    .Q(\dp.rf.rf[19][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][29]$_DFFE_PP_  (.D(_00344_),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\dp.rf.rf[19][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][2]$_DFFE_PP_  (.D(_00345_),
    .CLK(clknet_leaf_591_clk),
    .Q(\dp.rf.rf[19][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][30]$_DFFE_PP_  (.D(_00346_),
    .CLK(clknet_6_15__leaf_clk),
    .Q(\dp.rf.rf[19][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][31]$_DFFE_PP_  (.D(_00347_),
    .CLK(clknet_leaf_349_clk),
    .Q(\dp.rf.rf[19][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][3]$_DFFE_PP_  (.D(_00348_),
    .CLK(clknet_leaf_161_clk),
    .Q(\dp.rf.rf[19][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][4]$_DFFE_PP_  (.D(_00349_),
    .CLK(clknet_leaf_616_clk),
    .Q(\dp.rf.rf[19][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][5]$_DFFE_PP_  (.D(_00350_),
    .CLK(clknet_leaf_141_clk),
    .Q(\dp.rf.rf[19][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][6]$_DFFE_PP_  (.D(_00351_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\dp.rf.rf[19][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][7]$_DFFE_PP_  (.D(_00352_),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\dp.rf.rf[19][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][8]$_DFFE_PP_  (.D(_00353_),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\dp.rf.rf[19][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[19][9]$_DFFE_PP_  (.D(_00354_),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\dp.rf.rf[19][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][0]$_DFFE_PP_  (.D(_00355_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][10]$_DFFE_PP_  (.D(_00356_),
    .CLK(clknet_leaf_270_clk),
    .Q(\dp.rf.rf[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][11]$_DFFE_PP_  (.D(_00357_),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][12]$_DFFE_PP_  (.D(_00358_),
    .CLK(clknet_leaf_205_clk),
    .Q(\dp.rf.rf[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][13]$_DFFE_PP_  (.D(_00359_),
    .CLK(clknet_leaf_231_clk),
    .Q(\dp.rf.rf[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][14]$_DFFE_PP_  (.D(_00360_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\dp.rf.rf[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][15]$_DFFE_PP_  (.D(_00361_),
    .CLK(clknet_leaf_254_clk),
    .Q(\dp.rf.rf[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][16]$_DFFE_PP_  (.D(_00362_),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\dp.rf.rf[1][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][17]$_DFFE_PP_  (.D(_00363_),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\dp.rf.rf[1][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][18]$_DFFE_PP_  (.D(_00364_),
    .CLK(clknet_leaf_107_clk),
    .Q(\dp.rf.rf[1][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][19]$_DFFE_PP_  (.D(_00365_),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\dp.rf.rf[1][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][1]$_DFFE_PP_  (.D(_00366_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][20]$_DFFE_PP_  (.D(_00367_),
    .CLK(clknet_leaf_452_clk),
    .Q(\dp.rf.rf[1][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][21]$_DFFE_PP_  (.D(_00368_),
    .CLK(clknet_leaf_670_clk),
    .Q(\dp.rf.rf[1][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][22]$_DFFE_PP_  (.D(_00369_),
    .CLK(clknet_leaf_675_clk),
    .Q(\dp.rf.rf[1][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][23]$_DFFE_PP_  (.D(_00370_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[1][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][24]$_DFFE_PP_  (.D(_00371_),
    .CLK(clknet_leaf_647_clk),
    .Q(\dp.rf.rf[1][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][25]$_DFFE_PP_  (.D(_00372_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[1][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][26]$_DFFE_PP_  (.D(_00373_),
    .CLK(clknet_leaf_665_clk),
    .Q(\dp.rf.rf[1][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][27]$_DFFE_PP_  (.D(_00374_),
    .CLK(clknet_leaf_492_clk),
    .Q(\dp.rf.rf[1][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][28]$_DFFE_PP_  (.D(_00375_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[1][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][29]$_DFFE_PP_  (.D(_00376_),
    .CLK(clknet_leaf_545_clk),
    .Q(\dp.rf.rf[1][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][2]$_DFFE_PP_  (.D(_00377_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][30]$_DFFE_PP_  (.D(_00378_),
    .CLK(clknet_leaf_581_clk),
    .Q(\dp.rf.rf[1][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][31]$_DFFE_PP_  (.D(_00379_),
    .CLK(clknet_leaf_374_clk),
    .Q(\dp.rf.rf[1][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][3]$_DFFE_PP_  (.D(_00380_),
    .CLK(clknet_6_58__leaf_clk),
    .Q(\dp.rf.rf[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][4]$_DFFE_PP_  (.D(_00381_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\dp.rf.rf[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][5]$_DFFE_PP_  (.D(_00382_),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\dp.rf.rf[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][6]$_DFFE_PP_  (.D(_00383_),
    .CLK(clknet_leaf_424_clk),
    .Q(\dp.rf.rf[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][7]$_DFFE_PP_  (.D(_00384_),
    .CLK(clknet_leaf_113_clk),
    .Q(\dp.rf.rf[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][8]$_DFFE_PP_  (.D(_00385_),
    .CLK(clknet_leaf_454_clk),
    .Q(\dp.rf.rf[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[1][9]$_DFFE_PP_  (.D(_00386_),
    .CLK(clknet_leaf_639_clk),
    .Q(\dp.rf.rf[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][0]$_DFFE_PP_  (.D(_00387_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[20][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][10]$_DFFE_PP_  (.D(_00388_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\dp.rf.rf[20][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][11]$_DFFE_PP_  (.D(_00389_),
    .CLK(clknet_6_59__leaf_clk),
    .Q(\dp.rf.rf[20][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][12]$_DFFE_PP_  (.D(_00390_),
    .CLK(clknet_leaf_141_clk),
    .Q(\dp.rf.rf[20][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][13]$_DFFE_PP_  (.D(_00391_),
    .CLK(clknet_leaf_192_clk),
    .Q(\dp.rf.rf[20][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][14]$_DFFE_PP_  (.D(_00392_),
    .CLK(clknet_leaf_192_clk),
    .Q(\dp.rf.rf[20][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][15]$_DFFE_PP_  (.D(_00393_),
    .CLK(clknet_leaf_189_clk),
    .Q(\dp.rf.rf[20][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][16]$_DFFE_PP_  (.D(_00394_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[20][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][17]$_DFFE_PP_  (.D(_00395_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[20][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][18]$_DFFE_PP_  (.D(_00396_),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\dp.rf.rf[20][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][19]$_DFFE_PP_  (.D(_00397_),
    .CLK(clknet_leaf_96_clk),
    .Q(\dp.rf.rf[20][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][1]$_DFFE_PP_  (.D(_00398_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[20][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][20]$_DFFE_PP_  (.D(_00399_),
    .CLK(clknet_leaf_366_clk),
    .Q(\dp.rf.rf[20][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][21]$_DFFE_PP_  (.D(_00400_),
    .CLK(clknet_leaf_658_clk),
    .Q(\dp.rf.rf[20][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][22]$_DFFE_PP_  (.D(_00401_),
    .CLK(clknet_leaf_654_clk),
    .Q(\dp.rf.rf[20][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][23]$_DFFE_PP_  (.D(_00402_),
    .CLK(clknet_leaf_370_clk),
    .Q(\dp.rf.rf[20][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][24]$_DFFE_PP_  (.D(_00403_),
    .CLK(clknet_leaf_651_clk),
    .Q(\dp.rf.rf[20][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][25]$_DFFE_PP_  (.D(_00404_),
    .CLK(clknet_leaf_557_clk),
    .Q(\dp.rf.rf[20][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][26]$_DFFE_PP_  (.D(_00405_),
    .CLK(clknet_leaf_42_clk),
    .Q(\dp.rf.rf[20][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][27]$_DFFE_PP_  (.D(_00406_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[20][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][28]$_DFFE_PP_  (.D(_00407_),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\dp.rf.rf[20][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][29]$_DFFE_PP_  (.D(_00408_),
    .CLK(clknet_leaf_561_clk),
    .Q(\dp.rf.rf[20][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][2]$_DFFE_PP_  (.D(_00409_),
    .CLK(clknet_leaf_587_clk),
    .Q(\dp.rf.rf[20][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][30]$_DFFE_PP_  (.D(_00410_),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\dp.rf.rf[20][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][31]$_DFFE_PP_  (.D(_00411_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[20][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][3]$_DFFE_PP_  (.D(_00412_),
    .CLK(clknet_leaf_177_clk),
    .Q(\dp.rf.rf[20][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][4]$_DFFE_PP_  (.D(_00413_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\dp.rf.rf[20][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][5]$_DFFE_PP_  (.D(_00414_),
    .CLK(clknet_leaf_143_clk),
    .Q(\dp.rf.rf[20][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][6]$_DFFE_PP_  (.D(_00415_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[20][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][7]$_DFFE_PP_  (.D(_00416_),
    .CLK(clknet_leaf_95_clk),
    .Q(\dp.rf.rf[20][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][8]$_DFFE_PP_  (.D(_00417_),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\dp.rf.rf[20][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[20][9]$_DFFE_PP_  (.D(_00418_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\dp.rf.rf[20][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][0]$_DFFE_PP_  (.D(_00419_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[21][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][10]$_DFFE_PP_  (.D(_00420_),
    .CLK(clknet_leaf_317_clk),
    .Q(\dp.rf.rf[21][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][11]$_DFFE_PP_  (.D(_00421_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\dp.rf.rf[21][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][12]$_DFFE_PP_  (.D(_00422_),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\dp.rf.rf[21][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][13]$_DFFE_PP_  (.D(_00423_),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\dp.rf.rf[21][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][14]$_DFFE_PP_  (.D(_00424_),
    .CLK(clknet_leaf_211_clk),
    .Q(\dp.rf.rf[21][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][15]$_DFFE_PP_  (.D(_00425_),
    .CLK(clknet_leaf_194_clk),
    .Q(\dp.rf.rf[21][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][16]$_DFFE_PP_  (.D(_00426_),
    .CLK(clknet_leaf_334_clk),
    .Q(\dp.rf.rf[21][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][17]$_DFFE_PP_  (.D(_00427_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[21][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][18]$_DFFE_PP_  (.D(_00428_),
    .CLK(clknet_leaf_98_clk),
    .Q(\dp.rf.rf[21][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][19]$_DFFE_PP_  (.D(_00429_),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\dp.rf.rf[21][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][1]$_DFFE_PP_  (.D(_00430_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[21][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][20]$_DFFE_PP_  (.D(_00431_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\dp.rf.rf[21][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][21]$_DFFE_PP_  (.D(_00432_),
    .CLK(clknet_leaf_651_clk),
    .Q(\dp.rf.rf[21][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][22]$_DFFE_PP_  (.D(_00433_),
    .CLK(clknet_leaf_655_clk),
    .Q(\dp.rf.rf[21][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][23]$_DFFE_PP_  (.D(_00434_),
    .CLK(clknet_leaf_372_clk),
    .Q(\dp.rf.rf[21][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][24]$_DFFE_PP_  (.D(_00435_),
    .CLK(clknet_leaf_658_clk),
    .Q(\dp.rf.rf[21][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][25]$_DFFE_PP_  (.D(_00436_),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\dp.rf.rf[21][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][26]$_DFFE_PP_  (.D(_00437_),
    .CLK(clknet_leaf_42_clk),
    .Q(\dp.rf.rf[21][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][27]$_DFFE_PP_  (.D(_00438_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[21][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][28]$_DFFE_PP_  (.D(_00439_),
    .CLK(clknet_leaf_595_clk),
    .Q(\dp.rf.rf[21][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][29]$_DFFE_PP_  (.D(_00440_),
    .CLK(clknet_leaf_561_clk),
    .Q(\dp.rf.rf[21][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][2]$_DFFE_PP_  (.D(_00441_),
    .CLK(clknet_leaf_587_clk),
    .Q(\dp.rf.rf[21][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][30]$_DFFE_PP_  (.D(_00442_),
    .CLK(clknet_leaf_588_clk),
    .Q(\dp.rf.rf[21][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][31]$_DFFE_PP_  (.D(_00443_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[21][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][3]$_DFFE_PP_  (.D(_00444_),
    .CLK(clknet_leaf_174_clk),
    .Q(\dp.rf.rf[21][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][4]$_DFFE_PP_  (.D(_00445_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\dp.rf.rf[21][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][5]$_DFFE_PP_  (.D(_00446_),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\dp.rf.rf[21][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][6]$_DFFE_PP_  (.D(_00447_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[21][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][7]$_DFFE_PP_  (.D(_00448_),
    .CLK(clknet_leaf_95_clk),
    .Q(\dp.rf.rf[21][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][8]$_DFFE_PP_  (.D(_00449_),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\dp.rf.rf[21][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[21][9]$_DFFE_PP_  (.D(_00450_),
    .CLK(clknet_leaf_618_clk),
    .Q(\dp.rf.rf[21][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][0]$_DFFE_PP_  (.D(_00451_),
    .CLK(clknet_leaf_175_clk),
    .Q(\dp.rf.rf[22][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][10]$_DFFE_PP_  (.D(_00452_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\dp.rf.rf[22][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][11]$_DFFE_PP_  (.D(_00453_),
    .CLK(clknet_leaf_185_clk),
    .Q(\dp.rf.rf[22][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][12]$_DFFE_PP_  (.D(_00454_),
    .CLK(clknet_leaf_150_clk),
    .Q(\dp.rf.rf[22][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][13]$_DFFE_PP_  (.D(_00455_),
    .CLK(clknet_leaf_208_clk),
    .Q(\dp.rf.rf[22][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][14]$_DFFE_PP_  (.D(_00456_),
    .CLK(clknet_leaf_246_clk),
    .Q(\dp.rf.rf[22][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][15]$_DFFE_PP_  (.D(_00457_),
    .CLK(clknet_leaf_195_clk),
    .Q(\dp.rf.rf[22][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][16]$_DFFE_PP_  (.D(_00458_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[22][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][17]$_DFFE_PP_  (.D(_00459_),
    .CLK(clknet_leaf_326_clk),
    .Q(\dp.rf.rf[22][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][18]$_DFFE_PP_  (.D(_00460_),
    .CLK(clknet_leaf_92_clk),
    .Q(\dp.rf.rf[22][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][19]$_DFFE_PP_  (.D(_00461_),
    .CLK(clknet_leaf_84_clk),
    .Q(\dp.rf.rf[22][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][1]$_DFFE_PP_  (.D(_00462_),
    .CLK(clknet_leaf_526_clk),
    .Q(\dp.rf.rf[22][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][20]$_DFFE_PP_  (.D(_00463_),
    .CLK(clknet_leaf_360_clk),
    .Q(\dp.rf.rf[22][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][21]$_DFFE_PP_  (.D(_00464_),
    .CLK(clknet_leaf_665_clk),
    .Q(\dp.rf.rf[22][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][22]$_DFFE_PP_  (.D(_00465_),
    .CLK(clknet_leaf_657_clk),
    .Q(\dp.rf.rf[22][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][23]$_DFFE_PP_  (.D(_00466_),
    .CLK(clknet_leaf_369_clk),
    .Q(\dp.rf.rf[22][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][24]$_DFFE_PP_  (.D(_00467_),
    .CLK(clknet_leaf_673_clk),
    .Q(\dp.rf.rf[22][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][25]$_DFFE_PP_  (.D(_00468_),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\dp.rf.rf[22][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][26]$_DFFE_PP_  (.D(_00469_),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\dp.rf.rf[22][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][27]$_DFFE_PP_  (.D(_00470_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[22][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][28]$_DFFE_PP_  (.D(_00471_),
    .CLK(clknet_leaf_662_clk),
    .Q(\dp.rf.rf[22][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][29]$_DFFE_PP_  (.D(_00472_),
    .CLK(clknet_leaf_562_clk),
    .Q(\dp.rf.rf[22][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][2]$_DFFE_PP_  (.D(_00473_),
    .CLK(clknet_leaf_590_clk),
    .Q(\dp.rf.rf[22][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][30]$_DFFE_PP_  (.D(_00474_),
    .CLK(clknet_leaf_584_clk),
    .Q(\dp.rf.rf[22][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][31]$_DFFE_PP_  (.D(_00475_),
    .CLK(clknet_leaf_348_clk),
    .Q(\dp.rf.rf[22][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][3]$_DFFE_PP_  (.D(_00476_),
    .CLK(clknet_leaf_172_clk),
    .Q(\dp.rf.rf[22][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][4]$_DFFE_PP_  (.D(_00477_),
    .CLK(clknet_leaf_528_clk),
    .Q(\dp.rf.rf[22][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][5]$_DFFE_PP_  (.D(_00478_),
    .CLK(clknet_leaf_141_clk),
    .Q(\dp.rf.rf[22][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][6]$_DFFE_PP_  (.D(_00479_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[22][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][7]$_DFFE_PP_  (.D(_00480_),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\dp.rf.rf[22][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][8]$_DFFE_PP_  (.D(_00481_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[22][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[22][9]$_DFFE_PP_  (.D(_00482_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\dp.rf.rf[22][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][0]$_DFFE_PP_  (.D(_00483_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[23][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][10]$_DFFE_PP_  (.D(_00484_),
    .CLK(clknet_leaf_317_clk),
    .Q(\dp.rf.rf[23][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][11]$_DFFE_PP_  (.D(_00485_),
    .CLK(clknet_leaf_185_clk),
    .Q(\dp.rf.rf[23][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][12]$_DFFE_PP_  (.D(_00486_),
    .CLK(clknet_leaf_150_clk),
    .Q(\dp.rf.rf[23][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][13]$_DFFE_PP_  (.D(_00487_),
    .CLK(clknet_leaf_208_clk),
    .Q(\dp.rf.rf[23][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][14]$_DFFE_PP_  (.D(_00488_),
    .CLK(clknet_leaf_192_clk),
    .Q(\dp.rf.rf[23][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][15]$_DFFE_PP_  (.D(_00489_),
    .CLK(clknet_6_59__leaf_clk),
    .Q(\dp.rf.rf[23][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][16]$_DFFE_PP_  (.D(_00490_),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\dp.rf.rf[23][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][17]$_DFFE_PP_  (.D(_00491_),
    .CLK(clknet_leaf_326_clk),
    .Q(\dp.rf.rf[23][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][18]$_DFFE_PP_  (.D(_00492_),
    .CLK(clknet_leaf_96_clk),
    .Q(\dp.rf.rf[23][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][19]$_DFFE_PP_  (.D(_00493_),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\dp.rf.rf[23][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][1]$_DFFE_PP_  (.D(_00494_),
    .CLK(clknet_leaf_526_clk),
    .Q(\dp.rf.rf[23][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][20]$_DFFE_PP_  (.D(_00495_),
    .CLK(clknet_leaf_360_clk),
    .Q(\dp.rf.rf[23][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][21]$_DFFE_PP_  (.D(_00496_),
    .CLK(clknet_leaf_665_clk),
    .Q(\dp.rf.rf[23][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][22]$_DFFE_PP_  (.D(_00497_),
    .CLK(clknet_leaf_657_clk),
    .Q(\dp.rf.rf[23][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][23]$_DFFE_PP_  (.D(_00498_),
    .CLK(clknet_leaf_369_clk),
    .Q(\dp.rf.rf[23][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][24]$_DFFE_PP_  (.D(_00499_),
    .CLK(clknet_leaf_673_clk),
    .Q(\dp.rf.rf[23][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][25]$_DFFE_PP_  (.D(_00500_),
    .CLK(clknet_leaf_557_clk),
    .Q(\dp.rf.rf[23][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][26]$_DFFE_PP_  (.D(_00501_),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\dp.rf.rf[23][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][27]$_DFFE_PP_  (.D(_00502_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[23][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][28]$_DFFE_PP_  (.D(_00503_),
    .CLK(clknet_leaf_662_clk),
    .Q(\dp.rf.rf[23][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][29]$_DFFE_PP_  (.D(_00504_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[23][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][2]$_DFFE_PP_  (.D(_00505_),
    .CLK(clknet_leaf_590_clk),
    .Q(\dp.rf.rf[23][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][30]$_DFFE_PP_  (.D(_00506_),
    .CLK(clknet_leaf_584_clk),
    .Q(\dp.rf.rf[23][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][31]$_DFFE_PP_  (.D(_00507_),
    .CLK(clknet_leaf_348_clk),
    .Q(\dp.rf.rf[23][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][3]$_DFFE_PP_  (.D(_00508_),
    .CLK(clknet_leaf_172_clk),
    .Q(\dp.rf.rf[23][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][4]$_DFFE_PP_  (.D(_00509_),
    .CLK(clknet_leaf_528_clk),
    .Q(\dp.rf.rf[23][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][5]$_DFFE_PP_  (.D(_00510_),
    .CLK(clknet_leaf_139_clk),
    .Q(\dp.rf.rf[23][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][6]$_DFFE_PP_  (.D(_00511_),
    .CLK(clknet_leaf_358_clk),
    .Q(\dp.rf.rf[23][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][7]$_DFFE_PP_  (.D(_00512_),
    .CLK(clknet_leaf_92_clk),
    .Q(\dp.rf.rf[23][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][8]$_DFFE_PP_  (.D(_00513_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[23][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[23][9]$_DFFE_PP_  (.D(_00514_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\dp.rf.rf[23][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][0]$_DFFE_PP_  (.D(_00515_),
    .CLK(clknet_leaf_319_clk),
    .Q(\dp.rf.rf[24][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][10]$_DFFE_PP_  (.D(_00516_),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\dp.rf.rf[24][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][11]$_DFFE_PP_  (.D(_00517_),
    .CLK(clknet_leaf_283_clk),
    .Q(\dp.rf.rf[24][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][12]$_DFFE_PP_  (.D(_00518_),
    .CLK(clknet_leaf_139_clk),
    .Q(\dp.rf.rf[24][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][13]$_DFFE_PP_  (.D(_00519_),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\dp.rf.rf[24][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][14]$_DFFE_PP_  (.D(_00520_),
    .CLK(clknet_leaf_242_clk),
    .Q(\dp.rf.rf[24][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][15]$_DFFE_PP_  (.D(_00521_),
    .CLK(clknet_6_59__leaf_clk),
    .Q(\dp.rf.rf[24][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][16]$_DFFE_PP_  (.D(_00522_),
    .CLK(clknet_leaf_291_clk),
    .Q(\dp.rf.rf[24][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][17]$_DFFE_PP_  (.D(_00523_),
    .CLK(clknet_leaf_309_clk),
    .Q(\dp.rf.rf[24][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][18]$_DFFE_PP_  (.D(_00524_),
    .CLK(clknet_leaf_58_clk),
    .Q(\dp.rf.rf[24][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][19]$_DFFE_PP_  (.D(_00525_),
    .CLK(clknet_leaf_84_clk),
    .Q(\dp.rf.rf[24][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][1]$_DFFE_PP_  (.D(_00526_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[24][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][20]$_DFFE_PP_  (.D(_00527_),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\dp.rf.rf[24][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][21]$_DFFE_PP_  (.D(_00528_),
    .CLK(clknet_leaf_700_clk),
    .Q(\dp.rf.rf[24][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][22]$_DFFE_PP_  (.D(_00529_),
    .CLK(clknet_leaf_649_clk),
    .Q(\dp.rf.rf[24][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][23]$_DFFE_PP_  (.D(_00530_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[24][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][24]$_DFFE_PP_  (.D(_00531_),
    .CLK(clknet_leaf_638_clk),
    .Q(\dp.rf.rf[24][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][25]$_DFFE_PP_  (.D(_00532_),
    .CLK(clknet_leaf_396_clk),
    .Q(\dp.rf.rf[24][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][26]$_DFFE_PP_  (.D(_00533_),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\dp.rf.rf[24][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][27]$_DFFE_PP_  (.D(_00534_),
    .CLK(clknet_leaf_488_clk),
    .Q(\dp.rf.rf[24][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][28]$_DFFE_PP_  (.D(_00535_),
    .CLK(clknet_leaf_664_clk),
    .Q(\dp.rf.rf[24][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][29]$_DFFE_PP_  (.D(_00536_),
    .CLK(clknet_leaf_438_clk),
    .Q(\dp.rf.rf[24][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][2]$_DFFE_PP_  (.D(_00537_),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\dp.rf.rf[24][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][30]$_DFFE_PP_  (.D(_00538_),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\dp.rf.rf[24][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][31]$_DFFE_PP_  (.D(_00539_),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\dp.rf.rf[24][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][3]$_DFFE_PP_  (.D(_00540_),
    .CLK(clknet_leaf_179_clk),
    .Q(\dp.rf.rf[24][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][4]$_DFFE_PP_  (.D(_00541_),
    .CLK(clknet_leaf_623_clk),
    .Q(\dp.rf.rf[24][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][5]$_DFFE_PP_  (.D(_00542_),
    .CLK(clknet_leaf_216_clk),
    .Q(\dp.rf.rf[24][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][6]$_DFFE_PP_  (.D(_00543_),
    .CLK(clknet_leaf_408_clk),
    .Q(\dp.rf.rf[24][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][7]$_DFFE_PP_  (.D(_00544_),
    .CLK(clknet_leaf_56_clk),
    .Q(\dp.rf.rf[24][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][8]$_DFFE_PP_  (.D(_00545_),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\dp.rf.rf[24][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[24][9]$_DFFE_PP_  (.D(_00546_),
    .CLK(clknet_leaf_622_clk),
    .Q(\dp.rf.rf[24][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][0]$_DFFE_PP_  (.D(_00547_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[25][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][10]$_DFFE_PP_  (.D(_00548_),
    .CLK(clknet_leaf_284_clk),
    .Q(\dp.rf.rf[25][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][11]$_DFFE_PP_  (.D(_00549_),
    .CLK(clknet_leaf_283_clk),
    .Q(\dp.rf.rf[25][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][12]$_DFFE_PP_  (.D(_00550_),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\dp.rf.rf[25][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][13]$_DFFE_PP_  (.D(_00551_),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\dp.rf.rf[25][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][14]$_DFFE_PP_  (.D(_00552_),
    .CLK(clknet_6_62__leaf_clk),
    .Q(\dp.rf.rf[25][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][15]$_DFFE_PP_  (.D(_00553_),
    .CLK(clknet_leaf_187_clk),
    .Q(\dp.rf.rf[25][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][16]$_DFFE_PP_  (.D(_00554_),
    .CLK(clknet_leaf_291_clk),
    .Q(\dp.rf.rf[25][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][17]$_DFFE_PP_  (.D(_00555_),
    .CLK(clknet_leaf_308_clk),
    .Q(\dp.rf.rf[25][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][18]$_DFFE_PP_  (.D(_00556_),
    .CLK(clknet_leaf_89_clk),
    .Q(\dp.rf.rf[25][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][19]$_DFFE_PP_  (.D(_00557_),
    .CLK(clknet_leaf_85_clk),
    .Q(\dp.rf.rf[25][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][1]$_DFFE_PP_  (.D(_00558_),
    .CLK(clknet_leaf_513_clk),
    .Q(\dp.rf.rf[25][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][20]$_DFFE_PP_  (.D(_00559_),
    .CLK(clknet_leaf_411_clk),
    .Q(\dp.rf.rf[25][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][21]$_DFFE_PP_  (.D(_00560_),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\dp.rf.rf[25][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][22]$_DFFE_PP_  (.D(_00561_),
    .CLK(clknet_leaf_649_clk),
    .Q(\dp.rf.rf[25][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][23]$_DFFE_PP_  (.D(_00562_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[25][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][24]$_DFFE_PP_  (.D(_00563_),
    .CLK(clknet_leaf_638_clk),
    .Q(\dp.rf.rf[25][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][25]$_DFFE_PP_  (.D(_00564_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[25][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][26]$_DFFE_PP_  (.D(_00565_),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\dp.rf.rf[25][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][27]$_DFFE_PP_  (.D(_00566_),
    .CLK(clknet_leaf_486_clk),
    .Q(\dp.rf.rf[25][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][28]$_DFFE_PP_  (.D(_00567_),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\dp.rf.rf[25][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][29]$_DFFE_PP_  (.D(_00568_),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\dp.rf.rf[25][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][2]$_DFFE_PP_  (.D(_00569_),
    .CLK(clknet_leaf_25_clk),
    .Q(\dp.rf.rf[25][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][30]$_DFFE_PP_  (.D(_00570_),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\dp.rf.rf[25][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][31]$_DFFE_PP_  (.D(_00571_),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\dp.rf.rf[25][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][3]$_DFFE_PP_  (.D(_00572_),
    .CLK(clknet_leaf_179_clk),
    .Q(\dp.rf.rf[25][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][4]$_DFFE_PP_  (.D(_00573_),
    .CLK(clknet_leaf_626_clk),
    .Q(\dp.rf.rf[25][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][5]$_DFFE_PP_  (.D(_00574_),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\dp.rf.rf[25][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][6]$_DFFE_PP_  (.D(_00575_),
    .CLK(clknet_leaf_408_clk),
    .Q(\dp.rf.rf[25][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][7]$_DFFE_PP_  (.D(_00576_),
    .CLK(clknet_leaf_56_clk),
    .Q(\dp.rf.rf[25][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][8]$_DFFE_PP_  (.D(_00577_),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\dp.rf.rf[25][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[25][9]$_DFFE_PP_  (.D(_00578_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\dp.rf.rf[25][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][0]$_DFFE_PP_  (.D(_00579_),
    .CLK(clknet_leaf_324_clk),
    .Q(\dp.rf.rf[26][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][10]$_DFFE_PP_  (.D(_00580_),
    .CLK(clknet_leaf_281_clk),
    .Q(\dp.rf.rf[26][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][11]$_DFFE_PP_  (.D(_00581_),
    .CLK(clknet_leaf_282_clk),
    .Q(\dp.rf.rf[26][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][12]$_DFFE_PP_  (.D(_00582_),
    .CLK(clknet_leaf_121_clk),
    .Q(\dp.rf.rf[26][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][13]$_DFFE_PP_  (.D(_00583_),
    .CLK(clknet_leaf_215_clk),
    .Q(\dp.rf.rf[26][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][14]$_DFFE_PP_  (.D(_00584_),
    .CLK(clknet_leaf_243_clk),
    .Q(\dp.rf.rf[26][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][15]$_DFFE_PP_  (.D(_00585_),
    .CLK(clknet_leaf_190_clk),
    .Q(\dp.rf.rf[26][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][16]$_DFFE_PP_  (.D(_00586_),
    .CLK(clknet_leaf_290_clk),
    .Q(\dp.rf.rf[26][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][17]$_DFFE_PP_  (.D(_00587_),
    .CLK(clknet_leaf_294_clk),
    .Q(\dp.rf.rf[26][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][18]$_DFFE_PP_  (.D(_00588_),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\dp.rf.rf[26][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][19]$_DFFE_PP_  (.D(_00589_),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\dp.rf.rf[26][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][1]$_DFFE_PP_  (.D(_00590_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[26][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][20]$_DFFE_PP_  (.D(_00591_),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\dp.rf.rf[26][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][21]$_DFFE_PP_  (.D(_00592_),
    .CLK(clknet_leaf_697_clk),
    .Q(\dp.rf.rf[26][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][22]$_DFFE_PP_  (.D(_00593_),
    .CLK(clknet_6_1__leaf_clk),
    .Q(\dp.rf.rf[26][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][23]$_DFFE_PP_  (.D(_00594_),
    .CLK(clknet_leaf_430_clk),
    .Q(\dp.rf.rf[26][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][24]$_DFFE_PP_  (.D(_00595_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\dp.rf.rf[26][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][25]$_DFFE_PP_  (.D(_00596_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[26][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][26]$_DFFE_PP_  (.D(_00597_),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\dp.rf.rf[26][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][27]$_DFFE_PP_  (.D(_00598_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[26][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][28]$_DFFE_PP_  (.D(_00599_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[26][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][29]$_DFFE_PP_  (.D(_00600_),
    .CLK(clknet_leaf_438_clk),
    .Q(\dp.rf.rf[26][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][2]$_DFFE_PP_  (.D(_00601_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[26][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][30]$_DFFE_PP_  (.D(_00602_),
    .CLK(clknet_leaf_611_clk),
    .Q(\dp.rf.rf[26][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][31]$_DFFE_PP_  (.D(_00603_),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\dp.rf.rf[26][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][3]$_DFFE_PP_  (.D(_00604_),
    .CLK(clknet_leaf_179_clk),
    .Q(\dp.rf.rf[26][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][4]$_DFFE_PP_  (.D(_00605_),
    .CLK(clknet_leaf_623_clk),
    .Q(\dp.rf.rf[26][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][5]$_DFFE_PP_  (.D(_00606_),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\dp.rf.rf[26][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][6]$_DFFE_PP_  (.D(_00607_),
    .CLK(clknet_leaf_403_clk),
    .Q(\dp.rf.rf[26][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][7]$_DFFE_PP_  (.D(_00608_),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\dp.rf.rf[26][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][8]$_DFFE_PP_  (.D(_00609_),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\dp.rf.rf[26][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[26][9]$_DFFE_PP_  (.D(_00610_),
    .CLK(clknet_leaf_633_clk),
    .Q(\dp.rf.rf[26][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][0]$_DFFE_PP_  (.D(_00611_),
    .CLK(clknet_leaf_324_clk),
    .Q(\dp.rf.rf[27][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][10]$_DFFE_PP_  (.D(_00612_),
    .CLK(clknet_leaf_310_clk),
    .Q(\dp.rf.rf[27][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][11]$_DFFE_PP_  (.D(_00613_),
    .CLK(clknet_leaf_282_clk),
    .Q(\dp.rf.rf[27][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][12]$_DFFE_PP_  (.D(_00614_),
    .CLK(clknet_leaf_121_clk),
    .Q(\dp.rf.rf[27][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][13]$_DFFE_PP_  (.D(_00615_),
    .CLK(clknet_leaf_215_clk),
    .Q(\dp.rf.rf[27][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][14]$_DFFE_PP_  (.D(_00616_),
    .CLK(clknet_leaf_243_clk),
    .Q(\dp.rf.rf[27][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][15]$_DFFE_PP_  (.D(_00617_),
    .CLK(clknet_leaf_190_clk),
    .Q(\dp.rf.rf[27][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][16]$_DFFE_PP_  (.D(_00618_),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\dp.rf.rf[27][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][17]$_DFFE_PP_  (.D(_00619_),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\dp.rf.rf[27][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][18]$_DFFE_PP_  (.D(_00620_),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\dp.rf.rf[27][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][19]$_DFFE_PP_  (.D(_00621_),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\dp.rf.rf[27][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][1]$_DFFE_PP_  (.D(_00622_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[27][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][20]$_DFFE_PP_  (.D(_00623_),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\dp.rf.rf[27][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][21]$_DFFE_PP_  (.D(_00624_),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\dp.rf.rf[27][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][22]$_DFFE_PP_  (.D(_00625_),
    .CLK(clknet_leaf_645_clk),
    .Q(\dp.rf.rf[27][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][23]$_DFFE_PP_  (.D(_00626_),
    .CLK(clknet_leaf_430_clk),
    .Q(\dp.rf.rf[27][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][24]$_DFFE_PP_  (.D(_00627_),
    .CLK(clknet_leaf_645_clk),
    .Q(\dp.rf.rf[27][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][25]$_DFFE_PP_  (.D(_00628_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[27][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][26]$_DFFE_PP_  (.D(_00629_),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\dp.rf.rf[27][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][27]$_DFFE_PP_  (.D(_00630_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[27][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][28]$_DFFE_PP_  (.D(_00631_),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\dp.rf.rf[27][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][29]$_DFFE_PP_  (.D(_00632_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\dp.rf.rf[27][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][2]$_DFFE_PP_  (.D(_00633_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[27][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][30]$_DFFE_PP_  (.D(_00634_),
    .CLK(clknet_leaf_611_clk),
    .Q(\dp.rf.rf[27][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][31]$_DFFE_PP_  (.D(_00635_),
    .CLK(clknet_leaf_390_clk),
    .Q(\dp.rf.rf[27][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][3]$_DFFE_PP_  (.D(_00636_),
    .CLK(clknet_leaf_170_clk),
    .Q(\dp.rf.rf[27][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][4]$_DFFE_PP_  (.D(_00637_),
    .CLK(clknet_leaf_624_clk),
    .Q(\dp.rf.rf[27][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][5]$_DFFE_PP_  (.D(_00638_),
    .CLK(clknet_leaf_134_clk),
    .Q(\dp.rf.rf[27][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][6]$_DFFE_PP_  (.D(_00639_),
    .CLK(clknet_leaf_403_clk),
    .Q(\dp.rf.rf[27][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][7]$_DFFE_PP_  (.D(_00640_),
    .CLK(clknet_leaf_58_clk),
    .Q(\dp.rf.rf[27][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][8]$_DFFE_PP_  (.D(_00641_),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\dp.rf.rf[27][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[27][9]$_DFFE_PP_  (.D(_00642_),
    .CLK(clknet_leaf_633_clk),
    .Q(\dp.rf.rf[27][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][0]$_DFFE_PP_  (.D(_00643_),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\dp.rf.rf[28][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][10]$_DFFE_PP_  (.D(_00644_),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\dp.rf.rf[28][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][11]$_DFFE_PP_  (.D(_00645_),
    .CLK(clknet_leaf_284_clk),
    .Q(\dp.rf.rf[28][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][12]$_DFFE_PP_  (.D(_00646_),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\dp.rf.rf[28][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][13]$_DFFE_PP_  (.D(_00647_),
    .CLK(clknet_leaf_211_clk),
    .Q(\dp.rf.rf[28][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][14]$_DFFE_PP_  (.D(_00648_),
    .CLK(clknet_leaf_249_clk),
    .Q(\dp.rf.rf[28][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][15]$_DFFE_PP_  (.D(_00649_),
    .CLK(clknet_leaf_251_clk),
    .Q(\dp.rf.rf[28][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][16]$_DFFE_PP_  (.D(_00650_),
    .CLK(clknet_leaf_290_clk),
    .Q(\dp.rf.rf[28][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][17]$_DFFE_PP_  (.D(_00651_),
    .CLK(clknet_leaf_309_clk),
    .Q(\dp.rf.rf[28][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][18]$_DFFE_PP_  (.D(_00652_),
    .CLK(clknet_leaf_65_clk),
    .Q(\dp.rf.rf[28][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][19]$_DFFE_PP_  (.D(_00653_),
    .CLK(clknet_leaf_88_clk),
    .Q(\dp.rf.rf[28][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][1]$_DFFE_PP_  (.D(_00654_),
    .CLK(clknet_leaf_515_clk),
    .Q(\dp.rf.rf[28][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][20]$_DFFE_PP_  (.D(_00655_),
    .CLK(clknet_leaf_413_clk),
    .Q(\dp.rf.rf[28][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][21]$_DFFE_PP_  (.D(_00656_),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\dp.rf.rf[28][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][22]$_DFFE_PP_  (.D(_00657_),
    .CLK(clknet_6_1__leaf_clk),
    .Q(\dp.rf.rf[28][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][23]$_DFFE_PP_  (.D(_00658_),
    .CLK(clknet_leaf_383_clk),
    .Q(\dp.rf.rf[28][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][24]$_DFFE_PP_  (.D(_00659_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\dp.rf.rf[28][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][25]$_DFFE_PP_  (.D(_00660_),
    .CLK(clknet_leaf_385_clk),
    .Q(\dp.rf.rf[28][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][26]$_DFFE_PP_  (.D(_00661_),
    .CLK(clknet_leaf_712_clk),
    .Q(\dp.rf.rf[28][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][27]$_DFFE_PP_  (.D(_00662_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[28][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][28]$_DFFE_PP_  (.D(_00663_),
    .CLK(clknet_leaf_664_clk),
    .Q(\dp.rf.rf[28][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][29]$_DFFE_PP_  (.D(_00664_),
    .CLK(clknet_leaf_375_clk),
    .Q(\dp.rf.rf[28][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][2]$_DFFE_PP_  (.D(_00665_),
    .CLK(clknet_leaf_26_clk),
    .Q(\dp.rf.rf[28][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][30]$_DFFE_PP_  (.D(_00666_),
    .CLK(clknet_leaf_609_clk),
    .Q(\dp.rf.rf[28][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][31]$_DFFE_PP_  (.D(_00667_),
    .CLK(clknet_leaf_296_clk),
    .Q(\dp.rf.rf[28][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][3]$_DFFE_PP_  (.D(_00668_),
    .CLK(clknet_6_58__leaf_clk),
    .Q(\dp.rf.rf[28][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][4]$_DFFE_PP_  (.D(_00669_),
    .CLK(clknet_leaf_618_clk),
    .Q(\dp.rf.rf[28][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][5]$_DFFE_PP_  (.D(_00670_),
    .CLK(clknet_leaf_136_clk),
    .Q(\dp.rf.rf[28][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][6]$_DFFE_PP_  (.D(_00671_),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\dp.rf.rf[28][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][7]$_DFFE_PP_  (.D(_00672_),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\dp.rf.rf[28][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][8]$_DFFE_PP_  (.D(_00673_),
    .CLK(clknet_leaf_404_clk),
    .Q(\dp.rf.rf[28][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[28][9]$_DFFE_PP_  (.D(_00674_),
    .CLK(clknet_leaf_622_clk),
    .Q(\dp.rf.rf[28][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][0]$_DFFE_PP_  (.D(_00675_),
    .CLK(clknet_leaf_175_clk),
    .Q(\dp.rf.rf[29][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][10]$_DFFE_PP_  (.D(_00676_),
    .CLK(clknet_leaf_310_clk),
    .Q(\dp.rf.rf[29][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][11]$_DFFE_PP_  (.D(_00677_),
    .CLK(clknet_leaf_281_clk),
    .Q(\dp.rf.rf[29][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][12]$_DFFE_PP_  (.D(_00678_),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\dp.rf.rf[29][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][13]$_DFFE_PP_  (.D(_00679_),
    .CLK(clknet_leaf_232_clk),
    .Q(\dp.rf.rf[29][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][14]$_DFFE_PP_  (.D(_00680_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\dp.rf.rf[29][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][15]$_DFFE_PP_  (.D(_00681_),
    .CLK(clknet_leaf_187_clk),
    .Q(\dp.rf.rf[29][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][16]$_DFFE_PP_  (.D(_00682_),
    .CLK(clknet_leaf_295_clk),
    .Q(\dp.rf.rf[29][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][17]$_DFFE_PP_  (.D(_00683_),
    .CLK(clknet_leaf_308_clk),
    .Q(\dp.rf.rf[29][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][18]$_DFFE_PP_  (.D(_00684_),
    .CLK(clknet_leaf_65_clk),
    .Q(\dp.rf.rf[29][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][19]$_DFFE_PP_  (.D(_00685_),
    .CLK(clknet_leaf_87_clk),
    .Q(\dp.rf.rf[29][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][1]$_DFFE_PP_  (.D(_00686_),
    .CLK(clknet_leaf_515_clk),
    .Q(\dp.rf.rf[29][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][20]$_DFFE_PP_  (.D(_00687_),
    .CLK(clknet_leaf_413_clk),
    .Q(\dp.rf.rf[29][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][21]$_DFFE_PP_  (.D(_00688_),
    .CLK(clknet_leaf_697_clk),
    .Q(\dp.rf.rf[29][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][22]$_DFFE_PP_  (.D(_00689_),
    .CLK(clknet_6_1__leaf_clk),
    .Q(\dp.rf.rf[29][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][23]$_DFFE_PP_  (.D(_00690_),
    .CLK(clknet_leaf_383_clk),
    .Q(\dp.rf.rf[29][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][24]$_DFFE_PP_  (.D(_00691_),
    .CLK(clknet_leaf_654_clk),
    .Q(\dp.rf.rf[29][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][25]$_DFFE_PP_  (.D(_00692_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\dp.rf.rf[29][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][26]$_DFFE_PP_  (.D(_00693_),
    .CLK(clknet_leaf_712_clk),
    .Q(\dp.rf.rf[29][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][27]$_DFFE_PP_  (.D(_00694_),
    .CLK(clknet_leaf_486_clk),
    .Q(\dp.rf.rf[29][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][28]$_DFFE_PP_  (.D(_00695_),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\dp.rf.rf[29][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][29]$_DFFE_PP_  (.D(_00696_),
    .CLK(clknet_leaf_375_clk),
    .Q(\dp.rf.rf[29][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][2]$_DFFE_PP_  (.D(_00697_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[29][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][30]$_DFFE_PP_  (.D(_00698_),
    .CLK(clknet_leaf_609_clk),
    .Q(\dp.rf.rf[29][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][31]$_DFFE_PP_  (.D(_00699_),
    .CLK(clknet_leaf_393_clk),
    .Q(\dp.rf.rf[29][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][3]$_DFFE_PP_  (.D(_00700_),
    .CLK(clknet_leaf_177_clk),
    .Q(\dp.rf.rf[29][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][4]$_DFFE_PP_  (.D(_00701_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\dp.rf.rf[29][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][5]$_DFFE_PP_  (.D(_00702_),
    .CLK(clknet_leaf_134_clk),
    .Q(\dp.rf.rf[29][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][6]$_DFFE_PP_  (.D(_00703_),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\dp.rf.rf[29][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][7]$_DFFE_PP_  (.D(_00704_),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\dp.rf.rf[29][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][8]$_DFFE_PP_  (.D(_00705_),
    .CLK(clknet_leaf_404_clk),
    .Q(\dp.rf.rf[29][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[29][9]$_DFFE_PP_  (.D(_00706_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\dp.rf.rf[29][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][0]$_DFFE_PP_  (.D(_00707_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\dp.rf.rf[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][10]$_DFFE_PP_  (.D(_00708_),
    .CLK(clknet_leaf_271_clk),
    .Q(\dp.rf.rf[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][11]$_DFFE_PP_  (.D(_00709_),
    .CLK(clknet_leaf_267_clk),
    .Q(\dp.rf.rf[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][12]$_DFFE_PP_  (.D(_00710_),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\dp.rf.rf[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][13]$_DFFE_PP_  (.D(_00711_),
    .CLK(clknet_leaf_220_clk),
    .Q(\dp.rf.rf[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][14]$_DFFE_PP_  (.D(_00712_),
    .CLK(clknet_leaf_231_clk),
    .Q(\dp.rf.rf[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][15]$_DFFE_PP_  (.D(_00713_),
    .CLK(clknet_leaf_256_clk),
    .Q(\dp.rf.rf[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][16]$_DFFE_PP_  (.D(_00714_),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\dp.rf.rf[2][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][17]$_DFFE_PP_  (.D(_00715_),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\dp.rf.rf[2][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][18]$_DFFE_PP_  (.D(_00716_),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\dp.rf.rf[2][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][19]$_DFFE_PP_  (.D(_00717_),
    .CLK(clknet_leaf_114_clk),
    .Q(\dp.rf.rf[2][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][1]$_DFFE_PP_  (.D(_00718_),
    .CLK(clknet_leaf_502_clk),
    .Q(\dp.rf.rf[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][20]$_DFFE_PP_  (.D(_00719_),
    .CLK(clknet_leaf_449_clk),
    .Q(\dp.rf.rf[2][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][21]$_DFFE_PP_  (.D(_00720_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\dp.rf.rf[2][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][22]$_DFFE_PP_  (.D(_00721_),
    .CLK(clknet_leaf_680_clk),
    .Q(\dp.rf.rf[2][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][23]$_DFFE_PP_  (.D(_00722_),
    .CLK(clknet_leaf_481_clk),
    .Q(\dp.rf.rf[2][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][24]$_DFFE_PP_  (.D(_00723_),
    .CLK(clknet_leaf_678_clk),
    .Q(\dp.rf.rf[2][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][25]$_DFFE_PP_  (.D(_00724_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[2][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][26]$_DFFE_PP_  (.D(_00725_),
    .CLK(clknet_leaf_668_clk),
    .Q(\dp.rf.rf[2][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][27]$_DFFE_PP_  (.D(_00726_),
    .CLK(clknet_leaf_494_clk),
    .Q(\dp.rf.rf[2][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][28]$_DFFE_PP_  (.D(_00727_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[2][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][29]$_DFFE_PP_  (.D(_00728_),
    .CLK(clknet_leaf_545_clk),
    .Q(\dp.rf.rf[2][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][2]$_DFFE_PP_  (.D(_00729_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][30]$_DFFE_PP_  (.D(_00730_),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\dp.rf.rf[2][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][31]$_DFFE_PP_  (.D(_00731_),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\dp.rf.rf[2][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][3]$_DFFE_PP_  (.D(_00732_),
    .CLK(clknet_leaf_163_clk),
    .Q(\dp.rf.rf[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][4]$_DFFE_PP_  (.D(_00733_),
    .CLK(clknet_leaf_629_clk),
    .Q(\dp.rf.rf[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][5]$_DFFE_PP_  (.D(_00734_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\dp.rf.rf[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][6]$_DFFE_PP_  (.D(_00735_),
    .CLK(clknet_leaf_454_clk),
    .Q(\dp.rf.rf[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][7]$_DFFE_PP_  (.D(_00736_),
    .CLK(clknet_leaf_112_clk),
    .Q(\dp.rf.rf[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][8]$_DFFE_PP_  (.D(_00737_),
    .CLK(clknet_leaf_442_clk),
    .Q(\dp.rf.rf[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[2][9]$_DFFE_PP_  (.D(_00738_),
    .CLK(clknet_leaf_641_clk),
    .Q(\dp.rf.rf[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][0]$_DFFE_PP_  (.D(_00739_),
    .CLK(clknet_leaf_176_clk),
    .Q(\dp.rf.rf[30][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][10]$_DFFE_PP_  (.D(_00740_),
    .CLK(clknet_leaf_315_clk),
    .Q(\dp.rf.rf[30][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][11]$_DFFE_PP_  (.D(_00741_),
    .CLK(clknet_leaf_316_clk),
    .Q(\dp.rf.rf[30][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][12]$_DFFE_PP_  (.D(_00742_),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\dp.rf.rf[30][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][13]$_DFFE_PP_  (.D(_00743_),
    .CLK(clknet_leaf_216_clk),
    .Q(\dp.rf.rf[30][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][14]$_DFFE_PP_  (.D(_00744_),
    .CLK(clknet_leaf_244_clk),
    .Q(\dp.rf.rf[30][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][15]$_DFFE_PP_  (.D(_00745_),
    .CLK(clknet_leaf_189_clk),
    .Q(\dp.rf.rf[30][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][16]$_DFFE_PP_  (.D(_00746_),
    .CLK(clknet_leaf_296_clk),
    .Q(\dp.rf.rf[30][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][17]$_DFFE_PP_  (.D(_00747_),
    .CLK(clknet_leaf_307_clk),
    .Q(\dp.rf.rf[30][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][18]$_DFFE_PP_  (.D(_00748_),
    .CLK(clknet_leaf_64_clk),
    .Q(\dp.rf.rf[30][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][19]$_DFFE_PP_  (.D(_00749_),
    .CLK(clknet_leaf_89_clk),
    .Q(\dp.rf.rf[30][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][1]$_DFFE_PP_  (.D(_00750_),
    .CLK(clknet_leaf_516_clk),
    .Q(\dp.rf.rf[30][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][20]$_DFFE_PP_  (.D(_00751_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[30][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][21]$_DFFE_PP_  (.D(_00752_),
    .CLK(clknet_leaf_698_clk),
    .Q(\dp.rf.rf[30][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][22]$_DFFE_PP_  (.D(_00753_),
    .CLK(clknet_6_1__leaf_clk),
    .Q(\dp.rf.rf[30][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][23]$_DFFE_PP_  (.D(_00754_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\dp.rf.rf[30][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][24]$_DFFE_PP_  (.D(_00755_),
    .CLK(clknet_leaf_652_clk),
    .Q(\dp.rf.rf[30][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][25]$_DFFE_PP_  (.D(_00756_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\dp.rf.rf[30][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][26]$_DFFE_PP_  (.D(_00757_),
    .CLK(clknet_leaf_711_clk),
    .Q(\dp.rf.rf[30][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][27]$_DFFE_PP_  (.D(_00758_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[30][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][28]$_DFFE_PP_  (.D(_00759_),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\dp.rf.rf[30][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][29]$_DFFE_PP_  (.D(_00760_),
    .CLK(clknet_leaf_374_clk),
    .Q(\dp.rf.rf[30][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][2]$_DFFE_PP_  (.D(_00761_),
    .CLK(clknet_leaf_27_clk),
    .Q(\dp.rf.rf[30][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][30]$_DFFE_PP_  (.D(_00762_),
    .CLK(clknet_leaf_608_clk),
    .Q(\dp.rf.rf[30][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][31]$_DFFE_PP_  (.D(_00763_),
    .CLK(clknet_leaf_393_clk),
    .Q(\dp.rf.rf[30][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][3]$_DFFE_PP_  (.D(_00764_),
    .CLK(clknet_leaf_171_clk),
    .Q(\dp.rf.rf[30][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][4]$_DFFE_PP_  (.D(_00765_),
    .CLK(clknet_leaf_624_clk),
    .Q(\dp.rf.rf[30][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][5]$_DFFE_PP_  (.D(_00766_),
    .CLK(clknet_leaf_137_clk),
    .Q(\dp.rf.rf[30][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][6]$_DFFE_PP_  (.D(_00767_),
    .CLK(clknet_leaf_396_clk),
    .Q(\dp.rf.rf[30][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][7]$_DFFE_PP_  (.D(_00768_),
    .CLK(clknet_leaf_60_clk),
    .Q(\dp.rf.rf[30][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][8]$_DFFE_PP_  (.D(_00769_),
    .CLK(clknet_leaf_394_clk),
    .Q(\dp.rf.rf[30][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[30][9]$_DFFE_PP_  (.D(_00770_),
    .CLK(clknet_leaf_637_clk),
    .Q(\dp.rf.rf[30][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][0]$_DFFE_PP_  (.D(_00771_),
    .CLK(clknet_leaf_176_clk),
    .Q(\dp.rf.rf[31][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][10]$_DFFE_PP_  (.D(_00772_),
    .CLK(clknet_leaf_315_clk),
    .Q(\dp.rf.rf[31][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][11]$_DFFE_PP_  (.D(_00773_),
    .CLK(clknet_leaf_280_clk),
    .Q(\dp.rf.rf[31][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][12]$_DFFE_PP_  (.D(_00774_),
    .CLK(clknet_leaf_118_clk),
    .Q(\dp.rf.rf[31][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][13]$_DFFE_PP_  (.D(_00775_),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\dp.rf.rf[31][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][14]$_DFFE_PP_  (.D(_00776_),
    .CLK(clknet_leaf_244_clk),
    .Q(\dp.rf.rf[31][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][15]$_DFFE_PP_  (.D(_00777_),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\dp.rf.rf[31][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][16]$_DFFE_PP_  (.D(_00778_),
    .CLK(clknet_leaf_295_clk),
    .Q(\dp.rf.rf[31][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][17]$_DFFE_PP_  (.D(_00779_),
    .CLK(clknet_leaf_307_clk),
    .Q(\dp.rf.rf[31][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][18]$_DFFE_PP_  (.D(_00780_),
    .CLK(clknet_leaf_64_clk),
    .Q(\dp.rf.rf[31][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][19]$_DFFE_PP_  (.D(_00781_),
    .CLK(clknet_leaf_88_clk),
    .Q(\dp.rf.rf[31][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][1]$_DFFE_PP_  (.D(_00782_),
    .CLK(clknet_leaf_516_clk),
    .Q(\dp.rf.rf[31][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][20]$_DFFE_PP_  (.D(_00783_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[31][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][21]$_DFFE_PP_  (.D(_00784_),
    .CLK(clknet_leaf_698_clk),
    .Q(\dp.rf.rf[31][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][22]$_DFFE_PP_  (.D(_00785_),
    .CLK(clknet_6_1__leaf_clk),
    .Q(\dp.rf.rf[31][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][23]$_DFFE_PP_  (.D(_00786_),
    .CLK(clknet_leaf_380_clk),
    .Q(\dp.rf.rf[31][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][24]$_DFFE_PP_  (.D(_00787_),
    .CLK(clknet_leaf_652_clk),
    .Q(\dp.rf.rf[31][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][25]$_DFFE_PP_  (.D(_00788_),
    .CLK(clknet_leaf_385_clk),
    .Q(\dp.rf.rf[31][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][26]$_DFFE_PP_  (.D(_00789_),
    .CLK(clknet_leaf_711_clk),
    .Q(\dp.rf.rf[31][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][27]$_DFFE_PP_  (.D(_00790_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[31][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][28]$_DFFE_PP_  (.D(_00791_),
    .CLK(clknet_leaf_14_clk),
    .Q(\dp.rf.rf[31][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][29]$_DFFE_PP_  (.D(_00792_),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\dp.rf.rf[31][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][2]$_DFFE_PP_  (.D(_00793_),
    .CLK(clknet_leaf_28_clk),
    .Q(\dp.rf.rf[31][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][30]$_DFFE_PP_  (.D(_00794_),
    .CLK(clknet_leaf_608_clk),
    .Q(\dp.rf.rf[31][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][31]$_DFFE_PP_  (.D(_00795_),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\dp.rf.rf[31][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][3]$_DFFE_PP_  (.D(_00796_),
    .CLK(clknet_leaf_171_clk),
    .Q(\dp.rf.rf[31][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][4]$_DFFE_PP_  (.D(_00797_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\dp.rf.rf[31][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][5]$_DFFE_PP_  (.D(_00798_),
    .CLK(clknet_leaf_137_clk),
    .Q(\dp.rf.rf[31][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][6]$_DFFE_PP_  (.D(_00799_),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\dp.rf.rf[31][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][7]$_DFFE_PP_  (.D(_00800_),
    .CLK(clknet_leaf_60_clk),
    .Q(\dp.rf.rf[31][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][8]$_DFFE_PP_  (.D(_00801_),
    .CLK(clknet_leaf_394_clk),
    .Q(\dp.rf.rf[31][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[31][9]$_DFFE_PP_  (.D(_00802_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\dp.rf.rf[31][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][0]$_DFFE_PP_  (.D(_00803_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\dp.rf.rf[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][10]$_DFFE_PP_  (.D(_00804_),
    .CLK(clknet_leaf_271_clk),
    .Q(\dp.rf.rf[3][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][11]$_DFFE_PP_  (.D(_00805_),
    .CLK(clknet_leaf_267_clk),
    .Q(\dp.rf.rf[3][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][12]$_DFFE_PP_  (.D(_00806_),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\dp.rf.rf[3][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][13]$_DFFE_PP_  (.D(_00807_),
    .CLK(clknet_leaf_220_clk),
    .Q(\dp.rf.rf[3][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][14]$_DFFE_PP_  (.D(_00808_),
    .CLK(clknet_leaf_230_clk),
    .Q(\dp.rf.rf[3][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][15]$_DFFE_PP_  (.D(_00809_),
    .CLK(clknet_leaf_256_clk),
    .Q(\dp.rf.rf[3][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][16]$_DFFE_PP_  (.D(_00810_),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\dp.rf.rf[3][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][17]$_DFFE_PP_  (.D(_00811_),
    .CLK(clknet_leaf_308_clk),
    .Q(\dp.rf.rf[3][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][18]$_DFFE_PP_  (.D(_00812_),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\dp.rf.rf[3][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][19]$_DFFE_PP_  (.D(_00813_),
    .CLK(clknet_leaf_114_clk),
    .Q(\dp.rf.rf[3][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][1]$_DFFE_PP_  (.D(_00814_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][20]$_DFFE_PP_  (.D(_00815_),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\dp.rf.rf[3][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][21]$_DFFE_PP_  (.D(_00816_),
    .CLK(clknet_leaf_685_clk),
    .Q(\dp.rf.rf[3][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][22]$_DFFE_PP_  (.D(_00817_),
    .CLK(clknet_leaf_680_clk),
    .Q(\dp.rf.rf[3][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][23]$_DFFE_PP_  (.D(_00818_),
    .CLK(clknet_leaf_481_clk),
    .Q(\dp.rf.rf[3][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][24]$_DFFE_PP_  (.D(_00819_),
    .CLK(clknet_leaf_678_clk),
    .Q(\dp.rf.rf[3][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][25]$_DFFE_PP_  (.D(_00820_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[3][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][26]$_DFFE_PP_  (.D(_00821_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\dp.rf.rf[3][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][27]$_DFFE_PP_  (.D(_00822_),
    .CLK(clknet_leaf_494_clk),
    .Q(\dp.rf.rf[3][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][28]$_DFFE_PP_  (.D(_00823_),
    .CLK(clknet_leaf_11_clk),
    .Q(\dp.rf.rf[3][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][29]$_DFFE_PP_  (.D(_00824_),
    .CLK(clknet_leaf_546_clk),
    .Q(\dp.rf.rf[3][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][2]$_DFFE_PP_  (.D(_00825_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][30]$_DFFE_PP_  (.D(_00826_),
    .CLK(clknet_leaf_578_clk),
    .Q(\dp.rf.rf[3][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][31]$_DFFE_PP_  (.D(_00827_),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\dp.rf.rf[3][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][3]$_DFFE_PP_  (.D(_00828_),
    .CLK(clknet_leaf_163_clk),
    .Q(\dp.rf.rf[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][4]$_DFFE_PP_  (.D(_00829_),
    .CLK(clknet_leaf_629_clk),
    .Q(\dp.rf.rf[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][5]$_DFFE_PP_  (.D(_00830_),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\dp.rf.rf[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][6]$_DFFE_PP_  (.D(_00831_),
    .CLK(clknet_leaf_424_clk),
    .Q(\dp.rf.rf[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][7]$_DFFE_PP_  (.D(_00832_),
    .CLK(clknet_leaf_112_clk),
    .Q(\dp.rf.rf[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][8]$_DFFE_PP_  (.D(_00833_),
    .CLK(clknet_leaf_446_clk),
    .Q(\dp.rf.rf[3][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[3][9]$_DFFE_PP_  (.D(_00834_),
    .CLK(clknet_leaf_641_clk),
    .Q(\dp.rf.rf[3][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][0]$_DFFE_PP_  (.D(_00835_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\dp.rf.rf[4][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][10]$_DFFE_PP_  (.D(_00836_),
    .CLK(clknet_leaf_242_clk),
    .Q(\dp.rf.rf[4][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][11]$_DFFE_PP_  (.D(_00837_),
    .CLK(clknet_leaf_248_clk),
    .Q(\dp.rf.rf[4][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][12]$_DFFE_PP_  (.D(_00838_),
    .CLK(clknet_leaf_200_clk),
    .Q(\dp.rf.rf[4][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][13]$_DFFE_PP_  (.D(_00839_),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\dp.rf.rf[4][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][14]$_DFFE_PP_  (.D(_00840_),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\dp.rf.rf[4][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][15]$_DFFE_PP_  (.D(_00841_),
    .CLK(clknet_leaf_251_clk),
    .Q(\dp.rf.rf[4][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][16]$_DFFE_PP_  (.D(_00842_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\dp.rf.rf[4][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][17]$_DFFE_PP_  (.D(_00843_),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\dp.rf.rf[4][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][18]$_DFFE_PP_  (.D(_00844_),
    .CLK(clknet_leaf_103_clk),
    .Q(\dp.rf.rf[4][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][19]$_DFFE_PP_  (.D(_00845_),
    .CLK(clknet_leaf_102_clk),
    .Q(\dp.rf.rf[4][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][1]$_DFFE_PP_  (.D(_00846_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\dp.rf.rf[4][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][20]$_DFFE_PP_  (.D(_00847_),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\dp.rf.rf[4][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][21]$_DFFE_PP_  (.D(_00848_),
    .CLK(clknet_6_0__leaf_clk),
    .Q(\dp.rf.rf[4][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][22]$_DFFE_PP_  (.D(_00849_),
    .CLK(clknet_6_0__leaf_clk),
    .Q(\dp.rf.rf[4][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][23]$_DFFE_PP_  (.D(_00850_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[4][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][24]$_DFFE_PP_  (.D(_00851_),
    .CLK(clknet_leaf_673_clk),
    .Q(\dp.rf.rf[4][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][25]$_DFFE_PP_  (.D(_00852_),
    .CLK(clknet_leaf_546_clk),
    .Q(\dp.rf.rf[4][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][26]$_DFFE_PP_  (.D(_00853_),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\dp.rf.rf[4][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][27]$_DFFE_PP_  (.D(_00854_),
    .CLK(clknet_leaf_488_clk),
    .Q(\dp.rf.rf[4][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][28]$_DFFE_PP_  (.D(_00855_),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\dp.rf.rf[4][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][29]$_DFFE_PP_  (.D(_00856_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[4][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][2]$_DFFE_PP_  (.D(_00857_),
    .CLK(clknet_leaf_13_clk),
    .Q(\dp.rf.rf[4][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][30]$_DFFE_PP_  (.D(_00858_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[4][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][31]$_DFFE_PP_  (.D(_00859_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[4][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][3]$_DFFE_PP_  (.D(_00860_),
    .CLK(clknet_leaf_165_clk),
    .Q(\dp.rf.rf[4][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][4]$_DFFE_PP_  (.D(_00861_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\dp.rf.rf[4][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][5]$_DFFE_PP_  (.D(_00862_),
    .CLK(clknet_leaf_137_clk),
    .Q(\dp.rf.rf[4][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][6]$_DFFE_PP_  (.D(_00863_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[4][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][7]$_DFFE_PP_  (.D(_00864_),
    .CLK(clknet_leaf_103_clk),
    .Q(\dp.rf.rf[4][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][8]$_DFFE_PP_  (.D(_00865_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[4][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[4][9]$_DFFE_PP_  (.D(_00866_),
    .CLK(clknet_leaf_637_clk),
    .Q(\dp.rf.rf[4][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][0]$_DFFE_PP_  (.D(_00867_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\dp.rf.rf[5][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][10]$_DFFE_PP_  (.D(_00868_),
    .CLK(clknet_leaf_267_clk),
    .Q(\dp.rf.rf[5][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][11]$_DFFE_PP_  (.D(_00869_),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\dp.rf.rf[5][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][12]$_DFFE_PP_  (.D(_00870_),
    .CLK(clknet_6_32__leaf_clk),
    .Q(\dp.rf.rf[5][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][13]$_DFFE_PP_  (.D(_00871_),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\dp.rf.rf[5][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][14]$_DFFE_PP_  (.D(_00872_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\dp.rf.rf[5][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][15]$_DFFE_PP_  (.D(_00873_),
    .CLK(clknet_leaf_253_clk),
    .Q(\dp.rf.rf[5][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][16]$_DFFE_PP_  (.D(_00874_),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\dp.rf.rf[5][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][17]$_DFFE_PP_  (.D(_00875_),
    .CLK(clknet_leaf_330_clk),
    .Q(\dp.rf.rf[5][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][18]$_DFFE_PP_  (.D(_00876_),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\dp.rf.rf[5][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][19]$_DFFE_PP_  (.D(_00877_),
    .CLK(clknet_leaf_109_clk),
    .Q(\dp.rf.rf[5][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][1]$_DFFE_PP_  (.D(_00878_),
    .CLK(clknet_leaf_502_clk),
    .Q(\dp.rf.rf[5][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][20]$_DFFE_PP_  (.D(_00879_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[5][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][21]$_DFFE_PP_  (.D(_00880_),
    .CLK(clknet_leaf_670_clk),
    .Q(\dp.rf.rf[5][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][22]$_DFFE_PP_  (.D(_00881_),
    .CLK(clknet_leaf_675_clk),
    .Q(\dp.rf.rf[5][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][23]$_DFFE_PP_  (.D(_00882_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\dp.rf.rf[5][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][24]$_DFFE_PP_  (.D(_00883_),
    .CLK(clknet_6_1__leaf_clk),
    .Q(\dp.rf.rf[5][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][25]$_DFFE_PP_  (.D(_00884_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[5][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][26]$_DFFE_PP_  (.D(_00885_),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\dp.rf.rf[5][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][27]$_DFFE_PP_  (.D(_00886_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\dp.rf.rf[5][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][28]$_DFFE_PP_  (.D(_00887_),
    .CLK(clknet_leaf_12_clk),
    .Q(\dp.rf.rf[5][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][29]$_DFFE_PP_  (.D(_00888_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[5][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][2]$_DFFE_PP_  (.D(_00889_),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\dp.rf.rf[5][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][30]$_DFFE_PP_  (.D(_00890_),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\dp.rf.rf[5][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][31]$_DFFE_PP_  (.D(_00891_),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\dp.rf.rf[5][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][3]$_DFFE_PP_  (.D(_00892_),
    .CLK(clknet_leaf_165_clk),
    .Q(\dp.rf.rf[5][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][4]$_DFFE_PP_  (.D(_00893_),
    .CLK(clknet_leaf_626_clk),
    .Q(\dp.rf.rf[5][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][5]$_DFFE_PP_  (.D(_00894_),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\dp.rf.rf[5][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][6]$_DFFE_PP_  (.D(_00895_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[5][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][7]$_DFFE_PP_  (.D(_00896_),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\dp.rf.rf[5][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][8]$_DFFE_PP_  (.D(_00897_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[5][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[5][9]$_DFFE_PP_  (.D(_00898_),
    .CLK(clknet_leaf_639_clk),
    .Q(\dp.rf.rf[5][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][0]$_DFFE_PP_  (.D(_00899_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\dp.rf.rf[6][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][10]$_DFFE_PP_  (.D(_00900_),
    .CLK(clknet_6_62__leaf_clk),
    .Q(\dp.rf.rf[6][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][11]$_DFFE_PP_  (.D(_00901_),
    .CLK(clknet_leaf_248_clk),
    .Q(\dp.rf.rf[6][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][12]$_DFFE_PP_  (.D(_00902_),
    .CLK(clknet_leaf_145_clk),
    .Q(\dp.rf.rf[6][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][13]$_DFFE_PP_  (.D(_00903_),
    .CLK(clknet_leaf_221_clk),
    .Q(\dp.rf.rf[6][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][14]$_DFFE_PP_  (.D(_00904_),
    .CLK(clknet_leaf_232_clk),
    .Q(\dp.rf.rf[6][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][15]$_DFFE_PP_  (.D(_00905_),
    .CLK(clknet_leaf_250_clk),
    .Q(\dp.rf.rf[6][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][16]$_DFFE_PP_  (.D(_00906_),
    .CLK(clknet_leaf_427_clk),
    .Q(\dp.rf.rf[6][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][17]$_DFFE_PP_  (.D(_00907_),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\dp.rf.rf[6][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][18]$_DFFE_PP_  (.D(_00908_),
    .CLK(clknet_leaf_85_clk),
    .Q(\dp.rf.rf[6][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][19]$_DFFE_PP_  (.D(_00909_),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\dp.rf.rf[6][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][1]$_DFFE_PP_  (.D(_00910_),
    .CLK(clknet_leaf_507_clk),
    .Q(\dp.rf.rf[6][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][20]$_DFFE_PP_  (.D(_00911_),
    .CLK(clknet_leaf_448_clk),
    .Q(\dp.rf.rf[6][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][21]$_DFFE_PP_  (.D(_00912_),
    .CLK(clknet_leaf_688_clk),
    .Q(\dp.rf.rf[6][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][22]$_DFFE_PP_  (.D(_00913_),
    .CLK(clknet_leaf_684_clk),
    .Q(\dp.rf.rf[6][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][23]$_DFFE_PP_  (.D(_00914_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[6][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][24]$_DFFE_PP_  (.D(_00915_),
    .CLK(clknet_leaf_679_clk),
    .Q(\dp.rf.rf[6][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][25]$_DFFE_PP_  (.D(_00916_),
    .CLK(clknet_leaf_536_clk),
    .Q(\dp.rf.rf[6][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][26]$_DFFE_PP_  (.D(_00917_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[6][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][27]$_DFFE_PP_  (.D(_00918_),
    .CLK(clknet_leaf_497_clk),
    .Q(\dp.rf.rf[6][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][28]$_DFFE_PP_  (.D(_00919_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[6][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][29]$_DFFE_PP_  (.D(_00920_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\dp.rf.rf[6][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][2]$_DFFE_PP_  (.D(_00921_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[6][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][30]$_DFFE_PP_  (.D(_00922_),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\dp.rf.rf[6][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][31]$_DFFE_PP_  (.D(_00923_),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\dp.rf.rf[6][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][3]$_DFFE_PP_  (.D(_00924_),
    .CLK(clknet_leaf_153_clk),
    .Q(\dp.rf.rf[6][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][4]$_DFFE_PP_  (.D(_00925_),
    .CLK(clknet_leaf_630_clk),
    .Q(\dp.rf.rf[6][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][5]$_DFFE_PP_  (.D(_00926_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\dp.rf.rf[6][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][6]$_DFFE_PP_  (.D(_00927_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[6][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][7]$_DFFE_PP_  (.D(_00928_),
    .CLK(clknet_leaf_81_clk),
    .Q(\dp.rf.rf[6][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][8]$_DFFE_PP_  (.D(_00929_),
    .CLK(clknet_leaf_441_clk),
    .Q(\dp.rf.rf[6][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[6][9]$_DFFE_PP_  (.D(_00930_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\dp.rf.rf[6][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][0]$_DFFE_PP_  (.D(_00931_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\dp.rf.rf[7][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][10]$_DFFE_PP_  (.D(_00932_),
    .CLK(clknet_6_62__leaf_clk),
    .Q(\dp.rf.rf[7][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][11]$_DFFE_PP_  (.D(_00933_),
    .CLK(clknet_leaf_249_clk),
    .Q(\dp.rf.rf[7][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][12]$_DFFE_PP_  (.D(_00934_),
    .CLK(clknet_leaf_145_clk),
    .Q(\dp.rf.rf[7][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][13]$_DFFE_PP_  (.D(_00935_),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\dp.rf.rf[7][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][14]$_DFFE_PP_  (.D(_00936_),
    .CLK(clknet_leaf_232_clk),
    .Q(\dp.rf.rf[7][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][15]$_DFFE_PP_  (.D(_00937_),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\dp.rf.rf[7][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][16]$_DFFE_PP_  (.D(_00938_),
    .CLK(clknet_leaf_427_clk),
    .Q(\dp.rf.rf[7][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][17]$_DFFE_PP_  (.D(_00939_),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\dp.rf.rf[7][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][18]$_DFFE_PP_  (.D(_00940_),
    .CLK(clknet_leaf_81_clk),
    .Q(\dp.rf.rf[7][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][19]$_DFFE_PP_  (.D(_00941_),
    .CLK(clknet_leaf_109_clk),
    .Q(\dp.rf.rf[7][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][1]$_DFFE_PP_  (.D(_00942_),
    .CLK(clknet_leaf_507_clk),
    .Q(\dp.rf.rf[7][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][20]$_DFFE_PP_  (.D(_00943_),
    .CLK(clknet_leaf_448_clk),
    .Q(\dp.rf.rf[7][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][21]$_DFFE_PP_  (.D(_00944_),
    .CLK(clknet_leaf_687_clk),
    .Q(\dp.rf.rf[7][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][22]$_DFFE_PP_  (.D(_00945_),
    .CLK(clknet_leaf_685_clk),
    .Q(\dp.rf.rf[7][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][23]$_DFFE_PP_  (.D(_00946_),
    .CLK(clknet_leaf_484_clk),
    .Q(\dp.rf.rf[7][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][24]$_DFFE_PP_  (.D(_00947_),
    .CLK(clknet_leaf_679_clk),
    .Q(\dp.rf.rf[7][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][25]$_DFFE_PP_  (.D(_00948_),
    .CLK(clknet_leaf_536_clk),
    .Q(\dp.rf.rf[7][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][26]$_DFFE_PP_  (.D(_00949_),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\dp.rf.rf[7][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][27]$_DFFE_PP_  (.D(_00950_),
    .CLK(clknet_leaf_497_clk),
    .Q(\dp.rf.rf[7][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][28]$_DFFE_PP_  (.D(_00951_),
    .CLK(clknet_leaf_3_clk),
    .Q(\dp.rf.rf[7][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][29]$_DFFE_PP_  (.D(_00952_),
    .CLK(clknet_leaf_562_clk),
    .Q(\dp.rf.rf[7][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][2]$_DFFE_PP_  (.D(_00953_),
    .CLK(clknet_leaf_18_clk),
    .Q(\dp.rf.rf[7][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][30]$_DFFE_PP_  (.D(_00954_),
    .CLK(clknet_leaf_581_clk),
    .Q(\dp.rf.rf[7][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][31]$_DFFE_PP_  (.D(_00955_),
    .CLK(clknet_leaf_370_clk),
    .Q(\dp.rf.rf[7][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][3]$_DFFE_PP_  (.D(_00956_),
    .CLK(clknet_leaf_153_clk),
    .Q(\dp.rf.rf[7][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][4]$_DFFE_PP_  (.D(_00957_),
    .CLK(clknet_leaf_630_clk),
    .Q(\dp.rf.rf[7][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][5]$_DFFE_PP_  (.D(_00958_),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\dp.rf.rf[7][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][6]$_DFFE_PP_  (.D(_00959_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[7][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][7]$_DFFE_PP_  (.D(_00960_),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\dp.rf.rf[7][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][8]$_DFFE_PP_  (.D(_00961_),
    .CLK(clknet_leaf_442_clk),
    .Q(\dp.rf.rf[7][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[7][9]$_DFFE_PP_  (.D(_00962_),
    .CLK(clknet_leaf_642_clk),
    .Q(\dp.rf.rf[7][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][0]$_DFFE_PP_  (.D(_00963_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\dp.rf.rf[8][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][10]$_DFFE_PP_  (.D(_00964_),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[8][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][11]$_DFFE_PP_  (.D(_00965_),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\dp.rf.rf[8][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][12]$_DFFE_PP_  (.D(_00966_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\dp.rf.rf[8][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][13]$_DFFE_PP_  (.D(_00967_),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\dp.rf.rf[8][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][14]$_DFFE_PP_  (.D(_00968_),
    .CLK(clknet_leaf_238_clk),
    .Q(\dp.rf.rf[8][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][15]$_DFFE_PP_  (.D(_00969_),
    .CLK(clknet_leaf_276_clk),
    .Q(\dp.rf.rf[8][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][16]$_DFFE_PP_  (.D(_00970_),
    .CLK(clknet_leaf_418_clk),
    .Q(\dp.rf.rf[8][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][17]$_DFFE_PP_  (.D(_00971_),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\dp.rf.rf[8][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][18]$_DFFE_PP_  (.D(_00972_),
    .CLK(clknet_leaf_87_clk),
    .Q(\dp.rf.rf[8][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][19]$_DFFE_PP_  (.D(_00973_),
    .CLK(clknet_leaf_79_clk),
    .Q(\dp.rf.rf[8][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][1]$_DFFE_PP_  (.D(_00974_),
    .CLK(clknet_leaf_496_clk),
    .Q(\dp.rf.rf[8][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][20]$_DFFE_PP_  (.D(_00975_),
    .CLK(clknet_6_21__leaf_clk),
    .Q(\dp.rf.rf[8][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][21]$_DFFE_PP_  (.D(_00976_),
    .CLK(clknet_leaf_687_clk),
    .Q(\dp.rf.rf[8][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][22]$_DFFE_PP_  (.D(_00977_),
    .CLK(clknet_leaf_681_clk),
    .Q(\dp.rf.rf[8][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][23]$_DFFE_PP_  (.D(_00978_),
    .CLK(clknet_leaf_449_clk),
    .Q(\dp.rf.rf[8][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][24]$_DFFE_PP_  (.D(_00979_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\dp.rf.rf[8][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][25]$_DFFE_PP_  (.D(_00980_),
    .CLK(clknet_leaf_469_clk),
    .Q(\dp.rf.rf[8][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][26]$_DFFE_PP_  (.D(_00981_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\dp.rf.rf[8][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][27]$_DFFE_PP_  (.D(_00982_),
    .CLK(clknet_leaf_465_clk),
    .Q(\dp.rf.rf[8][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][28]$_DFFE_PP_  (.D(_00983_),
    .CLK(clknet_leaf_6_clk),
    .Q(\dp.rf.rf[8][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][29]$_DFFE_PP_  (.D(_00984_),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\dp.rf.rf[8][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][2]$_DFFE_PP_  (.D(_00985_),
    .CLK(clknet_leaf_22_clk),
    .Q(\dp.rf.rf[8][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][30]$_DFFE_PP_  (.D(_00986_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\dp.rf.rf[8][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][31]$_DFFE_PP_  (.D(_00987_),
    .CLK(clknet_leaf_432_clk),
    .Q(\dp.rf.rf[8][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][3]$_DFFE_PP_  (.D(_00988_),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\dp.rf.rf[8][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][4]$_DFFE_PP_  (.D(_00989_),
    .CLK(clknet_leaf_509_clk),
    .Q(\dp.rf.rf[8][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][5]$_DFFE_PP_  (.D(_00990_),
    .CLK(clknet_leaf_222_clk),
    .Q(\dp.rf.rf[8][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][6]$_DFFE_PP_  (.D(_00991_),
    .CLK(clknet_leaf_421_clk),
    .Q(\dp.rf.rf[8][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][7]$_DFFE_PP_  (.D(_00992_),
    .CLK(clknet_leaf_76_clk),
    .Q(\dp.rf.rf[8][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][8]$_DFFE_PP_  (.D(_00993_),
    .CLK(clknet_leaf_457_clk),
    .Q(\dp.rf.rf[8][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[8][9]$_DFFE_PP_  (.D(_00994_),
    .CLK(clknet_leaf_631_clk),
    .Q(\dp.rf.rf[8][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][0]$_DFFE_PP_  (.D(_00995_),
    .CLK(clknet_leaf_160_clk),
    .Q(\dp.rf.rf[9][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][10]$_DFFE_PP_  (.D(_00996_),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[9][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][11]$_DFFE_PP_  (.D(_00997_),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\dp.rf.rf[9][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][12]$_DFFE_PP_  (.D(_00998_),
    .CLK(clknet_leaf_125_clk),
    .Q(\dp.rf.rf[9][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][13]$_DFFE_PP_  (.D(_00999_),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\dp.rf.rf[9][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][14]$_DFFE_PP_  (.D(_01000_),
    .CLK(clknet_leaf_238_clk),
    .Q(\dp.rf.rf[9][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][15]$_DFFE_PP_  (.D(_01001_),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\dp.rf.rf[9][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][16]$_DFFE_PP_  (.D(_01002_),
    .CLK(clknet_leaf_418_clk),
    .Q(\dp.rf.rf[9][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][17]$_DFFE_PP_  (.D(_01003_),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\dp.rf.rf[9][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][18]$_DFFE_PP_  (.D(_01004_),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\dp.rf.rf[9][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][19]$_DFFE_PP_  (.D(_01005_),
    .CLK(clknet_leaf_79_clk),
    .Q(\dp.rf.rf[9][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][1]$_DFFE_PP_  (.D(_01006_),
    .CLK(clknet_leaf_496_clk),
    .Q(\dp.rf.rf[9][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][20]$_DFFE_PP_  (.D(_01007_),
    .CLK(clknet_leaf_459_clk),
    .Q(\dp.rf.rf[9][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][21]$_DFFE_PP_  (.D(_01008_),
    .CLK(clknet_leaf_688_clk),
    .Q(\dp.rf.rf[9][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][22]$_DFFE_PP_  (.D(_01009_),
    .CLK(clknet_leaf_681_clk),
    .Q(\dp.rf.rf[9][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][23]$_DFFE_PP_  (.D(_01010_),
    .CLK(clknet_6_21__leaf_clk),
    .Q(\dp.rf.rf[9][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][24]$_DFFE_PP_  (.D(_01011_),
    .CLK(clknet_leaf_688_clk),
    .Q(\dp.rf.rf[9][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][25]$_DFFE_PP_  (.D(_01012_),
    .CLK(clknet_leaf_468_clk),
    .Q(\dp.rf.rf[9][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][26]$_DFFE_PP_  (.D(_01013_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\dp.rf.rf[9][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][27]$_DFFE_PP_  (.D(_01014_),
    .CLK(clknet_leaf_465_clk),
    .Q(\dp.rf.rf[9][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][28]$_DFFE_PP_  (.D(_01015_),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\dp.rf.rf[9][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][29]$_DFFE_PP_  (.D(_01016_),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\dp.rf.rf[9][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][2]$_DFFE_PP_  (.D(_01017_),
    .CLK(clknet_leaf_20_clk),
    .Q(\dp.rf.rf[9][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][30]$_DFFE_PP_  (.D(_01018_),
    .CLK(clknet_leaf_534_clk),
    .Q(\dp.rf.rf[9][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][31]$_DFFE_PP_  (.D(_01019_),
    .CLK(clknet_leaf_432_clk),
    .Q(\dp.rf.rf[9][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][3]$_DFFE_PP_  (.D(_01020_),
    .CLK(clknet_leaf_170_clk),
    .Q(\dp.rf.rf[9][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][4]$_DFFE_PP_  (.D(_01021_),
    .CLK(clknet_leaf_509_clk),
    .Q(\dp.rf.rf[9][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][5]$_DFFE_PP_  (.D(_01022_),
    .CLK(clknet_leaf_131_clk),
    .Q(\dp.rf.rf[9][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][6]$_DFFE_PP_  (.D(_01023_),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\dp.rf.rf[9][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][7]$_DFFE_PP_  (.D(_01024_),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\dp.rf.rf[9][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][8]$_DFFE_PP_  (.D(_01025_),
    .CLK(clknet_leaf_457_clk),
    .Q(\dp.rf.rf[9][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \dp.rf.rf[9][9]$_DFFE_PP_  (.D(_01026_),
    .CLK(clknet_leaf_631_clk),
    .Q(\dp.rf.rf[9][9] ));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_991 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_49__f_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_6_49__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_50__f_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_6_50__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_51__f_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_6_51__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_52__f_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_6_52__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_53__f_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_6_53__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_54__f_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_6_54__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_55__f_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_6_55__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_56__f_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_6_56__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_57__f_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_6_57__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_58__f_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_6_58__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_59__f_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_6_59__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_60__f_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_6_60__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_61__f_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_6_61__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_62__f_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_6_62__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_6_63__f_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_6_63__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload0 (.I(clknet_6_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload1 (.I(clknet_6_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload2 (.I(clknet_6_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload3 (.I(clknet_6_5__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload4 (.I(clknet_6_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload5 (.I(clknet_6_7__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload6 (.I(clknet_6_9__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload7 (.I(clknet_6_10__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload8 (.I(clknet_6_11__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload9 (.I(clknet_6_12__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload10 (.I(clknet_6_14__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload11 (.I(clknet_6_15__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload12 (.I(clknet_6_16__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload13 (.I(clknet_6_18__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload14 (.I(clknet_6_19__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload15 (.I(clknet_6_21__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload16 (.I(clknet_6_22__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload17 (.I(clknet_6_23__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload18 (.I(clknet_6_24__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload19 (.I(clknet_6_26__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload20 (.I(clknet_6_27__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 clkload21 (.I(clknet_6_28__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload22 (.I(clknet_6_30__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload23 (.I(clknet_6_31__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload24 (.I(clknet_6_32__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload25 (.I(clknet_6_33__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload26 (.I(clknet_6_35__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload27 (.I(clknet_6_37__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload28 (.I(clknet_6_38__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload29 (.I(clknet_6_39__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload30 (.I(clknet_6_40__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload31 (.I(clknet_6_41__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload32 (.I(clknet_6_43__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload33 (.I(clknet_6_44__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload34 (.I(clknet_6_45__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload35 (.I(clknet_6_47__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload36 (.I(clknet_6_48__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload37 (.I(clknet_6_49__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload38 (.I(clknet_6_51__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload39 (.I(clknet_6_52__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload40 (.I(clknet_6_54__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload41 (.I(clknet_6_56__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload42 (.I(clknet_6_58__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload43 (.I(clknet_6_59__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload44 (.I(clknet_6_62__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload45 (.I(clknet_6_63__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload46 (.I(clknet_leaf_675_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload47 (.I(clknet_leaf_680_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload48 (.I(clknet_leaf_681_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload49 (.I(clknet_leaf_684_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload50 (.I(clknet_leaf_685_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload51 (.I(clknet_leaf_647_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload52 (.I(clknet_leaf_651_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload53 (.I(clknet_leaf_658_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload54 (.I(clknet_leaf_678_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload55 (.I(clknet_leaf_668_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload56 (.I(clknet_leaf_682_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload57 (.I(clknet_leaf_687_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload58 (.I(clknet_leaf_692_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload59 (.I(clknet_leaf_509_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload60 (.I(clknet_leaf_515_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload61 (.I(clknet_leaf_622_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload62 (.I(clknet_leaf_626_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload63 (.I(clknet_leaf_628_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload64 (.I(clknet_leaf_629_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload65 (.I(clknet_leaf_630_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload66 (.I(clknet_leaf_516_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload67 (.I(clknet_leaf_526_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload68 (.I(clknet_leaf_528_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload69 (.I(clknet_leaf_616_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload70 (.I(clknet_leaf_618_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload71 (.I(clknet_leaf_623_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload72 (.I(clknet_leaf_624_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload73 (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload74 (.I(clknet_leaf_705_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload75 (.I(clknet_leaf_711_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload76 (.I(clknet_leaf_712_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload77 (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload78 (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload79 (.I(clknet_leaf_662_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload80 (.I(clknet_leaf_664_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload81 (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload82 (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload83 (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload84 (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload85 (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload86 (.I(clknet_leaf_591_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload87 (.I(clknet_leaf_592_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload88 (.I(clknet_leaf_595_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload89 (.I(clknet_leaf_597_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload90 (.I(clknet_leaf_486_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload91 (.I(clknet_leaf_488_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload92 (.I(clknet_leaf_494_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload93 (.I(clknet_leaf_496_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload94 (.I(clknet_leaf_481_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload95 (.I(clknet_leaf_370_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload96 (.I(clknet_leaf_557_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload97 (.I(clknet_leaf_569_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload98 (.I(clknet_leaf_423_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload99 (.I(clknet_leaf_425_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload100 (.I(clknet_leaf_452_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload101 (.I(clknet_leaf_456_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload102 (.I(clknet_leaf_457_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload103 (.I(clknet_leaf_458_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload104 (.I(clknet_leaf_408_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload105 (.I(clknet_leaf_418_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload106 (.I(clknet_leaf_419_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload107 (.I(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload108 (.I(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload109 (.I(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload110 (.I(clknet_leaf_228_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload111 (.I(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload112 (.I(clknet_leaf_246_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload113 (.I(clknet_leaf_131_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload114 (.I(clknet_leaf_134_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload115 (.I(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload116 (.I(clknet_leaf_222_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload117 (.I(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload118 (.I(clknet_leaf_220_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload119 (.I(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload120 (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload121 (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload122 (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload123 (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload124 (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload125 (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload126 (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload127 (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload128 (.I(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload129 (.I(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload130 (.I(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload131 (.I(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload132 (.I(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload133 (.I(clknet_leaf_176_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload134 (.I(clknet_leaf_324_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload135 (.I(clknet_leaf_328_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload136 (.I(clknet_leaf_333_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload137 (.I(clknet_leaf_334_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload138 (.I(clknet_leaf_294_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload139 (.I(clknet_leaf_307_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload140 (.I(clknet_leaf_309_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload141 (.I(clknet_leaf_313_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload142 (.I(clknet_leaf_317_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload143 (.I(clknet_leaf_185_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload144 (.I(clknet_leaf_187_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload145 (.I(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload146 (.I(clknet_leaf_250_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload147 (.I(clknet_leaf_251_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload148 (.I(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload149 (.I(clknet_leaf_256_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload150 (.I(clknet_leaf_254_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload151 (.I(clknet_leaf_276_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload152 (.I(clknet_leaf_277_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload153 (.I(clknet_leaf_282_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload154 (.I(clknet_leaf_242_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload155 (.I(clknet_leaf_249_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload156 (.I(clknet_leaf_270_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload157 (.I(clknet_leaf_271_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 split1 (.I(net166),
    .Z(net165));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2 (.I(_01126_),
    .Z(net166));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer3 (.I(_01126_),
    .Z(net167));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer4 (.I(_01126_),
    .Z(net168));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_109_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_110_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_113_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_114_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_117_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_126_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_131_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_132_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_133_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_138_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1486 ();
endmodule
