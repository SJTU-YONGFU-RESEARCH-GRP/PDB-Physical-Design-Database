module simple_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \bit_count[3] ;
 wire \rx_shift_reg[0] ;
 wire \rx_shift_reg[1] ;
 wire \rx_shift_reg[2] ;
 wire \rx_shift_reg[3] ;
 wire \rx_shift_reg[4] ;
 wire \rx_shift_reg[5] ;
 wire \rx_shift_reg[6] ;
 wire \rx_shift_reg[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \tx_shift_reg[0] ;
 wire \tx_shift_reg[1] ;
 wire \tx_shift_reg[2] ;
 wire \tx_shift_reg[3] ;
 wire \tx_shift_reg[4] ;
 wire \tx_shift_reg[5] ;
 wire \tx_shift_reg[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 BUF_X2 _217_ (.A(\bit_count[3] ),
    .Z(_037_));
 INV_X1 _218_ (.A(_037_),
    .ZN(_038_));
 BUF_X4 _219_ (.A(\bit_count[2] ),
    .Z(_039_));
 NAND3_X2 _220_ (.A1(_038_),
    .A2(_039_),
    .A3(_198_),
    .ZN(_204_));
 INV_X1 _221_ (.A(_204_),
    .ZN(_207_));
 BUF_X1 _222_ (.A(rst_n),
    .Z(_040_));
 INV_X2 _223_ (.A(_040_),
    .ZN(_041_));
 CLKBUF_X3 _224_ (.A(_041_),
    .Z(_042_));
 CLKBUF_X3 _225_ (.A(\state[2] ),
    .Z(_043_));
 CLKBUF_X3 _226_ (.A(_043_),
    .Z(_044_));
 NAND2_X1 _227_ (.A1(_038_),
    .A2(_004_),
    .ZN(_045_));
 CLKBUF_X2 _228_ (.A(net20),
    .Z(_046_));
 INV_X1 _229_ (.A(_046_),
    .ZN(_047_));
 AND2_X1 _230_ (.A1(_047_),
    .A2(_205_),
    .ZN(_048_));
 OAI21_X1 _231_ (.A(_044_),
    .B1(_045_),
    .B2(_048_),
    .ZN(_049_));
 BUF_X4 _232_ (.A(\state[0] ),
    .Z(_050_));
 NAND2_X1 _233_ (.A1(net10),
    .A2(_050_),
    .ZN(_051_));
 AOI21_X1 _234_ (.A(_042_),
    .B1(_049_),
    .B2(_051_),
    .ZN(_002_));
 CLKBUF_X3 _235_ (.A(_040_),
    .Z(_052_));
 BUF_X1 _236_ (.A(\state[1] ),
    .Z(_053_));
 INV_X2 _237_ (.A(_053_),
    .ZN(_054_));
 INV_X1 _238_ (.A(_050_),
    .ZN(_055_));
 OR2_X1 _239_ (.A1(net10),
    .A2(_055_),
    .ZN(_056_));
 NAND3_X1 _240_ (.A1(_052_),
    .A2(_054_),
    .A3(_056_),
    .ZN(_001_));
 AND4_X1 _241_ (.A1(_047_),
    .A2(_052_),
    .A3(_044_),
    .A4(_208_),
    .ZN(_000_));
 NAND3_X1 _242_ (.A1(_039_),
    .A2(\bit_count[0] ),
    .A3(\bit_count[1] ),
    .ZN(_201_));
 OR2_X1 _243_ (.A1(_037_),
    .A2(_201_),
    .ZN(_214_));
 INV_X1 _244_ (.A(\bit_count[0] ),
    .ZN(_057_));
 NAND2_X1 _245_ (.A1(_044_),
    .A2(_057_),
    .ZN(_058_));
 MUX2_X2 _246_ (.A(\state[2] ),
    .B(net10),
    .S(_050_),
    .Z(_059_));
 INV_X1 _247_ (.A(_059_),
    .ZN(_060_));
 OAI21_X1 _248_ (.A(_200_),
    .B1(_047_),
    .B2(_037_),
    .ZN(_061_));
 AOI21_X2 _249_ (.A(_060_),
    .B1(_061_),
    .B2(_044_),
    .ZN(_062_));
 MUX2_X1 _250_ (.A(_057_),
    .B(_058_),
    .S(_062_),
    .Z(_063_));
 NOR2_X1 _251_ (.A1(_042_),
    .A2(_063_),
    .ZN(_005_));
 BUF_X2 _252_ (.A(_052_),
    .Z(_064_));
 INV_X2 _253_ (.A(\state[2] ),
    .ZN(_065_));
 BUF_X2 _254_ (.A(_199_),
    .Z(_066_));
 INV_X1 _255_ (.A(_066_),
    .ZN(_067_));
 NOR2_X1 _256_ (.A1(_065_),
    .A2(_067_),
    .ZN(_068_));
 MUX2_X1 _257_ (.A(\bit_count[1] ),
    .B(_068_),
    .S(_062_),
    .Z(_069_));
 AND2_X1 _258_ (.A1(_064_),
    .A2(_069_),
    .ZN(_006_));
 NAND3_X1 _259_ (.A1(_039_),
    .A2(_052_),
    .A3(_060_),
    .ZN(_070_));
 NAND2_X1 _260_ (.A1(_052_),
    .A2(_044_),
    .ZN(_071_));
 INV_X1 _261_ (.A(_039_),
    .ZN(_072_));
 NAND2_X1 _262_ (.A1(_072_),
    .A2(_056_),
    .ZN(_073_));
 INV_X1 _263_ (.A(_198_),
    .ZN(_074_));
 NOR2_X1 _264_ (.A1(_074_),
    .A2(_061_),
    .ZN(_075_));
 MUX2_X1 _265_ (.A(_072_),
    .B(_073_),
    .S(_075_),
    .Z(_076_));
 OAI21_X1 _266_ (.A(_070_),
    .B1(_071_),
    .B2(_076_),
    .ZN(_007_));
 NOR2_X1 _267_ (.A1(_065_),
    .A2(_200_),
    .ZN(_077_));
 NOR2_X1 _268_ (.A1(_060_),
    .A2(_077_),
    .ZN(_078_));
 NAND2_X1 _269_ (.A1(_043_),
    .A2(_203_),
    .ZN(_079_));
 NAND2_X1 _270_ (.A1(_047_),
    .A2(_078_),
    .ZN(_080_));
 AOI221_X1 _271_ (.A(_041_),
    .B1(_078_),
    .B2(_079_),
    .C1(_080_),
    .C2(_038_),
    .ZN(_008_));
 CLKBUF_X3 _272_ (.A(_053_),
    .Z(_081_));
 NAND2_X1 _273_ (.A1(_081_),
    .A2(\rx_shift_reg[0] ),
    .ZN(_082_));
 NAND2_X1 _274_ (.A1(_054_),
    .A2(net11),
    .ZN(_083_));
 AOI21_X1 _275_ (.A(_042_),
    .B1(_082_),
    .B2(_083_),
    .ZN(_009_));
 NAND2_X1 _276_ (.A1(_081_),
    .A2(\rx_shift_reg[1] ),
    .ZN(_084_));
 NAND2_X1 _277_ (.A1(_054_),
    .A2(net12),
    .ZN(_085_));
 AOI21_X1 _278_ (.A(_042_),
    .B1(_084_),
    .B2(_085_),
    .ZN(_010_));
 NAND2_X1 _279_ (.A1(_081_),
    .A2(\rx_shift_reg[2] ),
    .ZN(_086_));
 NAND2_X1 _280_ (.A1(_054_),
    .A2(net13),
    .ZN(_087_));
 AOI21_X1 _281_ (.A(_042_),
    .B1(_086_),
    .B2(_087_),
    .ZN(_011_));
 NAND2_X1 _282_ (.A1(_081_),
    .A2(\rx_shift_reg[3] ),
    .ZN(_088_));
 NAND2_X1 _283_ (.A1(_054_),
    .A2(net14),
    .ZN(_089_));
 AOI21_X1 _284_ (.A(_042_),
    .B1(_088_),
    .B2(_089_),
    .ZN(_012_));
 NAND2_X1 _285_ (.A1(_081_),
    .A2(\rx_shift_reg[4] ),
    .ZN(_090_));
 NAND2_X1 _286_ (.A1(_054_),
    .A2(net15),
    .ZN(_091_));
 AOI21_X1 _287_ (.A(_042_),
    .B1(_090_),
    .B2(_091_),
    .ZN(_013_));
 NAND2_X1 _288_ (.A1(_081_),
    .A2(\rx_shift_reg[5] ),
    .ZN(_092_));
 NAND2_X1 _289_ (.A1(_054_),
    .A2(net16),
    .ZN(_093_));
 AOI21_X1 _290_ (.A(_042_),
    .B1(_092_),
    .B2(_093_),
    .ZN(_014_));
 NAND2_X1 _291_ (.A1(_081_),
    .A2(\rx_shift_reg[6] ),
    .ZN(_094_));
 NAND2_X1 _292_ (.A1(_054_),
    .A2(net17),
    .ZN(_095_));
 AOI21_X1 _293_ (.A(_042_),
    .B1(_094_),
    .B2(_095_),
    .ZN(_015_));
 NAND2_X1 _294_ (.A1(_081_),
    .A2(\rx_shift_reg[7] ),
    .ZN(_096_));
 NAND2_X1 _295_ (.A1(_054_),
    .A2(net18),
    .ZN(_097_));
 AOI21_X1 _296_ (.A(_041_),
    .B1(_096_),
    .B2(_097_),
    .ZN(_016_));
 AND2_X1 _297_ (.A1(_040_),
    .A2(net1),
    .ZN(_098_));
 AND2_X1 _298_ (.A1(_052_),
    .A2(\rx_shift_reg[0] ),
    .ZN(_099_));
 INV_X1 _299_ (.A(_206_),
    .ZN(_100_));
 INV_X1 _300_ (.A(_216_),
    .ZN(_101_));
 AND4_X2 _301_ (.A1(_100_),
    .A2(_101_),
    .A3(_202_),
    .A4(_215_),
    .ZN(_102_));
 NOR4_X1 _302_ (.A1(_100_),
    .A2(_101_),
    .A3(_202_),
    .A4(_215_),
    .ZN(_103_));
 OR2_X1 _303_ (.A1(_102_),
    .A2(_103_),
    .ZN(_104_));
 NOR3_X1 _304_ (.A1(_100_),
    .A2(_066_),
    .A3(_079_),
    .ZN(_105_));
 OR2_X1 _305_ (.A1(_037_),
    .A2(_046_),
    .ZN(_106_));
 XOR2_X2 _306_ (.A(_039_),
    .B(_198_),
    .Z(_107_));
 NOR2_X1 _307_ (.A1(_106_),
    .A2(_107_),
    .ZN(_108_));
 NOR3_X2 _308_ (.A1(_212_),
    .A2(_210_),
    .A3(_003_),
    .ZN(_109_));
 NAND4_X1 _309_ (.A1(_104_),
    .A2(_105_),
    .A3(_108_),
    .A4(_109_),
    .ZN(_110_));
 MUX2_X1 _310_ (.A(_098_),
    .B(_099_),
    .S(_110_),
    .Z(_017_));
 NAND2_X1 _311_ (.A1(_052_),
    .A2(\rx_shift_reg[1] ),
    .ZN(_111_));
 INV_X1 _312_ (.A(_203_),
    .ZN(_112_));
 NOR2_X1 _313_ (.A1(_037_),
    .A2(_046_),
    .ZN(_113_));
 AND4_X1 _314_ (.A1(_043_),
    .A2(_112_),
    .A3(_113_),
    .A4(_107_),
    .ZN(_114_));
 NAND2_X1 _315_ (.A1(_066_),
    .A2(_114_),
    .ZN(_115_));
 NOR3_X1 _316_ (.A1(_037_),
    .A2(\bit_count[0] ),
    .A3(_115_),
    .ZN(_116_));
 NAND2_X1 _317_ (.A1(_057_),
    .A2(_098_),
    .ZN(_117_));
 NOR3_X1 _318_ (.A1(_212_),
    .A2(_210_),
    .A3(_117_),
    .ZN(_118_));
 NAND2_X1 _319_ (.A1(_102_),
    .A2(_118_),
    .ZN(_119_));
 OAI22_X1 _320_ (.A1(_111_),
    .A2(_116_),
    .B1(_119_),
    .B2(_115_),
    .ZN(_018_));
 AND2_X1 _321_ (.A1(_052_),
    .A2(\rx_shift_reg[2] ),
    .ZN(_120_));
 NAND4_X1 _322_ (.A1(_066_),
    .A2(_102_),
    .A3(_109_),
    .A4(_114_),
    .ZN(_121_));
 MUX2_X1 _323_ (.A(_098_),
    .B(_120_),
    .S(_121_),
    .Z(_019_));
 NAND2_X1 _324_ (.A1(_067_),
    .A2(_114_),
    .ZN(_122_));
 NOR3_X1 _325_ (.A1(_037_),
    .A2(\bit_count[0] ),
    .A3(_122_),
    .ZN(_123_));
 NAND2_X1 _326_ (.A1(_052_),
    .A2(\rx_shift_reg[3] ),
    .ZN(_124_));
 OAI22_X1 _327_ (.A1(_119_),
    .A2(_122_),
    .B1(_123_),
    .B2(_124_),
    .ZN(_020_));
 AND2_X1 _328_ (.A1(_040_),
    .A2(\rx_shift_reg[4] ),
    .ZN(_125_));
 NAND4_X1 _329_ (.A1(_067_),
    .A2(_102_),
    .A3(_109_),
    .A4(_114_),
    .ZN(_126_));
 MUX2_X1 _330_ (.A(_098_),
    .B(_125_),
    .S(_126_),
    .Z(_021_));
 NOR4_X4 _331_ (.A1(_065_),
    .A2(_203_),
    .A3(_106_),
    .A4(_107_),
    .ZN(_127_));
 NAND3_X1 _332_ (.A1(_057_),
    .A2(_066_),
    .A3(_127_),
    .ZN(_128_));
 NAND3_X1 _333_ (.A1(_064_),
    .A2(\rx_shift_reg[5] ),
    .A3(_128_),
    .ZN(_129_));
 NAND3_X1 _334_ (.A1(_102_),
    .A2(_118_),
    .A3(_127_),
    .ZN(_130_));
 OAI21_X1 _335_ (.A(_129_),
    .B1(_130_),
    .B2(_067_),
    .ZN(_022_));
 AND2_X1 _336_ (.A1(_040_),
    .A2(\rx_shift_reg[6] ),
    .ZN(_131_));
 NAND4_X1 _337_ (.A1(_066_),
    .A2(_102_),
    .A3(_109_),
    .A4(_127_),
    .ZN(_132_));
 MUX2_X1 _338_ (.A(_098_),
    .B(_131_),
    .S(_132_),
    .Z(_023_));
 NAND3_X1 _339_ (.A1(_057_),
    .A2(_067_),
    .A3(_127_),
    .ZN(_133_));
 NAND3_X1 _340_ (.A1(_064_),
    .A2(\rx_shift_reg[7] ),
    .A3(_133_),
    .ZN(_134_));
 OAI21_X1 _341_ (.A(_134_),
    .B1(_130_),
    .B2(_066_),
    .ZN(_024_));
 AOI21_X1 _342_ (.A(_081_),
    .B1(net19),
    .B2(_055_),
    .ZN(_135_));
 NOR2_X1 _343_ (.A1(_042_),
    .A2(_135_),
    .ZN(_025_));
 NOR2_X1 _344_ (.A1(_050_),
    .A2(_081_),
    .ZN(_136_));
 NAND4_X1 _345_ (.A1(_044_),
    .A2(_004_),
    .A3(_200_),
    .A4(_136_),
    .ZN(_137_));
 NOR3_X1 _346_ (.A1(_044_),
    .A2(_050_),
    .A3(_053_),
    .ZN(_138_));
 OAI21_X1 _347_ (.A(_046_),
    .B1(_077_),
    .B2(_138_),
    .ZN(_139_));
 AOI21_X1 _348_ (.A(_041_),
    .B1(_137_),
    .B2(_139_),
    .ZN(_026_));
 AND2_X1 _349_ (.A1(_055_),
    .A2(net21),
    .ZN(_140_));
 OR2_X1 _350_ (.A1(_001_),
    .A2(_140_),
    .ZN(_027_));
 INV_X1 _351_ (.A(_200_),
    .ZN(_141_));
 OAI21_X2 _352_ (.A(_043_),
    .B1(_141_),
    .B2(_113_),
    .ZN(_142_));
 NAND2_X4 _353_ (.A1(_059_),
    .A2(_142_),
    .ZN(_143_));
 NOR2_X1 _354_ (.A1(_044_),
    .A2(net9),
    .ZN(_144_));
 AOI21_X1 _355_ (.A(\tx_shift_reg[6] ),
    .B1(_208_),
    .B2(_046_),
    .ZN(_145_));
 AOI21_X1 _356_ (.A(_144_),
    .B1(_145_),
    .B2(_044_),
    .ZN(_146_));
 OAI21_X1 _357_ (.A(_052_),
    .B1(_143_),
    .B2(_146_),
    .ZN(_147_));
 NAND3_X1 _358_ (.A1(_046_),
    .A2(_044_),
    .A3(_208_),
    .ZN(_148_));
 NAND3_X1 _359_ (.A1(_059_),
    .A2(_142_),
    .A3(_148_),
    .ZN(_149_));
 INV_X1 _360_ (.A(net22),
    .ZN(_150_));
 AOI21_X1 _361_ (.A(_147_),
    .B1(_149_),
    .B2(_150_),
    .ZN(_028_));
 NAND2_X1 _362_ (.A1(_055_),
    .A2(net23),
    .ZN(_151_));
 NAND3_X1 _363_ (.A1(_064_),
    .A2(_056_),
    .A3(_151_),
    .ZN(_029_));
 NAND2_X1 _364_ (.A1(\tx_shift_reg[0] ),
    .A2(_143_),
    .ZN(_152_));
 NAND3_X1 _365_ (.A1(_065_),
    .A2(net2),
    .A3(_059_),
    .ZN(_153_));
 AOI21_X1 _366_ (.A(_041_),
    .B1(_152_),
    .B2(_153_),
    .ZN(_030_));
 MUX2_X1 _367_ (.A(net3),
    .B(\tx_shift_reg[0] ),
    .S(_043_),
    .Z(_154_));
 MUX2_X1 _368_ (.A(_154_),
    .B(\tx_shift_reg[1] ),
    .S(_143_),
    .Z(_155_));
 AND2_X1 _369_ (.A1(_064_),
    .A2(_155_),
    .ZN(_031_));
 MUX2_X1 _370_ (.A(net4),
    .B(\tx_shift_reg[1] ),
    .S(_043_),
    .Z(_156_));
 MUX2_X1 _371_ (.A(_156_),
    .B(\tx_shift_reg[2] ),
    .S(_143_),
    .Z(_157_));
 AND2_X1 _372_ (.A1(_064_),
    .A2(_157_),
    .ZN(_032_));
 MUX2_X1 _373_ (.A(net5),
    .B(\tx_shift_reg[2] ),
    .S(_043_),
    .Z(_158_));
 MUX2_X1 _374_ (.A(_158_),
    .B(\tx_shift_reg[3] ),
    .S(_143_),
    .Z(_159_));
 AND2_X1 _375_ (.A1(_064_),
    .A2(_159_),
    .ZN(_033_));
 MUX2_X1 _376_ (.A(net6),
    .B(\tx_shift_reg[3] ),
    .S(_043_),
    .Z(_160_));
 MUX2_X1 _377_ (.A(_160_),
    .B(\tx_shift_reg[4] ),
    .S(_143_),
    .Z(_161_));
 AND2_X1 _378_ (.A1(_064_),
    .A2(_161_),
    .ZN(_034_));
 MUX2_X1 _379_ (.A(net7),
    .B(\tx_shift_reg[4] ),
    .S(_043_),
    .Z(_162_));
 MUX2_X1 _380_ (.A(_162_),
    .B(\tx_shift_reg[5] ),
    .S(_143_),
    .Z(_163_));
 AND2_X1 _381_ (.A1(_064_),
    .A2(_163_),
    .ZN(_035_));
 MUX2_X1 _382_ (.A(net8),
    .B(\tx_shift_reg[5] ),
    .S(_043_),
    .Z(_164_));
 MUX2_X1 _383_ (.A(_164_),
    .B(\tx_shift_reg[6] ),
    .S(_143_),
    .Z(_165_));
 AND2_X1 _384_ (.A1(_064_),
    .A2(_165_),
    .ZN(_036_));
 HA_X1 _385_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_198_),
    .S(_199_));
 HA_X1 _386_ (.A(_200_),
    .B(_201_),
    .CO(_202_),
    .S(_203_));
 HA_X1 _387_ (.A(_200_),
    .B(_204_),
    .CO(_205_),
    .S(_206_));
 HA_X1 _388_ (.A(_200_),
    .B(_207_),
    .CO(_208_),
    .S(_209_));
 HA_X1 _389_ (.A(\bit_count[3] ),
    .B(_204_),
    .CO(_210_),
    .S(_211_));
 HA_X1 _390_ (.A(\bit_count[3] ),
    .B(_207_),
    .CO(_212_),
    .S(_213_));
 HA_X1 _391_ (.A(_200_),
    .B(_214_),
    .CO(_215_),
    .S(_216_));
 DFF_X2 \bit_count[0]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\bit_count[0] ),
    .QN(_003_));
 DFF_X1 \bit_count[1]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\bit_count[1] ),
    .QN(_194_));
 DFF_X1 \bit_count[2]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\bit_count[2] ),
    .QN(_193_));
 DFF_X2 \bit_count[3]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\bit_count[3] ),
    .QN(_200_));
 DFF_X1 \rx_data[0]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net11),
    .QN(_192_));
 DFF_X1 \rx_data[1]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net12),
    .QN(_191_));
 DFF_X1 \rx_data[2]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net13),
    .QN(_190_));
 DFF_X1 \rx_data[3]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net14),
    .QN(_189_));
 DFF_X1 \rx_data[4]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_188_));
 DFF_X1 \rx_data[5]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net16),
    .QN(_187_));
 DFF_X1 \rx_data[6]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net17),
    .QN(_186_));
 DFF_X1 \rx_data[7]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net18),
    .QN(_185_));
 DFF_X1 \rx_shift_reg[0]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[0] ),
    .QN(_184_));
 DFF_X1 \rx_shift_reg[1]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[1] ),
    .QN(_183_));
 DFF_X1 \rx_shift_reg[2]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[2] ),
    .QN(_182_));
 DFF_X1 \rx_shift_reg[3]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[3] ),
    .QN(_181_));
 DFF_X1 \rx_shift_reg[4]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[4] ),
    .QN(_180_));
 DFF_X1 \rx_shift_reg[5]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[5] ),
    .QN(_179_));
 DFF_X1 \rx_shift_reg[6]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[6] ),
    .QN(_178_));
 DFF_X1 \rx_shift_reg[7]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[7] ),
    .QN(_177_));
 DFF_X1 \rx_valid$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net19),
    .QN(_176_));
 DFF_X1 \spi_clk$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net20),
    .QN(_004_));
 DFF_X1 \spi_cs_n$_SDFFE_PN1P_  (.D(_027_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net21),
    .QN(_175_));
 DFF_X1 \spi_mosi$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net22),
    .QN(_195_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[0] ),
    .QN(_196_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[1] ),
    .QN(_197_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[2] ),
    .QN(_174_));
 DFF_X1 \tx_ready$_SDFFE_PN1P_  (.D(_029_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net23),
    .QN(_173_));
 DFF_X1 \tx_shift_reg[0]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[0] ),
    .QN(_172_));
 DFF_X1 \tx_shift_reg[1]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[1] ),
    .QN(_171_));
 DFF_X1 \tx_shift_reg[2]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[2] ),
    .QN(_170_));
 DFF_X1 \tx_shift_reg[3]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[3] ),
    .QN(_169_));
 DFF_X1 \tx_shift_reg[4]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\tx_shift_reg[4] ),
    .QN(_168_));
 DFF_X1 \tx_shift_reg[5]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[5] ),
    .QN(_167_));
 DFF_X1 \tx_shift_reg[6]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[6] ),
    .QN(_166_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_67 ();
 BUF_X1 input1 (.A(spi_miso),
    .Z(net1));
 BUF_X1 input2 (.A(tx_data[0]),
    .Z(net2));
 BUF_X1 input3 (.A(tx_data[1]),
    .Z(net3));
 BUF_X1 input4 (.A(tx_data[2]),
    .Z(net4));
 BUF_X1 input5 (.A(tx_data[3]),
    .Z(net5));
 BUF_X1 input6 (.A(tx_data[4]),
    .Z(net6));
 BUF_X1 input7 (.A(tx_data[5]),
    .Z(net7));
 BUF_X1 input8 (.A(tx_data[6]),
    .Z(net8));
 BUF_X1 input9 (.A(tx_data[7]),
    .Z(net9));
 BUF_X1 input10 (.A(tx_valid),
    .Z(net10));
 BUF_X1 output11 (.A(net11),
    .Z(rx_data[0]));
 BUF_X1 output12 (.A(net12),
    .Z(rx_data[1]));
 BUF_X1 output13 (.A(net13),
    .Z(rx_data[2]));
 BUF_X1 output14 (.A(net14),
    .Z(rx_data[3]));
 BUF_X1 output15 (.A(net15),
    .Z(rx_data[4]));
 BUF_X1 output16 (.A(net16),
    .Z(rx_data[5]));
 BUF_X1 output17 (.A(net17),
    .Z(rx_data[6]));
 BUF_X1 output18 (.A(net18),
    .Z(rx_data[7]));
 BUF_X1 output19 (.A(net19),
    .Z(rx_valid));
 BUF_X1 output20 (.A(net20),
    .Z(spi_clk));
 BUF_X1 output21 (.A(net21),
    .Z(spi_cs_n));
 BUF_X1 output22 (.A(net22),
    .Z(spi_mosi));
 BUF_X1 output23 (.A(net23),
    .Z(tx_ready));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_2__leaf_clk));
 CLKBUF_X1 clkload1 (.A(clknet_2_3__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X4 FILLER_0_65 ();
 FILLCELL_X2 FILLER_0_69 ();
 FILLCELL_X4 FILLER_0_74 ();
 FILLCELL_X2 FILLER_0_78 ();
 FILLCELL_X16 FILLER_0_83 ();
 FILLCELL_X4 FILLER_0_99 ();
 FILLCELL_X2 FILLER_0_103 ();
 FILLCELL_X1 FILLER_0_105 ();
 FILLCELL_X16 FILLER_0_109 ();
 FILLCELL_X2 FILLER_0_125 ();
 FILLCELL_X8 FILLER_0_133 ();
 FILLCELL_X32 FILLER_0_144 ();
 FILLCELL_X32 FILLER_0_176 ();
 FILLCELL_X32 FILLER_0_208 ();
 FILLCELL_X16 FILLER_0_240 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_88 ();
 FILLCELL_X4 FILLER_1_99 ();
 FILLCELL_X2 FILLER_1_103 ();
 FILLCELL_X1 FILLER_1_105 ();
 FILLCELL_X2 FILLER_1_113 ();
 FILLCELL_X1 FILLER_1_115 ();
 FILLCELL_X4 FILLER_1_123 ();
 FILLCELL_X2 FILLER_1_127 ();
 FILLCELL_X1 FILLER_1_129 ();
 FILLCELL_X2 FILLER_1_137 ();
 FILLCELL_X1 FILLER_1_139 ();
 FILLCELL_X32 FILLER_1_147 ();
 FILLCELL_X32 FILLER_1_179 ();
 FILLCELL_X32 FILLER_1_211 ();
 FILLCELL_X8 FILLER_1_243 ();
 FILLCELL_X4 FILLER_1_251 ();
 FILLCELL_X1 FILLER_1_255 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X2 FILLER_2_65 ();
 FILLCELL_X1 FILLER_2_67 ();
 FILLCELL_X1 FILLER_2_72 ();
 FILLCELL_X8 FILLER_2_87 ();
 FILLCELL_X8 FILLER_2_99 ();
 FILLCELL_X2 FILLER_2_107 ();
 FILLCELL_X1 FILLER_2_109 ();
 FILLCELL_X4 FILLER_2_131 ();
 FILLCELL_X1 FILLER_2_135 ();
 FILLCELL_X32 FILLER_2_147 ();
 FILLCELL_X32 FILLER_2_179 ();
 FILLCELL_X32 FILLER_2_211 ();
 FILLCELL_X8 FILLER_2_243 ();
 FILLCELL_X4 FILLER_2_251 ();
 FILLCELL_X1 FILLER_2_255 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X1 FILLER_3_65 ();
 FILLCELL_X8 FILLER_3_83 ();
 FILLCELL_X32 FILLER_3_108 ();
 FILLCELL_X1 FILLER_3_140 ();
 FILLCELL_X32 FILLER_3_158 ();
 FILLCELL_X32 FILLER_3_190 ();
 FILLCELL_X32 FILLER_3_222 ();
 FILLCELL_X2 FILLER_3_254 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X16 FILLER_4_225 ();
 FILLCELL_X8 FILLER_4_241 ();
 FILLCELL_X4 FILLER_4_249 ();
 FILLCELL_X2 FILLER_4_253 ();
 FILLCELL_X1 FILLER_4_255 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X16 FILLER_5_97 ();
 FILLCELL_X8 FILLER_5_113 ();
 FILLCELL_X4 FILLER_5_121 ();
 FILLCELL_X2 FILLER_5_125 ();
 FILLCELL_X32 FILLER_5_141 ();
 FILLCELL_X32 FILLER_5_173 ();
 FILLCELL_X32 FILLER_5_205 ();
 FILLCELL_X16 FILLER_5_237 ();
 FILLCELL_X2 FILLER_5_253 ();
 FILLCELL_X1 FILLER_5_255 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X4 FILLER_6_97 ();
 FILLCELL_X2 FILLER_6_101 ();
 FILLCELL_X8 FILLER_6_114 ();
 FILLCELL_X32 FILLER_6_143 ();
 FILLCELL_X32 FILLER_6_175 ();
 FILLCELL_X32 FILLER_6_207 ();
 FILLCELL_X16 FILLER_6_239 ();
 FILLCELL_X1 FILLER_6_255 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X8 FILLER_7_81 ();
 FILLCELL_X4 FILLER_7_89 ();
 FILLCELL_X2 FILLER_7_93 ();
 FILLCELL_X1 FILLER_7_95 ();
 FILLCELL_X32 FILLER_7_113 ();
 FILLCELL_X32 FILLER_7_145 ();
 FILLCELL_X32 FILLER_7_177 ();
 FILLCELL_X32 FILLER_7_209 ();
 FILLCELL_X8 FILLER_7_241 ();
 FILLCELL_X4 FILLER_7_249 ();
 FILLCELL_X2 FILLER_7_253 ();
 FILLCELL_X1 FILLER_7_255 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X16 FILLER_8_225 ();
 FILLCELL_X8 FILLER_8_241 ();
 FILLCELL_X4 FILLER_8_249 ();
 FILLCELL_X2 FILLER_8_253 ();
 FILLCELL_X1 FILLER_8_255 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X16 FILLER_9_225 ();
 FILLCELL_X8 FILLER_9_241 ();
 FILLCELL_X4 FILLER_9_249 ();
 FILLCELL_X2 FILLER_9_253 ();
 FILLCELL_X1 FILLER_9_255 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X16 FILLER_10_33 ();
 FILLCELL_X8 FILLER_10_49 ();
 FILLCELL_X4 FILLER_10_57 ();
 FILLCELL_X32 FILLER_10_81 ();
 FILLCELL_X32 FILLER_10_113 ();
 FILLCELL_X32 FILLER_10_145 ();
 FILLCELL_X32 FILLER_10_177 ();
 FILLCELL_X32 FILLER_10_209 ();
 FILLCELL_X8 FILLER_10_241 ();
 FILLCELL_X4 FILLER_10_249 ();
 FILLCELL_X2 FILLER_10_253 ();
 FILLCELL_X1 FILLER_10_255 ();
 FILLCELL_X16 FILLER_11_1 ();
 FILLCELL_X8 FILLER_11_17 ();
 FILLCELL_X1 FILLER_11_25 ();
 FILLCELL_X32 FILLER_11_29 ();
 FILLCELL_X16 FILLER_11_61 ();
 FILLCELL_X32 FILLER_11_84 ();
 FILLCELL_X8 FILLER_11_116 ();
 FILLCELL_X4 FILLER_11_124 ();
 FILLCELL_X1 FILLER_11_128 ();
 FILLCELL_X32 FILLER_11_133 ();
 FILLCELL_X32 FILLER_11_165 ();
 FILLCELL_X32 FILLER_11_197 ();
 FILLCELL_X16 FILLER_11_229 ();
 FILLCELL_X8 FILLER_11_245 ();
 FILLCELL_X2 FILLER_11_253 ();
 FILLCELL_X1 FILLER_11_255 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X2 FILLER_12_13 ();
 FILLCELL_X1 FILLER_12_15 ();
 FILLCELL_X8 FILLER_12_19 ();
 FILLCELL_X1 FILLER_12_27 ();
 FILLCELL_X16 FILLER_12_31 ();
 FILLCELL_X2 FILLER_12_66 ();
 FILLCELL_X1 FILLER_12_72 ();
 FILLCELL_X1 FILLER_12_102 ();
 FILLCELL_X8 FILLER_12_112 ();
 FILLCELL_X4 FILLER_12_120 ();
 FILLCELL_X1 FILLER_12_124 ();
 FILLCELL_X8 FILLER_12_142 ();
 FILLCELL_X32 FILLER_12_154 ();
 FILLCELL_X32 FILLER_12_186 ();
 FILLCELL_X32 FILLER_12_218 ();
 FILLCELL_X4 FILLER_12_250 ();
 FILLCELL_X2 FILLER_12_254 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X8 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_105 ();
 FILLCELL_X1 FILLER_13_109 ();
 FILLCELL_X8 FILLER_13_115 ();
 FILLCELL_X32 FILLER_13_130 ();
 FILLCELL_X32 FILLER_13_162 ();
 FILLCELL_X32 FILLER_13_194 ();
 FILLCELL_X16 FILLER_13_226 ();
 FILLCELL_X8 FILLER_13_242 ();
 FILLCELL_X4 FILLER_13_250 ();
 FILLCELL_X2 FILLER_13_254 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X4 FILLER_14_65 ();
 FILLCELL_X1 FILLER_14_96 ();
 FILLCELL_X4 FILLER_14_99 ();
 FILLCELL_X1 FILLER_14_109 ();
 FILLCELL_X4 FILLER_14_115 ();
 FILLCELL_X1 FILLER_14_119 ();
 FILLCELL_X2 FILLER_14_130 ();
 FILLCELL_X1 FILLER_14_132 ();
 FILLCELL_X4 FILLER_14_136 ();
 FILLCELL_X2 FILLER_14_140 ();
 FILLCELL_X1 FILLER_14_142 ();
 FILLCELL_X1 FILLER_14_148 ();
 FILLCELL_X32 FILLER_14_153 ();
 FILLCELL_X16 FILLER_14_185 ();
 FILLCELL_X8 FILLER_14_201 ();
 FILLCELL_X2 FILLER_14_209 ();
 FILLCELL_X1 FILLER_14_211 ();
 FILLCELL_X4 FILLER_14_229 ();
 FILLCELL_X2 FILLER_14_233 ();
 FILLCELL_X16 FILLER_14_238 ();
 FILLCELL_X2 FILLER_14_254 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X4 FILLER_15_65 ();
 FILLCELL_X2 FILLER_15_69 ();
 FILLCELL_X1 FILLER_15_71 ();
 FILLCELL_X2 FILLER_15_80 ();
 FILLCELL_X16 FILLER_15_93 ();
 FILLCELL_X4 FILLER_15_109 ();
 FILLCELL_X2 FILLER_15_113 ();
 FILLCELL_X1 FILLER_15_134 ();
 FILLCELL_X16 FILLER_15_161 ();
 FILLCELL_X4 FILLER_15_177 ();
 FILLCELL_X1 FILLER_15_181 ();
 FILLCELL_X8 FILLER_15_202 ();
 FILLCELL_X1 FILLER_15_210 ();
 FILLCELL_X8 FILLER_15_215 ();
 FILLCELL_X2 FILLER_15_223 ();
 FILLCELL_X1 FILLER_15_225 ();
 FILLCELL_X16 FILLER_15_229 ();
 FILLCELL_X8 FILLER_15_245 ();
 FILLCELL_X2 FILLER_15_253 ();
 FILLCELL_X1 FILLER_15_255 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X16 FILLER_16_33 ();
 FILLCELL_X8 FILLER_16_49 ();
 FILLCELL_X4 FILLER_16_57 ();
 FILLCELL_X2 FILLER_16_61 ();
 FILLCELL_X1 FILLER_16_80 ();
 FILLCELL_X8 FILLER_16_89 ();
 FILLCELL_X4 FILLER_16_97 ();
 FILLCELL_X2 FILLER_16_101 ();
 FILLCELL_X4 FILLER_16_106 ();
 FILLCELL_X1 FILLER_16_110 ();
 FILLCELL_X2 FILLER_16_114 ();
 FILLCELL_X1 FILLER_16_116 ();
 FILLCELL_X8 FILLER_16_125 ();
 FILLCELL_X2 FILLER_16_133 ();
 FILLCELL_X8 FILLER_16_142 ();
 FILLCELL_X4 FILLER_16_150 ();
 FILLCELL_X16 FILLER_16_157 ();
 FILLCELL_X4 FILLER_16_173 ();
 FILLCELL_X2 FILLER_16_177 ();
 FILLCELL_X1 FILLER_16_179 ();
 FILLCELL_X16 FILLER_16_200 ();
 FILLCELL_X8 FILLER_16_216 ();
 FILLCELL_X4 FILLER_16_224 ();
 FILLCELL_X2 FILLER_16_228 ();
 FILLCELL_X1 FILLER_16_230 ();
 FILLCELL_X2 FILLER_16_251 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X2 FILLER_17_65 ();
 FILLCELL_X1 FILLER_17_76 ();
 FILLCELL_X4 FILLER_17_89 ();
 FILLCELL_X2 FILLER_17_95 ();
 FILLCELL_X1 FILLER_17_97 ();
 FILLCELL_X16 FILLER_17_101 ();
 FILLCELL_X8 FILLER_17_117 ();
 FILLCELL_X2 FILLER_17_125 ();
 FILLCELL_X1 FILLER_17_127 ();
 FILLCELL_X16 FILLER_17_150 ();
 FILLCELL_X8 FILLER_17_166 ();
 FILLCELL_X4 FILLER_17_174 ();
 FILLCELL_X2 FILLER_17_178 ();
 FILLCELL_X1 FILLER_17_180 ();
 FILLCELL_X1 FILLER_17_185 ();
 FILLCELL_X1 FILLER_17_190 ();
 FILLCELL_X1 FILLER_17_195 ();
 FILLCELL_X4 FILLER_17_218 ();
 FILLCELL_X2 FILLER_17_222 ();
 FILLCELL_X4 FILLER_17_227 ();
 FILLCELL_X2 FILLER_17_231 ();
 FILLCELL_X16 FILLER_17_237 ();
 FILLCELL_X2 FILLER_17_253 ();
 FILLCELL_X1 FILLER_17_255 ();
 FILLCELL_X16 FILLER_18_1 ();
 FILLCELL_X8 FILLER_18_17 ();
 FILLCELL_X2 FILLER_18_25 ();
 FILLCELL_X32 FILLER_18_30 ();
 FILLCELL_X4 FILLER_18_62 ();
 FILLCELL_X2 FILLER_18_66 ();
 FILLCELL_X1 FILLER_18_68 ();
 FILLCELL_X4 FILLER_18_90 ();
 FILLCELL_X2 FILLER_18_94 ();
 FILLCELL_X1 FILLER_18_96 ();
 FILLCELL_X2 FILLER_18_101 ();
 FILLCELL_X4 FILLER_18_107 ();
 FILLCELL_X8 FILLER_18_115 ();
 FILLCELL_X2 FILLER_18_123 ();
 FILLCELL_X4 FILLER_18_142 ();
 FILLCELL_X2 FILLER_18_146 ();
 FILLCELL_X1 FILLER_18_148 ();
 FILLCELL_X32 FILLER_18_159 ();
 FILLCELL_X8 FILLER_18_191 ();
 FILLCELL_X4 FILLER_18_199 ();
 FILLCELL_X2 FILLER_18_203 ();
 FILLCELL_X1 FILLER_18_205 ();
 FILLCELL_X1 FILLER_18_211 ();
 FILLCELL_X32 FILLER_18_215 ();
 FILLCELL_X8 FILLER_18_247 ();
 FILLCELL_X1 FILLER_18_255 ();
 FILLCELL_X16 FILLER_19_1 ();
 FILLCELL_X8 FILLER_19_17 ();
 FILLCELL_X2 FILLER_19_25 ();
 FILLCELL_X1 FILLER_19_27 ();
 FILLCELL_X32 FILLER_19_31 ();
 FILLCELL_X1 FILLER_19_63 ();
 FILLCELL_X16 FILLER_19_71 ();
 FILLCELL_X8 FILLER_19_87 ();
 FILLCELL_X1 FILLER_19_95 ();
 FILLCELL_X2 FILLER_19_101 ();
 FILLCELL_X1 FILLER_19_103 ();
 FILLCELL_X16 FILLER_19_111 ();
 FILLCELL_X4 FILLER_19_127 ();
 FILLCELL_X2 FILLER_19_131 ();
 FILLCELL_X1 FILLER_19_144 ();
 FILLCELL_X32 FILLER_19_165 ();
 FILLCELL_X16 FILLER_19_197 ();
 FILLCELL_X8 FILLER_19_213 ();
 FILLCELL_X1 FILLER_19_221 ();
 FILLCELL_X4 FILLER_19_225 ();
 FILLCELL_X2 FILLER_19_229 ();
 FILLCELL_X2 FILLER_19_235 ();
 FILLCELL_X4 FILLER_19_240 ();
 FILLCELL_X8 FILLER_19_247 ();
 FILLCELL_X1 FILLER_19_255 ();
 FILLCELL_X16 FILLER_20_1 ();
 FILLCELL_X8 FILLER_20_17 ();
 FILLCELL_X8 FILLER_20_28 ();
 FILLCELL_X1 FILLER_20_36 ();
 FILLCELL_X2 FILLER_20_54 ();
 FILLCELL_X1 FILLER_20_56 ();
 FILLCELL_X1 FILLER_20_60 ();
 FILLCELL_X16 FILLER_20_69 ();
 FILLCELL_X8 FILLER_20_85 ();
 FILLCELL_X8 FILLER_20_96 ();
 FILLCELL_X4 FILLER_20_104 ();
 FILLCELL_X1 FILLER_20_108 ();
 FILLCELL_X1 FILLER_20_112 ();
 FILLCELL_X8 FILLER_20_118 ();
 FILLCELL_X16 FILLER_20_144 ();
 FILLCELL_X1 FILLER_20_160 ();
 FILLCELL_X4 FILLER_20_173 ();
 FILLCELL_X2 FILLER_20_177 ();
 FILLCELL_X16 FILLER_20_182 ();
 FILLCELL_X4 FILLER_20_198 ();
 FILLCELL_X4 FILLER_20_223 ();
 FILLCELL_X1 FILLER_20_227 ();
 FILLCELL_X8 FILLER_20_245 ();
 FILLCELL_X2 FILLER_20_253 ();
 FILLCELL_X1 FILLER_20_255 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X1 FILLER_21_65 ();
 FILLCELL_X16 FILLER_21_68 ();
 FILLCELL_X8 FILLER_21_84 ();
 FILLCELL_X2 FILLER_21_92 ();
 FILLCELL_X8 FILLER_21_98 ();
 FILLCELL_X4 FILLER_21_106 ();
 FILLCELL_X1 FILLER_21_110 ();
 FILLCELL_X8 FILLER_21_118 ();
 FILLCELL_X4 FILLER_21_126 ();
 FILLCELL_X1 FILLER_21_130 ();
 FILLCELL_X8 FILLER_21_133 ();
 FILLCELL_X4 FILLER_21_141 ();
 FILLCELL_X2 FILLER_21_145 ();
 FILLCELL_X1 FILLER_21_147 ();
 FILLCELL_X1 FILLER_21_170 ();
 FILLCELL_X1 FILLER_21_174 ();
 FILLCELL_X8 FILLER_21_189 ();
 FILLCELL_X1 FILLER_21_197 ();
 FILLCELL_X8 FILLER_21_205 ();
 FILLCELL_X4 FILLER_21_213 ();
 FILLCELL_X2 FILLER_21_217 ();
 FILLCELL_X1 FILLER_21_219 ();
 FILLCELL_X2 FILLER_21_224 ();
 FILLCELL_X1 FILLER_21_226 ();
 FILLCELL_X4 FILLER_21_230 ();
 FILLCELL_X1 FILLER_21_234 ();
 FILLCELL_X16 FILLER_21_238 ();
 FILLCELL_X2 FILLER_21_254 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_33 ();
 FILLCELL_X4 FILLER_22_41 ();
 FILLCELL_X2 FILLER_22_45 ();
 FILLCELL_X4 FILLER_22_71 ();
 FILLCELL_X2 FILLER_22_79 ();
 FILLCELL_X1 FILLER_22_81 ();
 FILLCELL_X16 FILLER_22_98 ();
 FILLCELL_X1 FILLER_22_114 ();
 FILLCELL_X1 FILLER_22_118 ();
 FILLCELL_X16 FILLER_22_144 ();
 FILLCELL_X2 FILLER_22_160 ();
 FILLCELL_X1 FILLER_22_162 ();
 FILLCELL_X8 FILLER_22_166 ();
 FILLCELL_X4 FILLER_22_174 ();
 FILLCELL_X16 FILLER_22_188 ();
 FILLCELL_X4 FILLER_22_204 ();
 FILLCELL_X1 FILLER_22_208 ();
 FILLCELL_X8 FILLER_22_220 ();
 FILLCELL_X2 FILLER_22_228 ();
 FILLCELL_X8 FILLER_22_247 ();
 FILLCELL_X1 FILLER_22_255 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X8 FILLER_23_65 ();
 FILLCELL_X4 FILLER_23_73 ();
 FILLCELL_X2 FILLER_23_77 ();
 FILLCELL_X16 FILLER_23_103 ();
 FILLCELL_X8 FILLER_23_119 ();
 FILLCELL_X4 FILLER_23_127 ();
 FILLCELL_X2 FILLER_23_131 ();
 FILLCELL_X1 FILLER_23_133 ();
 FILLCELL_X4 FILLER_23_138 ();
 FILLCELL_X1 FILLER_23_142 ();
 FILLCELL_X32 FILLER_23_147 ();
 FILLCELL_X32 FILLER_23_179 ();
 FILLCELL_X2 FILLER_23_211 ();
 FILLCELL_X1 FILLER_23_237 ();
 FILLCELL_X2 FILLER_23_241 ();
 FILLCELL_X1 FILLER_23_243 ();
 FILLCELL_X8 FILLER_23_247 ();
 FILLCELL_X1 FILLER_23_255 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X2 FILLER_24_129 ();
 FILLCELL_X4 FILLER_24_136 ();
 FILLCELL_X2 FILLER_24_140 ();
 FILLCELL_X1 FILLER_24_142 ();
 FILLCELL_X16 FILLER_24_151 ();
 FILLCELL_X2 FILLER_24_174 ();
 FILLCELL_X32 FILLER_24_180 ();
 FILLCELL_X32 FILLER_24_212 ();
 FILLCELL_X8 FILLER_24_244 ();
 FILLCELL_X4 FILLER_24_252 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X1 FILLER_25_9 ();
 FILLCELL_X16 FILLER_25_13 ();
 FILLCELL_X4 FILLER_25_29 ();
 FILLCELL_X2 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_60 ();
 FILLCELL_X32 FILLER_25_92 ();
 FILLCELL_X4 FILLER_25_124 ();
 FILLCELL_X2 FILLER_25_128 ();
 FILLCELL_X16 FILLER_25_150 ();
 FILLCELL_X4 FILLER_25_166 ();
 FILLCELL_X1 FILLER_25_170 ();
 FILLCELL_X8 FILLER_25_188 ();
 FILLCELL_X2 FILLER_25_196 ();
 FILLCELL_X32 FILLER_25_209 ();
 FILLCELL_X8 FILLER_25_241 ();
 FILLCELL_X4 FILLER_25_249 ();
 FILLCELL_X2 FILLER_25_253 ();
 FILLCELL_X1 FILLER_25_255 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X4 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_73 ();
 FILLCELL_X8 FILLER_26_105 ();
 FILLCELL_X2 FILLER_26_113 ();
 FILLCELL_X1 FILLER_26_115 ();
 FILLCELL_X8 FILLER_26_136 ();
 FILLCELL_X1 FILLER_26_144 ();
 FILLCELL_X32 FILLER_26_148 ();
 FILLCELL_X4 FILLER_26_180 ();
 FILLCELL_X8 FILLER_26_187 ();
 FILLCELL_X4 FILLER_26_195 ();
 FILLCELL_X2 FILLER_26_199 ();
 FILLCELL_X8 FILLER_26_218 ();
 FILLCELL_X2 FILLER_26_226 ();
 FILLCELL_X16 FILLER_26_231 ();
 FILLCELL_X8 FILLER_26_247 ();
 FILLCELL_X1 FILLER_26_255 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X4 FILLER_27_65 ();
 FILLCELL_X8 FILLER_27_72 ();
 FILLCELL_X4 FILLER_27_80 ();
 FILLCELL_X2 FILLER_27_84 ();
 FILLCELL_X1 FILLER_27_86 ();
 FILLCELL_X32 FILLER_27_111 ();
 FILLCELL_X32 FILLER_27_150 ();
 FILLCELL_X2 FILLER_27_182 ();
 FILLCELL_X1 FILLER_27_184 ();
 FILLCELL_X1 FILLER_27_189 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X1 FILLER_27_225 ();
 FILLCELL_X2 FILLER_27_250 ();
 FILLCELL_X1 FILLER_27_255 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X16 FILLER_28_33 ();
 FILLCELL_X8 FILLER_28_49 ();
 FILLCELL_X2 FILLER_28_57 ();
 FILLCELL_X1 FILLER_28_59 ();
 FILLCELL_X32 FILLER_28_77 ();
 FILLCELL_X16 FILLER_28_109 ();
 FILLCELL_X8 FILLER_28_125 ();
 FILLCELL_X2 FILLER_28_133 ();
 FILLCELL_X1 FILLER_28_135 ();
 FILLCELL_X16 FILLER_28_153 ();
 FILLCELL_X8 FILLER_28_169 ();
 FILLCELL_X4 FILLER_28_177 ();
 FILLCELL_X1 FILLER_28_181 ();
 FILLCELL_X32 FILLER_28_199 ();
 FILLCELL_X16 FILLER_28_231 ();
 FILLCELL_X8 FILLER_28_247 ();
 FILLCELL_X1 FILLER_28_255 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X16 FILLER_29_225 ();
 FILLCELL_X8 FILLER_29_241 ();
 FILLCELL_X4 FILLER_29_249 ();
 FILLCELL_X2 FILLER_29_253 ();
 FILLCELL_X1 FILLER_29_255 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X16 FILLER_30_225 ();
 FILLCELL_X8 FILLER_30_241 ();
 FILLCELL_X4 FILLER_30_249 ();
 FILLCELL_X2 FILLER_30_253 ();
 FILLCELL_X1 FILLER_30_255 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X16 FILLER_31_225 ();
 FILLCELL_X8 FILLER_31_241 ();
 FILLCELL_X4 FILLER_31_249 ();
 FILLCELL_X2 FILLER_31_253 ();
 FILLCELL_X1 FILLER_31_255 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X4 FILLER_32_65 ();
 FILLCELL_X2 FILLER_32_69 ();
 FILLCELL_X32 FILLER_32_74 ();
 FILLCELL_X32 FILLER_32_106 ();
 FILLCELL_X32 FILLER_32_138 ();
 FILLCELL_X32 FILLER_32_170 ();
 FILLCELL_X32 FILLER_32_202 ();
 FILLCELL_X16 FILLER_32_234 ();
 FILLCELL_X4 FILLER_32_250 ();
 FILLCELL_X2 FILLER_32_254 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X4 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_104 ();
 FILLCELL_X8 FILLER_33_136 ();
 FILLCELL_X4 FILLER_33_144 ();
 FILLCELL_X2 FILLER_33_148 ();
 FILLCELL_X1 FILLER_33_150 ();
 FILLCELL_X32 FILLER_33_154 ();
 FILLCELL_X8 FILLER_33_186 ();
 FILLCELL_X4 FILLER_33_194 ();
 FILLCELL_X32 FILLER_33_201 ();
 FILLCELL_X16 FILLER_33_233 ();
 FILLCELL_X4 FILLER_33_249 ();
 FILLCELL_X2 FILLER_33_253 ();
 FILLCELL_X1 FILLER_33_255 ();
endmodule
