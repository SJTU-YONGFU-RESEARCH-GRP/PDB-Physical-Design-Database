
* cell fifo
* pin full
* pin wr_en
* pin rd_en
* pin empty
* pin PWELL
* pin NWELL
* pin clk
* pin din[1]
* pin din[2]
* pin rst_n
* pin dout[6]
* pin dout[1]
* pin dout[7]
* pin dout[0]
* pin din[4]
* pin din[7]
* pin din[6]
* pin din[0]
* pin din[3]
* pin din[5]
* pin dout[3]
* pin dout[5]
* pin dout[4]
* pin dout[2]
.SUBCKT fifo 1 2 3 4 5 6 82 191 207 323 324 325 338 381 538 546 557 558 581 582
+ 583 584 585 586
* net 1 full
* net 2 wr_en
* net 3 rd_en
* net 4 empty
* net 5 PWELL
* net 6 NWELL
* net 82 clk
* net 191 din[1]
* net 207 din[2]
* net 323 rst_n
* net 324 dout[6]
* net 325 dout[1]
* net 338 dout[7]
* net 381 dout[0]
* net 538 din[4]
* net 546 din[7]
* net 557 din[6]
* net 558 din[0]
* net 581 din[3]
* net 582 din[5]
* net 583 dout[3]
* net 584 dout[5]
* net 585 dout[4]
* net 586 dout[2]
* cell instance $1 m0 *1 266.19,4.2
X$1 78 5 6 1 BUF_X1
* cell instance $8 r0 *1 272.08,1.4
X$8 2 6 8 5 BUF_X4
* cell instance $17 r0 *1 279.11,1.4
X$17 3 6 7 5 BUF_X4
* cell instance $20 r0 *1 276.26,1.4
X$20 9 5 6 4 BUF_X1
* cell instance $25 m0 *1 268.09,217
X$25 28 24 16 5 6 21 MUX2_X1
* cell instance $26 m0 *1 264.86,217
X$26 5 616 37 34 15 6 DFF_X1
* cell instance $28 m0 *1 269.61,217
X$28 5 602 11 35 27 6 DFF_X1
* cell instance $29 m0 *1 272.84,217
X$29 11 17 18 5 6 59 MUX2_X1
* cell instance $30 m0 *1 274.17,217
X$30 18 25 28 5 6 19 MUX2_X1
* cell instance $33 m0 *1 277.21,217
X$33 32 25 29 5 6 20 MUX2_X1
* cell instance $34 m0 *1 278.54,217
X$34 30 17 32 5 6 70 MUX2_X1
* cell instance $35 m0 *1 279.87,217
X$35 29 12 30 5 6 31 MUX2_X1
* cell instance $38 m0 *1 282.15,217
X$38 5 604 30 31 27 6 DFF_X1
* cell instance $73 m0 *1 250.99,217
X$73 10 24 46 5 6 45 MUX2_X1
* cell instance $77 r0 *1 250.8,217
X$77 5 669 46 45 13 6 DFF_X1
* cell instance $79 m0 *1 260.11,217
X$79 26 25 10 5 6 14 MUX2_X1
* cell instance $80 m0 *1 258.78,217
X$80 23 17 26 5 6 33 MUX2_X1
* cell instance $87 r0 *1 265.62,217
X$87 28 36 37 5 6 34 MUX2_X1
* cell instance $90 r0 *1 268.66,217
X$90 37 38 16 5 6 61 MUX2_X1
* cell instance $93 r0 *1 276.83,217
X$93 5 730 32 20 27 6 DFF_X1
* cell instance $99 r0 *1 285.95,217
X$99 5 724 40 47 42 6 DFF_X1
* cell instance $100 r0 *1 289.18,217
X$100 5 722 43 41 42 6 DFF_X1
* cell instance $103 r0 *1 294.12,217
X$103 5 694 52 44 42 6 DFF_X1
* cell instance $2039 r0 *1 230.47,278.6
X$2039 582 5 6 406 BUF_X2
* cell instance $2053 m0 *1 254.41,278.6
X$2053 5 655 570 579 473 6 DFF_X1
* cell instance $2057 m0 *1 259.54,278.6
X$2057 5 658 547 571 473 6 DFF_X1
* cell instance $12661 m0 *1 232.18,281.4
X$12661 581 5 6 469 BUF_X2
* cell instance $12874 m0 *1 235.22,273
X$12874 538 5 6 405 CLKBUF_X2
* cell instance $12884 r0 *1 248.9,273
X$12884 560 243 561 5 6 472 MUX2_X1
* cell instance $12888 m0 *1 252.13,273
X$12888 5 631 515 539 473 6 DFF_X1
* cell instance $12892 r0 *1 258.02,273
X$12892 540 39 564 5 6 474 MUX2_X1
* cell instance $12896 r0 *1 260.68,273
X$12896 547 353 548 5 6 564 MUX2_X1
* cell instance $12902 r0 *1 267.14,273
X$12902 5 675 542 566 473 6 DFF_X1
* cell instance $12904 m0 *1 268.28,273
X$12904 549 243 542 5 6 541 MUX2_X1
* cell instance $12906 r0 *1 270.37,273
X$12906 542 230 29 5 6 566 MUX2_X1
* cell instance $12908 r0 *1 272.46,273
X$12908 469 5 6 29 BUF_X2
* cell instance $12909 r0 *1 273.22,273
X$12909 5 681 550 567 453 6 DFF_X1
* cell instance $12915 r0 *1 280.82,273
X$12915 552 292 97 5 6 551 MUX2_X1
* cell instance $12918 r0 *1 282.34,273
X$12918 573 353 552 5 6 543 MUX2_X1
* cell instance $12922 r0 *1 287.28,273
X$12922 437 288 569 5 6 568 MUX2_X1
* cell instance $12924 r0 *1 288.61,273
X$12924 574 17 569 5 6 553 MUX2_X1
* cell instance $12925 r0 *1 289.94,273
X$12925 553 39 543 5 6 486 MUX2_X1
* cell instance $12929 r0 *1 293.36,273
X$12929 437 5 6 97 BUF_X2
* cell instance $12932 r0 *1 294.5,273
X$12932 555 230 97 5 6 554 MUX2_X1
* cell instance $12933 r0 *1 295.83,273
X$12933 545 243 555 5 6 544 MUX2_X1
* cell instance $12934 r0 *1 297.16,273
X$12934 437 280 545 5 6 556 MUX2_X1
* cell instance $12940 r0 *1 302.86,273
X$12940 557 5 6 437 CLKBUF_X2
* cell instance $16515 r0 *1 241.87,488.6
X$16515 468 5 6 583 BUF_X1
* cell instance $16516 r0 *1 242.44,488.6
X$16516 428 5 6 586 BUF_X1
* cell instance $16517 r0 *1 243.01,488.6
X$16517 433 5 6 584 BUF_X1
* cell instance $16519 r0 *1 245.1,488.6
X$16519 467 5 6 585 BUF_X1
* cell instance $17151 m0 *1 246.24,231
X$17151 5 621 155 139 84 6 DFF_X1
* cell instance $17155 r0 *1 249.85,231
X$17155 155 6 128 5 BUF_X4
* cell instance $17157 r0 *1 251.18,231
X$17157 128 146 130 5 6 129 OR3_X1
* cell instance $17158 m0 *1 251.75,231
X$17158 90 129 131 5 139 6 AOI21_X1
* cell instance $17159 r0 *1 252.13,231
X$17159 130 146 128 6 131 5 OAI21_X1
* cell instance $17165 r0 *1 256.88,231
X$17165 137 5 6 13 CLKBUF_X3
* cell instance $17168 m0 *1 257.64,231
X$17168 141 5 6 132 BUF_X2
* cell instance $17169 r0 *1 257.83,231
X$17169 13 5 6 INV_X4
* cell instance $17172 r0 *1 259.16,231
X$17172 109 128 5 6 183 XNOR2_X2
* cell instance $17174 r0 *1 261.44,231
X$17174 158 144 109 5 6 108 NAND3_X1
* cell instance $17179 r0 *1 264.67,231
X$17179 147 135 146 5 6 145 NOR3_X1
* cell instance $17180 m0 *1 264.86,231
X$17180 8 5 6 135 INV_X1
* cell instance $17181 m0 *1 265.24,231
X$17181 8 96 104 6 5 130 OAI21_X2
* cell instance $17183 r0 *1 266.19,231
X$17183 164 5 6 78 INV_X2
* cell instance $17187 r0 *1 267.9,231
X$17187 8 150 5 163 6 NAND2_X4
* cell instance $17188 r0 *1 269.61,231
X$17188 150 5 6 90 INV_X2
* cell instance $17189 r0 *1 270.18,231
X$17189 90 91 5 6 165 OR2_X1
* cell instance $17192 r0 *1 272.08,231
X$17192 157 91 158 5 6 187 MUX2_X1
* cell instance $17194 r0 *1 273.41,231
X$17194 5 136 152 143 27 6 DFF_X1
* cell instance $17195 m0 *1 275.69,231
X$17195 136 91 144 5 6 156 MUX2_X1
* cell instance $17196 r0 *1 276.64,231
X$17196 151 156 6 5 143 AND2_X1
* cell instance $17201 r0 *1 280.06,231
X$17201 137 5 6 27 CLKBUF_X3
* cell instance $17202 r0 *1 281.01,231
X$17202 27 5 6 741 INV_X1
* cell instance $17207 r0 *1 286.33,231
X$17207 154 25 153 5 6 140 MUX2_X1
* cell instance $17208 r0 *1 287.66,231
X$17208 5 704 154 140 42 6 DFF_X1
* cell instance $17211 r0 *1 291.27,231
X$17211 137 5 6 42 CLKBUF_X3
* cell instance $17212 r0 *1 292.22,231
X$17212 42 5 6 742 INV_X1
* cell instance $20892 m0 *1 237.88,261.8
X$20892 405 216 442 5 6 441 MUX2_X1
* cell instance $20942 r0 *1 236.55,261.8
X$20942 5 693 442 441 431 6 DFF_X1
* cell instance $20947 m0 *1 243.58,261.8
X$20947 442 158 454 5 6 423 MUX2_X1
* cell instance $20949 m0 *1 245.1,261.8
X$20949 137 5 6 340 CLKBUF_X3
* cell instance $20951 m0 *1 246.24,261.8
X$20951 406 216 432 5 6 443 MUX2_X1
* cell instance $20952 m0 *1 247.57,261.8
X$20952 5 617 432 443 431 6 DFF_X1
* cell instance $20955 r0 *1 241.49,261.8
X$20955 5 705 454 466 340 6 DFF_X1
* cell instance $20956 r0 *1 244.72,261.8
X$20956 454 241 57 5 6 466 MUX2_X1
* cell instance $20957 r0 *1 246.05,261.8
X$20957 340 5 6 739 INV_X2
* cell instance $20960 r0 *1 251.18,261.8
X$20960 5 683 444 445 358 6 DFF_X1
* cell instance $20961 m0 *1 252.51,261.8
X$20961 444 241 116 5 6 445 MUX2_X1
* cell instance $20962 m0 *1 251.18,261.8
X$20962 432 158 444 5 6 408 MUX2_X1
* cell instance $20966 m0 *1 258.59,261.8
X$20966 114 433 151 5 6 449 NAND3_X1
* cell instance $20967 m0 *1 259.35,261.8
X$20967 409 458 6 5 447 AND2_X1
* cell instance $20969 m0 *1 260.3,261.8
X$20969 137 5 6 358 CLKBUF_X3
* cell instance $20970 m0 *1 261.25,261.8
X$20970 283 447 449 6 448 5 OAI21_X1
* cell instance $20977 r0 *1 257.07,261.8
X$20977 391 455 6 5 456 AND2_X1
* cell instance $20978 r0 *1 257.83,261.8
X$20978 114 467 151 5 6 457 NAND3_X1
* cell instance $20980 r0 *1 258.78,261.8
X$20980 5 448 358 590 433 6 DFF_X2
* cell instance $20986 r0 *1 268.28,261.8
X$20986 114 468 151 5 6 459 NAND3_X1
* cell instance $20988 m0 *1 269.42,261.8
X$20988 469 226 450 5 6 451 MUX2_X1
* cell instance $20990 m0 *1 270.75,261.8
X$20990 5 656 450 451 453 6 DFF_X1
* cell instance $20996 r0 *1 273.41,261.8
X$20996 469 216 434 5 6 461 MUX2_X1
* cell instance $20998 m0 *1 275.31,261.8
X$20998 434 158 435 5 6 452 MUX2_X1
* cell instance $21000 m0 *1 276.64,261.8
X$21000 435 241 29 5 6 446 MUX2_X1
* cell instance $21004 m0 *1 280.44,261.8
X$21004 171 6 353 5 BUF_X4
* cell instance $21005 m0 *1 281.77,261.8
X$21005 5 654 413 412 316 6 DFF_X1
* cell instance $21009 r0 *1 276.07,261.8
X$21009 5 686 435 446 453 6 DFF_X1
* cell instance $21011 r0 *1 279.49,261.8
X$21011 137 5 6 453 CLKBUF_X3
* cell instance $21012 r0 *1 280.44,261.8
X$21012 453 5 6 740 INV_X1
* cell instance $21016 m0 *1 285.57,261.8
X$21016 437 216 414 5 6 436 MUX2_X1
* cell instance $21019 m0 *1 288.42,261.8
X$21019 437 226 415 5 6 438 MUX2_X1
* cell instance $21023 m0 *1 294.5,261.8
X$21023 137 5 6 318 CLKBUF_X3
* cell instance $21024 m0 *1 295.45,261.8
X$21024 318 5 6 CLKBUF_X1
* cell instance $21029 m0 *1 301.53,261.8
X$21029 420 171 439 5 6 440 MUX2_X1
* cell instance $21061 r0 *1 285.76,261.8
X$21061 5 727 414 436 462 6 DFF_X1
* cell instance $21064 r0 *1 289.94,261.8
X$21064 172 6 65 5 BUF_X4
* cell instance $21068 r0 *1 292.6,261.8
X$21068 137 5 6 462 CLKBUF_X3
* cell instance $21071 r0 *1 294.12,261.8
X$21071 273 465 206 485 5 6 463 AOI22_X1
* cell instance $21073 r0 *1 295.83,261.8
X$21073 440 172 478 5 6 465 MUX2_X1
* cell instance $21232 m0 *1 243.39,253.4
X$21232 5 638 312 352 340 6 DFF_X1
* cell instance $21237 m0 *1 254.41,253.4
X$21237 5 640 354 364 358 6 DFF_X1
* cell instance $21238 m0 *1 257.64,253.4
X$21238 354 353 333 5 6 372 MUX2_X1
* cell instance $21239 m0 *1 258.97,253.4
X$21239 372 39 356 5 6 355 MUX2_X1
* cell instance $21244 r0 *1 259.54,253.4
X$21244 373 247 357 5 6 356 MUX2_X1
* cell instance $21245 m0 *1 260.87,253.4
X$21245 357 292 10 5 6 385 MUX2_X1
* cell instance $21247 m0 *1 262.2,253.4
X$21247 5 643 357 385 358 6 DFF_X1
* cell instance $21250 r0 *1 260.87,253.4
X$21250 10 317 373 5 6 402 MUX2_X1
* cell instance $21255 r0 *1 267.71,253.4
X$21255 5 668 359 384 358 6 DFF_X1
* cell instance $21257 m0 *1 268.85,253.4
X$21257 28 315 359 5 6 384 MUX2_X1
* cell instance $21260 m0 *1 272.27,253.4
X$21260 359 353 350 5 6 371 MUX2_X1
* cell instance $21263 m0 *1 275.12,253.4
X$21263 371 39 375 5 6 331 MUX2_X1
* cell instance $21265 m0 *1 276.64,253.4
X$21265 370 292 28 5 6 369 MUX2_X1
* cell instance $21266 m0 *1 277.97,253.4
X$21266 5 606 370 369 316 6 DFF_X1
* cell instance $21269 m0 *1 282.15,253.4
X$21269 368 241 50 5 6 376 MUX2_X1
* cell instance $21276 r0 *1 273.6,253.4
X$21276 28 317 374 5 6 386 MUX2_X1
* cell instance $21278 r0 *1 275.12,253.4
X$21278 374 247 370 5 6 375 MUX2_X1
* cell instance $21283 r0 *1 281.96,253.4
X$21283 5 725 368 376 316 6 DFF_X1
* cell instance $21286 r0 *1 286.14,253.4
X$21286 377 158 368 5 6 367 MUX2_X1
* cell instance $21291 r0 *1 291.84,253.4
X$21291 378 247 383 5 6 379 MUX2_X1
* cell instance $21292 m0 *1 293.55,253.4
X$21292 134 68 197 365 5 6 360 AOI22_X1
* cell instance $21293 m0 *1 292.22,253.4
X$21293 379 144 367 5 6 365 MUX2_X1
* cell instance $21294 m0 *1 294.5,253.4
X$21294 360 463 6 5 361 AND2_X1
* cell instance $21295 m0 *1 295.26,253.4
X$21295 50 233 383 5 6 363 MUX2_X1
* cell instance $21296 m0 *1 296.59,253.4
X$21296 5 612 383 363 318 6 DFF_X1
* cell instance $21297 m0 *1 299.82,253.4
X$21297 5 334 318 587 347 6 DFF_X2
* cell instance $21298 m0 *1 303.43,253.4
X$21298 283 382 336 6 380 5 OAI21_X1
* cell instance $21300 m0 *1 304.38,253.4
X$21300 283 361 337 6 362 5 OAI21_X1
* cell instance $21337 r0 *1 304.57,253.4
X$21337 5 362 318 591 343 6 DFF_X2
* cell instance $21377 r0 *1 483.74,253.4
X$21377 347 5 6 381 BUF_X1
* cell instance $21498 r0 *1 233.51,247.8
X$21498 223 289 342 5 6 341 MUX2_X1
* cell instance $21507 r0 *1 244.34,247.8
X$21507 313 144 257 5 6 314 MUX2_X1
* cell instance $21511 m0 *1 250.04,247.8
X$21511 303 230 10 5 6 327 MUX2_X1
* cell instance $21515 r0 *1 250.42,247.8
X$21515 5 663 303 327 211 6 DFF_X1
* cell instance $21518 r0 *1 257.45,247.8
X$21518 134 56 197 314 5 6 348 AOI22_X1
* cell instance $21520 m0 *1 259.54,247.8
X$21520 164 185 291 5 315 6 NAND3_X4
* cell instance $21524 r0 *1 259.92,247.8
X$21524 164 227 291 5 317 6 NAND3_X4
* cell instance $21526 m0 *1 264.1,247.8
X$21526 164 185 259 5 289 6 NAND3_X4
* cell instance $21528 m0 *1 266.57,247.8
X$21528 164 227 259 5 280 6 NAND3_X4
* cell instance $21532 m0 *1 269.42,247.8
X$21532 82 5 6 137 CLKBUF_X3
* cell instance $21535 m0 *1 280.25,247.8
X$21535 5 615 293 309 316 6 DFF_X1
* cell instance $21536 m0 *1 283.48,247.8
X$21536 328 17 293 5 6 308 MUX2_X1
* cell instance $21538 m0 *1 285,247.8
X$21538 244 288 294 5 6 310 MUX2_X1
* cell instance $21540 m0 *1 286.52,247.8
X$21540 5 614 294 310 318 6 DFF_X1
* cell instance $21546 r0 *1 280.06,247.8
X$21546 5 698 328 330 316 6 DFF_X1
* cell instance $21547 r0 *1 283.29,247.8
X$21547 153 317 328 5 6 330 MUX2_X1
* cell instance $21549 r0 *1 284.81,247.8
X$21549 153 315 319 5 6 326 MUX2_X1
* cell instance $21550 r0 *1 286.14,247.8
X$21550 5 692 319 326 318 6 DFF_X1
* cell instance $21551 r0 *1 289.37,247.8
X$21551 319 17 294 5 6 320 MUX2_X1
* cell instance $21553 m0 *1 290.13,247.8
X$21553 320 39 308 5 6 307 MUX2_X1
* cell instance $21555 m0 *1 292.03,247.8
X$21555 244 5 6 153 BUF_X2
* cell instance $21558 m0 *1 292.98,247.8
X$21558 273 304 307 206 5 6 306 AOI22_X1
* cell instance $21560 m0 *1 294.5,247.8
X$21560 305 306 6 5 321 AND2_X1
* cell instance $21563 m0 *1 296.02,247.8
X$21563 301 172 282 5 6 304 MUX2_X1
* cell instance $21566 m0 *1 299.06,247.8
X$21566 295 171 265 5 6 301 MUX2_X1
* cell instance $21567 m0 *1 300.39,247.8
X$21567 244 289 295 5 6 296 MUX2_X1
* cell instance $21606 r0 *1 306.09,247.8
X$21606 323 5 6 150 CLKBUF_X3
* cell instance $21710 m0 *1 231.04,250.6
X$21710 5 642 342 341 340 6 DFF_X1
* cell instance $21757 r0 *1 232.75,250.6
X$21757 5 731 332 339 340 6 DFF_X1
* cell instance $21758 m0 *1 234.84,250.6
X$21758 342 243 332 5 6 345 MUX2_X1
* cell instance $21763 m0 *1 238.64,250.6
X$21763 223 226 311 5 6 344 MUX2_X1
* cell instance $21766 r0 *1 235.98,250.6
X$21766 223 260 332 5 6 339 MUX2_X1
* cell instance $21769 r0 *1 238.26,250.6
X$21769 5 716 311 344 340 6 DFF_X1
* cell instance $21772 m0 *1 242.82,250.6
X$21772 311 247 312 5 6 313 MUX2_X1
* cell instance $21777 r0 *1 243.39,250.6
X$21777 10 233 312 5 6 352 MUX2_X1
* cell instance $21780 r0 *1 246.62,250.6
X$21780 223 5 6 10 BUF_X2
* cell instance $21785 r0 *1 250.23,250.6
X$21785 223 288 333 5 6 346 MUX2_X1
* cell instance $21787 m0 *1 250.61,250.6
X$21787 345 65 290 5 6 329 MUX2_X1
* cell instance $21798 r0 *1 251.94,250.6
X$21798 5 662 333 346 211 6 DFF_X1
* cell instance $21800 r0 *1 255.36,250.6
X$21800 10 315 354 5 6 364 MUX2_X1
* cell instance $21803 r0 *1 257.83,250.6
X$21803 348 349 6 5 366 AND2_X1
* cell instance $21805 r0 *1 258.78,250.6
X$21805 273 329 206 355 5 6 349 AOI22_X1
* cell instance $21809 r0 *1 269.23,250.6
X$21809 208 288 350 5 6 351 MUX2_X1
* cell instance $21810 r0 *1 270.56,250.6
X$21810 5 689 350 351 316 6 DFF_X1
* cell instance $21818 r0 *1 300.2,250.6
X$21818 321 283 335 6 334 5 OAI21_X1
* cell instance $21821 r0 *1 301.53,250.6
X$21821 114 347 151 5 6 335 NAND3_X1
* cell instance $21822 r0 *1 302.29,250.6
X$21822 5 380 318 592 322 6 DFF_X2
* cell instance $21823 m0 *1 304.19,250.6
X$21823 114 322 150 5 6 336 NAND3_X1
* cell instance $21828 m0 *1 323.19,250.6
X$21828 558 5 6 244 BUF_X2
* cell instance $21857 r0 *1 305.9,250.6
X$21857 114 343 150 5 6 337 NAND3_X1
* cell instance $21899 r0 *1 484.12,250.6
X$21899 343 5 6 338 BUF_X1
* cell instance $21901 m0 *1 486.4,250.6
X$21901 322 5 6 324 BUF_X1
* cell instance $21903 m0 *1 486.97,250.6
X$21903 284 5 6 325 BUF_X1
* cell instance $22027 r0 *1 236.36,256.2
X$22027 5 700 387 398 340 6 DFF_X1
* cell instance $22030 r0 *1 240.16,256.2
X$22030 5 665 400 399 340 6 DFF_X1
* cell instance $22035 m0 *1 243.2,256.2
X$22035 57 233 400 5 6 399 MUX2_X1
* cell instance $22038 r0 *1 243.39,256.2
X$22038 387 247 400 5 6 422 MUX2_X1
* cell instance $22040 m0 *1 248.9,256.2
X$22040 116 233 388 5 6 404 MUX2_X1
* cell instance $22043 m0 *1 250.42,256.2
X$22043 5 639 388 404 340 6 DFF_X1
* cell instance $22046 m0 *1 261.25,256.2
X$22046 5 629 373 402 358 6 DFF_X1
* cell instance $22049 m0 *1 272.08,256.2
X$22049 5 632 374 386 316 6 DFF_X1
* cell instance $22053 m0 *1 284.62,256.2
X$22053 5 608 377 397 318 6 DFF_X1
* cell instance $22055 m0 *1 289.37,256.2
X$22055 396 226 378 5 6 395 MUX2_X1
* cell instance $22056 m0 *1 290.7,256.2
X$22056 5 630 378 395 318 6 DFF_X1
* cell instance $22102 r0 *1 285.76,256.2
X$22102 396 216 377 5 6 397 MUX2_X1
* cell instance $22462 m0 *1 237.5,259
X$22462 405 226 387 5 6 398 MUX2_X1
* cell instance $22468 m0 *1 244.34,259
X$22468 422 144 423 5 6 389 MUX2_X1
* cell instance $22470 m0 *1 246.43,259
X$22470 5 641 407 424 340 6 DFF_X1
* cell instance $22471 m0 *1 249.66,259
X$22471 407 247 388 5 6 425 MUX2_X1
* cell instance $22477 r0 *1 245.29,259
X$22477 137 5 6 431 CLKBUF_X3
* cell instance $22480 r0 *1 247.19,259
X$22480 406 226 407 5 6 424 MUX2_X1
* cell instance $22483 m0 *1 252.13,259
X$22483 425 144 408 5 6 403 MUX2_X1
* cell instance $22488 r0 *1 255.74,259
X$22488 5 390 358 588 428 6 DFF_X2
* cell instance $22489 m0 *1 256.31,259
X$22489 134 89 197 389 5 6 391 AOI22_X1
* cell instance $22491 m0 *1 257.26,259
X$22491 283 366 392 6 390 5 OAI21_X1
* cell instance $22492 m0 *1 258.02,259
X$22492 114 428 151 5 6 392 NAND3_X1
* cell instance $22493 m0 *1 258.78,259
X$22493 134 204 197 403 5 6 409 AOI22_X1
* cell instance $22497 m0 *1 270.37,259
X$22497 5 633 410 429 316 6 DFF_X1
* cell instance $22505 r0 *1 270.94,259
X$22505 29 233 410 5 6 429 MUX2_X1
* cell instance $22506 r0 *1 272.27,259
X$22506 450 247 410 5 6 430 MUX2_X1
* cell instance $22509 r0 *1 274.17,259
X$22509 430 144 452 5 6 411 MUX2_X1
* cell instance $22510 m0 *1 274.93,259
X$22510 134 72 197 411 5 6 401 AOI22_X1
* cell instance $22515 m0 *1 285.19,259
X$22515 171 6 247 5 BUF_X4
* cell instance $22518 m0 *1 293.36,259
X$22518 134 120 197 426 5 6 394 AOI22_X1
* cell instance $22519 m0 *1 294.31,259
X$22519 394 417 6 5 382 AND2_X1
* cell instance $22520 m0 *1 295.07,259
X$22520 97 233 393 5 6 418 MUX2_X1
* cell instance $22526 r0 *1 278.92,259
X$22526 316 5 6 735 INV_X2
* cell instance $22527 r0 *1 279.49,259
X$22527 137 5 6 316 CLKBUF_X3
* cell instance $22529 r0 *1 280.82,259
X$22529 171 6 158 5 BUF_X4
* cell instance $22530 r0 *1 282.15,259
X$22530 413 241 97 5 6 412 MUX2_X1
* cell instance $22534 r0 *1 285.95,259
X$22534 414 158 413 5 6 427 MUX2_X1
* cell instance $22537 r0 *1 288.42,259
X$22537 5 664 415 438 462 6 DFF_X1
* cell instance $22538 r0 *1 291.65,259
X$22538 415 247 393 5 6 416 MUX2_X1
* cell instance $22539 r0 *1 292.98,259
X$22539 416 144 427 5 6 426 MUX2_X1
* cell instance $22543 r0 *1 295.64,259
X$22543 5 715 393 418 318 6 DFF_X1
* cell instance $22546 r0 *1 300.01,259
X$22546 5 720 420 419 318 6 DFF_X1
* cell instance $22548 m0 *1 300.58,259
X$22548 396 289 420 5 6 419 MUX2_X1
* cell instance $22549 m0 *1 302.48,259
X$22549 396 260 439 5 6 421 MUX2_X1
* cell instance $22587 r0 *1 303.24,259
X$22587 5 718 439 421 318 6 DFF_X1
* cell instance $22693 m0 *1 231.61,267.4
X$22693 5 646 507 484 431 6 DFF_X1
* cell instance $22694 m0 *1 234.84,267.4
X$22694 406 260 507 5 6 484 MUX2_X1
* cell instance $22744 r0 *1 236.55,267.4
X$22744 5 695 471 508 431 6 DFF_X1
* cell instance $22745 m0 *1 237.5,267.4
X$22745 405 289 471 5 6 508 MUX2_X1
* cell instance $22751 m0 *1 241.49,267.4
X$22751 405 260 495 5 6 527 MUX2_X1
* cell instance $22752 m0 *1 242.82,267.4
X$22752 471 243 495 5 6 490 MUX2_X1
* cell instance $22753 m0 *1 244.15,267.4
X$22753 405 5 6 57 BUF_X2
* cell instance $22756 r0 *1 239.78,267.4
X$22756 5 726 495 527 431 6 DFF_X1
* cell instance $22761 r0 *1 245.86,267.4
X$22761 405 280 514 5 6 528 MUX2_X1
* cell instance $22764 r0 *1 247.76,267.4
X$22764 514 243 497 5 6 496 MUX2_X1
* cell instance $22766 m0 *1 248.33,267.4
X$22766 490 65 496 5 6 494 MUX2_X1
* cell instance $22768 m0 *1 258.78,267.4
X$22768 273 494 206 500 5 6 455 AOI22_X1
* cell instance $22769 m0 *1 259.73,267.4
X$22769 5 618 475 489 358 6 DFF_X1
* cell instance $22774 m0 *1 271.51,267.4
X$22774 273 511 206 510 5 6 460 AOI22_X1
* cell instance $22778 m0 *1 280.25,267.4
X$22778 5 613 502 509 453 6 DFF_X1
* cell instance $22782 r0 *1 249.09,267.4
X$22782 497 230 57 5 6 529 MUX2_X1
* cell instance $22787 r0 *1 255.55,267.4
X$22787 57 315 498 5 6 530 MUX2_X1
* cell instance $22789 r0 *1 257.26,267.4
X$22789 498 353 515 5 6 499 MUX2_X1
* cell instance $22791 r0 *1 258.78,267.4
X$22791 499 39 512 5 6 500 MUX2_X1
* cell instance $22793 r0 *1 260.87,267.4
X$22793 57 317 516 5 6 533 MUX2_X1
* cell instance $22794 r0 *1 262.2,267.4
X$22794 516 353 475 5 6 512 MUX2_X1
* cell instance $22798 r0 *1 268.47,267.4
X$22798 525 65 541 5 6 511 MUX2_X1
* cell instance $22802 r0 *1 271.13,267.4
X$22802 29 317 535 5 6 534 MUX2_X1
* cell instance $22804 r0 *1 273.98,267.4
X$22804 501 39 518 5 6 510 MUX2_X1
* cell instance $22809 r0 *1 279.68,267.4
X$22809 5 672 519 536 453 6 DFF_X1
* cell instance $22810 r0 *1 282.91,267.4
X$22810 502 292 50 5 6 509 MUX2_X1
* cell instance $22814 r0 *1 285.57,267.4
X$22814 5 667 503 520 462 6 DFF_X1
* cell instance $22816 m0 *1 286.14,267.4
X$22816 50 315 503 5 6 520 MUX2_X1
* cell instance $22817 m0 *1 288.23,267.4
X$22817 503 17 476 5 6 504 MUX2_X1
* cell instance $22823 r0 *1 288.99,267.4
X$22823 504 39 532 5 6 485 MUX2_X1
* cell instance $22827 r0 *1 294.31,267.4
X$22827 396 5 6 50 BUF_X2
* cell instance $22828 r0 *1 295.07,267.4
X$22828 396 280 477 5 6 505 MUX2_X1
* cell instance $22830 m0 *1 295.26,267.4
X$22830 5 601 477 505 462 6 DFF_X1
* cell instance $22832 m0 *1 299.44,267.4
X$22832 5 610 506 479 462 6 DFF_X1
* cell instance $22867 r0 *1 300.39,267.4
X$22867 437 289 506 5 6 479 MUX2_X1
* cell instance $22977 m0 *1 234.08,270.2
X$22977 469 289 524 5 6 523 MUX2_X1
* cell instance $22978 m0 *1 235.41,270.2
X$22978 524 243 513 5 6 525 MUX2_X1
* cell instance $22979 m0 *1 236.74,270.2
X$22979 469 260 513 5 6 526 MUX2_X1
* cell instance $22984 m0 *1 244.53,270.2
X$22984 5 636 514 528 431 6 DFF_X1
* cell instance $23045 r0 *1 232.18,270.2
X$23045 5 713 524 523 431 6 DFF_X1
* cell instance $23046 r0 *1 235.41,270.2
X$23046 5 670 513 526 431 6 DFF_X1
* cell instance $23050 m0 *1 248.9,270.2
X$23050 5 628 497 529 431 6 DFF_X1
* cell instance $23053 m0 *1 254.6,270.2
X$23053 5 634 498 530 473 6 DFF_X1
* cell instance $23058 r0 *1 251.94,270.2
X$23058 405 288 515 5 6 539 MUX2_X1
* cell instance $23061 m0 *1 258.97,270.2
X$23061 5 624 516 533 473 6 DFF_X1
* cell instance $23065 m0 *1 268.85,270.2
X$23065 5 627 535 534 473 6 DFF_X1
* cell instance $23070 r0 *1 271.7,270.2
X$23070 5 679 517 537 453 6 DFF_X1
* cell instance $23071 m0 *1 274.55,270.2
X$23071 517 292 29 5 6 537 MUX2_X1
* cell instance $23072 m0 *1 273.22,270.2
X$23072 535 353 517 5 6 518 MUX2_X1
* cell instance $23078 m0 *1 280.82,270.2
X$23078 50 317 519 5 6 536 MUX2_X1
* cell instance $23079 m0 *1 282.34,270.2
X$23079 519 353 502 5 6 532 MUX2_X1
* cell instance $23088 m0 *1 289.18,270.2
X$23088 5 653 476 531 462 6 DFF_X1
* cell instance $23089 m0 *1 287.85,270.2
X$23089 396 288 476 5 6 531 MUX2_X1
* cell instance $23092 m0 *1 294.69,270.2
X$23092 521 230 50 5 6 522 MUX2_X1
* cell instance $23093 m0 *1 296.02,270.2
X$23093 5 647 521 522 462 6 DFF_X1
* cell instance $23097 m0 *1 303.24,270.2
X$23097 546 5 6 396 CLKBUF_X2
* cell instance $23220 m0 *1 231.04,264.6
X$23220 5 648 470 482 431 6 DFF_X1
* cell instance $23228 m0 *1 257.26,264.6
X$23228 283 456 457 6 493 5 OAI21_X1
* cell instance $23290 r0 *1 233.13,264.6
X$23290 406 289 470 5 6 482 MUX2_X1
* cell instance $23292 r0 *1 234.84,264.6
X$23292 470 243 507 5 6 492 MUX2_X1
* cell instance $23297 r0 *1 249.47,264.6
X$23297 492 65 472 5 6 491 MUX2_X1
* cell instance $23301 r0 *1 254.98,264.6
X$23301 5 493 473 593 467 6 DFF_X2
* cell instance $23302 m0 *1 258.59,264.6
X$23302 273 491 206 474 5 6 458 AOI22_X1
* cell instance $23305 m0 *1 260.3,264.6
X$23305 358 5 6 734 INV_X2
* cell instance $23309 r0 *1 258.59,264.6
X$23309 473 5 6 CLKBUF_X1
* cell instance $23310 r0 *1 259.16,264.6
X$23310 137 5 6 473 CLKBUF_X3
* cell instance $23312 r0 *1 260.3,264.6
X$23312 475 292 57 5 6 489 MUX2_X1
* cell instance $23316 r0 *1 266.38,264.6
X$23316 5 488 473 595 468 6 DFF_X2
* cell instance $23318 m0 *1 268.09,264.6
X$23318 283 487 459 6 488 5 OAI21_X1
* cell instance $23322 m0 *1 271.7,264.6
X$23322 401 460 6 5 487 AND2_X1
* cell instance $23325 m0 *1 273.22,264.6
X$23325 5 650 434 461 453 6 DFF_X1
* cell instance $23337 m0 *1 293.74,264.6
X$23337 273 483 206 486 5 6 417 AOI22_X1
* cell instance $23341 m0 *1 295.64,264.6
X$23341 481 172 544 5 6 483 MUX2_X1
* cell instance $23346 r0 *1 295.83,264.6
X$23346 477 243 521 5 6 478 MUX2_X1
* cell instance $23349 m0 *1 302.48,264.6
X$23349 437 260 464 5 6 480 MUX2_X1
* cell instance $23350 m0 *1 301.15,264.6
X$23350 506 171 464 5 6 481 MUX2_X1
* cell instance $23389 r0 *1 302.29,264.6
X$23389 5 661 464 480 462 6 DFF_X1
* cell instance $23542 r0 *1 244.15,275.8
X$23542 5 696 560 559 431 6 DFF_X1
* cell instance $23543 m0 *1 245.67,275.8
X$23543 406 280 560 5 6 559 MUX2_X1
* cell instance $23548 m0 *1 249.47,275.8
X$23548 561 230 116 5 6 577 MUX2_X1
* cell instance $23549 m0 *1 250.8,275.8
X$23549 406 5 6 116 CLKBUF_X3
* cell instance $23554 m0 *1 257.26,275.8
X$23554 570 353 562 5 6 540 MUX2_X1
* cell instance $23556 m0 *1 258.78,275.8
X$23556 5 622 548 563 473 6 DFF_X1
* cell instance $23557 m0 *1 262.01,275.8
X$23557 548 292 116 5 6 563 MUX2_X1
* cell instance $23560 r0 *1 247.38,275.8
X$23560 5 685 561 577 431 6 DFF_X1
* cell instance $23562 r0 *1 250.8,275.8
X$23562 406 288 562 5 6 578 MUX2_X1
* cell instance $23563 r0 *1 252.13,275.8
X$23563 5 677 562 578 473 6 DFF_X1
* cell instance $23566 r0 *1 256.5,275.8
X$23566 116 315 570 5 6 579 MUX2_X1
* cell instance $23570 r0 *1 259.92,275.8
X$23570 116 317 547 5 6 571 MUX2_X1
* cell instance $23572 m0 *1 266.57,275.8
X$23572 5 625 549 565 473 6 DFF_X1
* cell instance $23573 m0 *1 265.24,275.8
X$23573 469 280 549 5 6 565 MUX2_X1
* cell instance $23575 m0 *1 272.84,275.8
X$23575 29 315 550 5 6 567 MUX2_X1
* cell instance $23580 r0 *1 271.51,275.8
X$23580 469 288 572 5 6 580 MUX2_X1
* cell instance $23581 r0 *1 272.84,275.8
X$23581 5 673 572 580 453 6 DFF_X1
* cell instance $23583 m0 *1 274.55,275.8
X$23583 550 353 572 5 6 501 MUX2_X1
* cell instance $23585 m0 *1 280.44,275.8
X$23585 5 607 552 551 453 6 DFF_X1
* cell instance $23592 r0 *1 280.25,275.8
X$23592 5 676 573 576 453 6 DFF_X1
* cell instance $23596 r0 *1 283.48,275.8
X$23596 97 317 573 5 6 576 MUX2_X1
* cell instance $23598 r0 *1 285.19,275.8
X$23598 97 315 574 5 6 575 MUX2_X1
* cell instance $23600 m0 *1 286.33,275.8
X$23600 5 623 569 568 462 6 DFF_X1
* cell instance $23603 r0 *1 286.52,275.8
X$23603 5 687 574 575 462 6 DFF_X1
* cell instance $23605 m0 *1 293.93,275.8
X$23605 5 600 555 554 462 6 DFF_X1
* cell instance $23607 m0 *1 297.16,275.8
X$23607 5 649 545 556 462 6 DFF_X1
* cell instance $33403 r0 *1 233.13,242.2
X$33403 5 688 276 285 211 6 DFF_X1
* cell instance $33408 r0 *1 239.21,242.2
X$33408 5 671 269 268 211 6 DFF_X1
* cell instance $33413 m0 *1 251.94,242.2
X$33413 151 251 6 5 272 AND2_X1
* cell instance $33414 m0 *1 252.7,242.2
X$33414 252 130 194 5 6 251 MUX2_X1
* cell instance $33416 m0 *1 254.22,242.2
X$33416 212 225 252 6 5 253 HA_X1
* cell instance $33417 m0 *1 256.12,242.2
X$33417 212 194 596 6 5 271 HA_X1
* cell instance $33419 m0 *1 258.21,242.2
X$33419 253 6 185 5 BUF_X4
* cell instance $33421 m0 *1 259.73,242.2
X$33421 5 159 128 163 291 6 NOR3_X4
* cell instance $33423 m0 *1 262.58,242.2
X$33423 228 128 5 6 242 OR2_X2
* cell instance $33425 m0 *1 263.72,242.2
X$33425 148 242 241 5 6 NOR2_X4
* cell instance $33426 m0 *1 265.43,242.2
X$33426 242 163 256 5 6 NOR2_X4
* cell instance $33427 m0 *1 267.14,242.2
X$33427 217 185 256 5 226 6 NAND3_X4
* cell instance $33432 m0 *1 275.12,242.2
X$33432 5 644 255 231 167 6 DFF_X1
* cell instance $33435 r0 *1 242.44,242.2
X$33435 223 216 269 5 6 268 MUX2_X1
* cell instance $33439 r0 *1 251.56,242.2
X$33439 5 272 211 225 194 6 DFF_X2
* cell instance $33443 r0 *1 257.83,242.2
X$33443 271 6 229 5 BUF_X4
* cell instance $33447 r0 *1 260.49,242.2
X$33447 213 5 6 273 CLKBUF_X3
* cell instance $33449 r0 *1 261.82,242.2
X$33449 5 159 128 148 292 6 NOR3_X4
* cell instance $33450 r0 *1 264.48,242.2
X$33450 240 163 259 5 6 NOR2_X4
* cell instance $33453 r0 *1 267.14,242.2
X$33453 217 229 259 5 260 6 NAND3_X4
* cell instance $33457 r0 *1 274.36,242.2
X$33457 274 38 255 5 6 261 MUX2_X1
* cell instance $33459 m0 *1 281.96,242.2
X$33459 245 241 153 5 6 254 MUX2_X1
* cell instance $33465 r0 *1 283.48,242.2
X$33465 5 710 245 254 167 6 DFF_X1
* cell instance $33466 m0 *1 285.76,242.2
X$33466 232 247 245 5 6 249 MUX2_X1
* cell instance $33467 m0 *1 284.43,242.2
X$33467 244 216 232 5 6 236 MUX2_X1
* cell instance $33468 m0 *1 287.09,242.2
X$33468 244 226 246 5 6 250 MUX2_X1
* cell instance $33469 m0 *1 288.42,242.2
X$33469 5 626 246 250 173 6 DFF_X1
* cell instance $33470 m0 *1 291.65,242.2
X$33470 246 247 235 5 6 248 MUX2_X1
* cell instance $33471 m0 *1 292.98,242.2
X$33471 248 144 249 5 6 270 MUX2_X1
* cell instance $33476 r0 *1 293.93,242.2
X$33476 134 199 270 197 5 6 305 AOI22_X1
* cell instance $33477 m0 *1 294.88,242.2
X$33477 267 230 153 5 6 263 MUX2_X1
* cell instance $33517 r0 *1 294.88,242.2
X$33517 5 707 267 263 173 6 DFF_X1
* cell instance $33518 r0 *1 298.11,242.2
X$33518 244 260 265 5 6 264 MUX2_X1
* cell instance $33670 m0 *1 247.38,233.8
X$33670 5 660 176 180 84 6 DFF_X1
* cell instance $33672 m0 *1 251.37,233.8
X$33672 176 6 159 5 BUF_X4
* cell instance $33673 m0 *1 252.7,233.8
X$33673 159 130 161 5 6 181 OR3_X1
* cell instance $33674 m0 *1 253.65,233.8
X$33674 90 181 178 5 180 6 AOI21_X1
* cell instance $33675 m0 *1 254.41,233.8
X$33675 161 130 159 6 178 5 OAI21_X1
* cell instance $33682 r0 *1 253.65,233.8
X$33682 160 5 6 146 INV_X1
* cell instance $33685 m0 *1 257.26,233.8
X$33685 15 5 6 INV_X4
* cell instance $33687 m0 *1 258.21,233.8
X$33687 137 5 6 15 CLKBUF_X3
* cell instance $33688 m0 *1 259.16,233.8
X$33688 132 159 5 6 162 XNOR2_X2
* cell instance $33691 m0 *1 262.01,233.8
X$33691 128 159 5 6 147 NAND2_X2
* cell instance $33692 m0 *1 262.96,233.8
X$33692 147 148 25 5 6 NOR2_X4
* cell instance $33693 m0 *1 264.67,233.8
X$33693 163 146 5 6 149 NOR2_X1
* cell instance $33694 m0 *1 265.24,233.8
X$33694 149 104 96 6 5 148 OAI21_X4
* cell instance $33697 r0 *1 257.64,233.8
X$33697 5 183 162 196 205 96 6 NAND4_X4
* cell instance $33700 r0 *1 261.63,233.8
X$33700 132 5 6 221 INV_X1
* cell instance $33705 r0 *1 264.86,233.8
X$33705 147 163 186 5 6 NOR2_X4
* cell instance $33706 r0 *1 266.57,233.8
X$33706 164 185 186 5 36 6 NAND3_X4
* cell instance $33707 m0 *1 268.28,233.8
X$33707 104 96 5 6 214 OR2_X1
* cell instance $33712 m0 *1 273.03,233.8
X$33712 151 187 6 5 166 AND2_X1
* cell instance $33714 m0 *1 274.55,233.8
X$33714 152 188 157 6 5 112 HA_X1
* cell instance $33716 m0 *1 276.64,233.8
X$33716 152 6 172 5 BUF_X4
* cell instance $33724 r0 *1 273.41,233.8
X$33724 5 691 188 166 167 6 DFF_X1
* cell instance $33727 r0 *1 278.92,233.8
X$33727 167 5 6 736 INV_X2
* cell instance $33728 r0 *1 279.49,233.8
X$33728 116 36 168 5 6 190 MUX2_X1
* cell instance $33729 m0 *1 280.82,233.8
X$33729 5 651 169 189 167 6 DFF_X1
* cell instance $33731 m0 *1 284.05,233.8
X$33731 116 24 169 5 6 189 MUX2_X1
* cell instance $33734 m0 *1 287.66,233.8
X$33734 5 599 184 170 42 6 DFF_X1
* cell instance $33738 r0 *1 280.82,233.8
X$33738 5 711 168 190 167 6 DFF_X1
* cell instance $33739 r0 *1 284.05,233.8
X$33739 168 38 169 5 6 202 MUX2_X1
* cell instance $33743 r0 *1 287.85,233.8
X$33743 153 12 184 5 6 170 MUX2_X1
* cell instance $33744 r0 *1 289.18,233.8
X$33744 172 6 39 5 BUF_X4
* cell instance $33745 r0 *1 290.51,233.8
X$33745 184 171 154 5 6 182 MUX2_X1
* cell instance $33747 r0 *1 292.22,233.8
X$33747 173 5 6 738 INV_X2
* cell instance $33748 r0 *1 292.79,233.8
X$33748 137 5 6 173 CLKBUF_X3
* cell instance $33749 m0 *1 294.88,233.8
X$33749 5 659 177 179 173 6 DFF_X1
* cell instance $33750 m0 *1 293.55,233.8
X$33750 153 24 177 5 6 179 MUX2_X1
* cell instance $33782 r0 *1 293.74,233.8
X$33782 174 171 177 5 6 200 MUX2_X1
* cell instance $33783 r0 *1 295.07,233.8
X$33783 153 36 174 5 6 175 MUX2_X1
* cell instance $33786 r0 *1 298.3,233.8
X$33786 5 709 174 175 173 6 DFF_X1
* cell instance $33962 m0 *1 249.09,225.4
X$33962 5 611 75 86 13 6 DFF_X1
* cell instance $33969 m0 *1 258.97,225.4
X$33969 5 620 92 101 13 6 DFF_X1
* cell instance $33973 m0 *1 266,225.4
X$33973 103 90 5 6 77 NOR2_X1
* cell instance $33977 r0 *1 260.68,225.4
X$33977 90 102 110 5 101 6 AOI21_X1
* cell instance $33979 r0 *1 261.63,225.4
X$33979 92 6 109 5 BUF_X4
* cell instance $33984 m0 *1 267.14,225.4
X$33984 80 79 5 6 103 XOR2_X1
* cell instance $33987 m0 *1 269.23,225.4
X$33987 93 80 6 95 5 XOR2_X2
* cell instance $33991 r0 *1 267.33,225.4
X$33991 80 93 5 6 104 XNOR2_X2
* cell instance $33992 r0 *1 269.23,225.4
X$33992 93 91 113 5 6 107 OR3_X1
* cell instance $33993 r0 *1 270.18,225.4
X$33993 90 107 115 5 94 6 AOI21_X1
* cell instance $33995 r0 *1 271.13,225.4
X$33995 7 96 95 6 5 91 OAI21_X4
* cell instance $33997 m0 *1 272.08,225.4
X$33997 96 95 9 5 6 NOR2_X4
* cell instance $34001 m0 *1 286.9,225.4
X$34001 5 657 81 105 42 6 DFF_X1
* cell instance $34042 r0 *1 279.68,225.4
X$34042 5 706 126 127 27 6 DFF_X1
* cell instance $34043 r0 *1 282.91,225.4
X$34043 5 684 117 122 27 6 DFF_X1
* cell instance $34049 r0 *1 287.09,225.4
X$34049 97 12 98 5 6 106 MUX2_X1
* cell instance $34050 r0 *1 288.42,225.4
X$34050 81 25 97 5 6 105 MUX2_X1
* cell instance $34051 r0 *1 289.75,225.4
X$34051 98 17 81 5 6 121 MUX2_X1
* cell instance $34054 r0 *1 293.36,225.4
X$34054 97 24 99 5 6 100 MUX2_X1
* cell instance $34055 r0 *1 294.69,225.4
X$34055 5 729 99 100 42 6 DFF_X1
* cell instance $34208 m0 *1 260.3,228.2
X$34208 91 111 109 6 110 5 OAI21_X1
* cell instance $34209 m0 *1 261.06,228.2
X$34209 109 111 91 5 6 102 OR3_X1
* cell instance $34212 m0 *1 266.57,228.2
X$34212 112 5 6 111 INV_X1
* cell instance $34213 m0 *1 266.95,228.2
X$34213 104 96 145 6 79 5 OAI21_X1
* cell instance $34220 r0 *1 253.84,228.2
X$34220 5 666 141 123 15 6 DFF_X1
* cell instance $34221 r0 *1 257.07,228.2
X$34221 90 124 142 5 123 6 AOI21_X1
* cell instance $34222 r0 *1 257.83,228.2
X$34222 108 114 132 6 142 5 OAI21_X1
* cell instance $34224 r0 *1 258.78,228.2
X$34224 132 91 108 5 6 124 OR3_X1
* cell instance $34225 r0 *1 259.73,228.2
X$34225 109 132 6 5 133 AND2_X1
* cell instance $34226 r0 *1 260.49,228.2
X$34226 133 6 134 5 BUF_X4
* cell instance $34231 r0 *1 269.23,228.2
X$34231 134 112 5 6 113 NAND2_X1
* cell instance $34233 m0 *1 269.61,228.2
X$34233 113 114 93 6 115 5 OAI21_X1
* cell instance $34239 r0 *1 274.36,228.2
X$34239 91 6 114 5 BUF_X4
* cell instance $34241 m0 *1 279.3,228.2
X$34241 116 12 126 5 6 127 MUX2_X1
* cell instance $34245 m0 *1 282.91,228.2
X$34245 126 17 117 5 6 125 MUX2_X1
* cell instance $34246 m0 *1 284.24,228.2
X$34246 117 25 116 5 6 122 MUX2_X1
* cell instance $34255 r0 *1 291.27,228.2
X$34255 97 36 118 5 6 138 MUX2_X1
* cell instance $34257 m0 *1 292.03,228.2
X$34257 119 65 121 5 6 120 MUX2_X1
* cell instance $34258 r0 *1 292.6,228.2
X$34258 5 732 118 138 42 6 DFF_X1
* cell instance $34260 m0 *1 293.74,228.2
X$34260 118 38 99 5 6 119 MUX2_X1
* cell instance $34545 m0 *1 231.99,245
X$34545 5 645 275 299 211 6 DFF_X1
* cell instance $34547 r0 *1 232.94,245
X$34547 208 289 275 5 6 299 MUX2_X1
* cell instance $34552 m0 *1 235.6,245
X$34552 275 243 276 5 6 258 MUX2_X1
* cell instance $34555 r0 *1 235.6,245
X$34555 208 260 276 5 6 285 MUX2_X1
* cell instance $34560 m0 *1 244.34,245
X$34560 269 158 277 5 6 257 MUX2_X1
* cell instance $34563 m0 *1 247.38,245
X$34563 5 635 278 302 211 6 DFF_X1
* cell instance $34567 m0 *1 259.92,245
X$34567 164 229 291 5 288 6 NAND3_X4
* cell instance $34569 m0 *1 265.43,245
X$34569 164 229 256 5 233 6 NAND3_X4
* cell instance $34570 m0 *1 267.9,245
X$34570 5 217 164 6 BUF_X16
* cell instance $34574 r0 *1 242.06,245
X$34574 5 699 277 300 211 6 DFF_X1
* cell instance $34575 r0 *1 245.29,245
X$34575 277 241 10 5 6 300 MUX2_X1
* cell instance $34579 r0 *1 249.09,245
X$34579 223 280 278 5 6 302 MUX2_X1
* cell instance $34580 r0 *1 250.42,245
X$34580 278 38 303 5 6 290 MUX2_X1
* cell instance $34585 m0 *1 274.36,245
X$34585 258 65 261 5 6 262 MUX2_X1
* cell instance $34586 m0 *1 273.03,245
X$34586 208 280 274 5 6 279 MUX2_X1
* cell instance $34590 r0 *1 273.6,245
X$34590 5 701 274 279 167 6 DFF_X1
* cell instance $34591 m0 *1 277.02,245
X$34591 238 287 6 5 266 AND2_X1
* cell instance $34592 m0 *1 276.07,245
X$34592 273 262 206 331 5 6 287 AOI22_X1
* cell instance $34604 r0 *1 282.72,245
X$34604 293 292 153 5 6 309 MUX2_X1
* cell instance $34611 r0 *1 295.26,245
X$34611 5 702 281 286 173 6 DFF_X1
* cell instance $34612 m0 *1 296.97,245
X$34612 281 171 267 5 6 282 MUX2_X1
* cell instance $34613 m0 *1 295.64,245
X$34613 244 280 281 5 6 286 MUX2_X1
* cell instance $34614 m0 *1 298.3,245
X$34614 5 619 265 264 173 6 DFF_X1
* cell instance $34652 r0 *1 300.01,245
X$34652 5 703 295 296 173 6 DFF_X1
* cell instance $34653 r0 *1 303.24,245
X$34653 283 266 298 6 297 5 OAI21_X1
* cell instance $34654 r0 *1 304,245
X$34654 114 284 151 5 6 298 NAND3_X1
* cell instance $34658 r0 *1 306.09,245
X$34658 5 297 173 594 284 6 DFF_X2
* cell instance $34801 r0 *1 232.75,239.4
X$34801 207 5 6 223 CLKBUF_X2
* cell instance $34804 m0 *1 238.83,239.4
X$34804 208 226 210 5 6 209 MUX2_X1
* cell instance $34809 m0 *1 244.91,239.4
X$34809 201 241 28 5 6 218 MUX2_X1
* cell instance $34810 m0 *1 241.68,239.4
X$34810 5 609 224 237 211 6 DFF_X1
* cell instance $34816 r0 *1 243.2,239.4
X$34816 28 233 224 5 6 237 MUX2_X1
* cell instance $34819 r0 *1 245.48,239.4
X$34819 137 5 6 211 CLKBUF_X3
* cell instance $34820 r0 *1 246.43,239.4
X$34820 208 5 6 28 BUF_X2
* cell instance $34821 r0 *1 247.19,239.4
X$34821 211 5 6 737 INV_X2
* cell instance $34823 m0 *1 253.65,239.4
X$34823 5 222 15 212 203 6 DFF_X2
* cell instance $34828 m0 *1 262.58,239.4
X$34828 159 5 6 228 INV_X1
* cell instance $34831 m0 *1 272.08,239.4
X$34831 198 6 38 5 BUF_X4
* cell instance $34836 r0 *1 255.36,239.4
X$34836 203 225 598 6 5 239 HA_X1
* cell instance $34840 r0 *1 258.59,239.4
X$34840 239 6 227 5 BUF_X4
* cell instance $34843 r0 *1 263.15,239.4
X$34843 128 228 5 6 240 NAND2_X2
* cell instance $34844 r0 *1 264.1,239.4
X$34844 240 148 230 5 6 NOR2_X4
* cell instance $34846 r0 *1 266.57,239.4
X$34846 217 227 256 5 216 6 NAND3_X4
* cell instance $34849 r0 *1 275.5,239.4
X$34849 255 230 28 5 6 231 MUX2_X1
* cell instance $34851 m0 *1 276.07,239.4
X$34851 198 6 243 5 BUF_X4
* cell instance $34894 r0 *1 282.34,239.4
X$34894 5 712 232 236 167 6 DFF_X1
* cell instance $34899 r0 *1 288.42,239.4
X$34899 153 233 235 5 6 234 MUX2_X1
* cell instance $34900 r0 *1 289.75,239.4
X$34900 5 723 235 234 173 6 DFF_X1
* cell instance $35008 m0 *1 237.88,236.6
X$35008 5 652 193 192 84 6 DFF_X1
* cell instance $35011 m0 *1 242.82,236.6
X$35011 5 637 201 218 84 6 DFF_X1
* cell instance $35013 m0 *1 246.24,236.6
X$35013 84 5 6 733 INV_X2
* cell instance $35017 m0 *1 252.13,236.6
X$35017 203 194 597 6 5 160 HA_X1
* cell instance $35018 m0 *1 254.03,236.6
X$35018 203 194 128 5 6 161 NAND3_X1
* cell instance $35080 r0 *1 231.61,236.6
X$35080 191 5 6 208 BUF_X2
* cell instance $35085 r0 *1 238.07,236.6
X$35085 208 216 193 5 6 192 MUX2_X1
* cell instance $35086 r0 *1 239.4,236.6
X$35086 5 682 210 209 84 6 DFF_X1
* cell instance $35089 r0 *1 243.2,236.6
X$35089 210 158 224 5 6 219 MUX2_X1
* cell instance $35090 r0 *1 244.53,236.6
X$35090 193 158 201 5 6 220 MUX2_X1
* cell instance $35091 r0 *1 245.86,236.6
X$35091 219 144 220 5 6 215 MUX2_X1
* cell instance $35092 r0 *1 247.19,236.6
X$35092 137 5 6 84 CLKBUF_X3
* cell instance $35095 r0 *1 254.41,236.6
X$35095 212 130 203 5 6 195 MUX2_X1
* cell instance $35096 r0 *1 255.74,236.6
X$35096 151 195 6 5 222 AND2_X1
* cell instance $35098 m0 *1 258.59,236.6
X$35098 198 194 5 6 205 XNOR2_X2
* cell instance $35099 m0 *1 256.69,236.6
X$35099 172 203 5 6 196 XNOR2_X2
* cell instance $35103 r0 *1 260.11,236.6
X$35103 109 221 6 5 213 AND2_X1
* cell instance $35104 r0 *1 260.87,236.6
X$35104 221 109 197 5 6 NOR2_X4
* cell instance $35105 m0 *1 261.06,236.6
X$35105 132 109 206 5 6 NOR2_X4
* cell instance $35110 m0 *1 266.38,236.6
X$35110 164 229 186 5 24 6 NAND3_X4
* cell instance $35111 m0 *1 263.91,236.6
X$35111 164 227 186 5 12 6 NAND3_X4
* cell instance $35115 m0 *1 275.88,236.6
X$35115 188 5 6 198 BUF_X2
* cell instance $35116 m0 *1 276.64,236.6
X$35116 198 6 171 5 BUF_X4
* cell instance $35120 m0 *1 280.44,236.6
X$35120 137 5 6 167 CLKBUF_X3
* cell instance $35123 r0 *1 268.66,236.6
X$35123 5 217 6 214 BUF_X8
* cell instance $35124 r0 *1 271.13,236.6
X$35124 165 5 6 283 CLKBUF_X3
* cell instance $35127 r0 *1 272.65,236.6
X$35127 134 60 197 215 5 6 238 AOI22_X1
* cell instance $35131 m0 *1 282.53,236.6
X$35131 202 65 125 5 6 204 MUX2_X1
* cell instance $35138 m0 *1 288.99,236.6
X$35138 171 6 17 5 BUF_X4
* cell instance $35141 m0 *1 293.36,236.6
X$35141 200 172 182 5 6 199 MUX2_X1
* cell instance $35144 m0 *1 302.29,236.6
X$35144 150 5 6 151 CLKBUF_X3
* cell instance $35181 r0 *1 290.32,236.6
X$35181 172 6 144 5 BUF_X4
* cell instance $36001 r0 *1 255.36,214.2
X$36001 10 12 23 5 6 22 MUX2_X1
* cell instance $36002 r0 *1 256.69,214.2
X$36002 5 690 23 22 13 6 DFF_X1
* cell instance $36003 r0 *1 259.92,214.2
X$36003 5 719 26 14 15 6 DFF_X1
* cell instance $36007 r0 *1 265.62,214.2
X$36007 5 721 16 21 15 6 DFF_X1
* cell instance $36011 r0 *1 271.32,214.2
X$36011 28 12 11 5 6 35 MUX2_X1
* cell instance $36013 r0 *1 274.17,214.2
X$36013 5 717 18 19 27 6 DFF_X1
* cell instance $36592 m0 *1 246.62,219.8
X$36592 5 605 48 54 84 6 DFF_X1
* cell instance $36593 m0 *1 249.85,219.8
X$36593 10 36 48 5 6 54 MUX2_X1
* cell instance $36597 m0 *1 251.75,219.8
X$36597 48 38 46 5 6 55 MUX2_X1
* cell instance $36602 m0 *1 257.07,219.8
X$36602 55 39 33 5 6 56 MUX2_X1
* cell instance $36610 r0 *1 257.07,219.8
X$36610 5 678 63 58 13 6 DFF_X1
* cell instance $36611 r0 *1 260.3,219.8
X$36611 63 25 57 5 6 58 MUX2_X1
* cell instance $36614 m0 *1 271.89,219.8
X$36614 61 39 59 5 6 60 MUX2_X1
* cell instance $36622 r0 *1 277.02,219.8
X$36622 73 38 49 5 6 66 MUX2_X1
* cell instance $36628 m0 *1 286.71,219.8
X$36628 50 12 40 5 6 47 MUX2_X1
* cell instance $36631 m0 *1 288.61,219.8
X$36631 43 25 50 5 6 41 MUX2_X1
* cell instance $36635 m0 *1 290.89,219.8
X$36635 40 38 43 5 6 51 MUX2_X1
* cell instance $36638 m0 *1 293.17,219.8
X$36638 50 24 52 5 6 44 MUX2_X1
* cell instance $36674 r0 *1 292.79,219.8
X$36674 53 38 52 5 6 69 MUX2_X1
* cell instance $36675 r0 *1 294.12,219.8
X$36675 50 36 53 5 6 67 MUX2_X1
* cell instance $36676 r0 *1 295.45,219.8
X$36676 5 728 53 67 42 6 DFF_X1
* cell instance $36837 r0 *1 245.48,222.6
X$36837 5 697 74 83 84 6 DFF_X1
* cell instance $36838 r0 *1 248.71,222.6
X$36838 57 36 74 5 6 83 MUX2_X1
* cell instance $36839 r0 *1 250.04,222.6
X$36839 57 24 75 5 6 86 MUX2_X1
* cell instance $36841 r0 *1 251.56,222.6
X$36841 74 38 75 5 6 87 MUX2_X1
* cell instance $36845 r0 *1 255.36,222.6
X$36845 87 65 71 5 6 89 MUX2_X1
* cell instance $36848 r0 *1 257.64,222.6
X$36848 5 708 62 76 13 6 DFF_X1
* cell instance $36849 m0 *1 257.83,222.6
X$36849 57 12 62 5 6 76 MUX2_X1
* cell instance $36851 m0 *1 259.16,222.6
X$36851 62 17 63 5 6 71 MUX2_X1
* cell instance $36859 r0 *1 265.05,222.6
X$36859 5 77 13 589 80 6 DFF_X2
* cell instance $36862 m0 *1 269.23,222.6
X$36862 5 603 88 94 27 6 DFF_X1
* cell instance $36864 m0 *1 274.17,222.6
X$36864 29 36 73 5 6 85 MUX2_X1
* cell instance $36867 m0 *1 276.45,222.6
X$36867 29 24 49 5 6 64 MUX2_X1
* cell instance $36868 m0 *1 277.78,222.6
X$36868 66 65 70 5 6 72 MUX2_X1
* cell instance $36872 m0 *1 292.03,222.6
X$36872 69 65 51 5 6 68 MUX2_X1
* cell instance $36912 r0 *1 270.56,222.6
X$36912 88 5 6 93 BUF_X2
* cell instance $36915 r0 *1 273.22,222.6
X$36915 5 714 73 85 27 6 DFF_X1
* cell instance $36918 r0 *1 277.02,222.6
X$36918 5 674 49 64 27 6 DFF_X1
* cell instance $36924 r0 *1 286.71,222.6
X$36924 5 680 98 106 42 6 DFF_X1
.ENDS fifo

* cell XOR2_X1
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT XOR2_X1 1 3 4 5 6
* net 1 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 8 1 2 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 7 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 6 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 7 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 2 1 4 4 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 4 3 2 4 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.555,0.2975 NMOS_VTL
M$8 6 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.745,0.2975 NMOS_VTL
M$9 9 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.935,0.2975 NMOS_VTL
M$10 4 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XOR2_X1

* cell NAND2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 6 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 5 2 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X1

* cell XOR2_X2
* pin B
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT XOR2_X2 1 2 4 5 7
* net 1 B
* net 2 A
* net 4 NWELL,VDD
* net 5 Z
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.2,0.995 PMOS_VTL
M$1 8 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.39,0.995 PMOS_VTL
M$2 4 1 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.58,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.77,0.995 PMOS_VTL
M$4 5 2 6 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.96,0.995 PMOS_VTL
M$5 6 1 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.2,0.2975 NMOS_VTL
M$9 3 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.39,0.2975 NMOS_VTL
M$10 7 1 3 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.58,0.2975 NMOS_VTL
M$11 5 3 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $12 r0 *1 0.77,0.2975 NMOS_VTL
M$12 10 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.96,0.2975 NMOS_VTL
M$13 7 1 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.15,0.2975 NMOS_VTL
M$14 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.34,0.2975 NMOS_VTL
M$15 5 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
.ENDS XOR2_X2

* cell INV_X4
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT INV_X4 1 2 3
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 2 2 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
.ENDS INV_X4

* cell NAND2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 4 1 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 5 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND2_X4

* cell NOR3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 6 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 4 2 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR3_X1

* cell NAND2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.195,0.2975 NMOS_VTL
M$5 7 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.385,0.2975 NMOS_VTL
M$6 5 2 7 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.575,0.2975 NMOS_VTL
M$7 6 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.765,0.2975 NMOS_VTL
M$8 3 1 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X2

* cell OAI21_X4
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X4 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 11 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 7 3 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 5 2 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 9 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 7 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 8 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 5 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 6 1 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 7 2 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $18 r0 *1 1.12,0.2975 NMOS_VTL
M$18 4 3 7 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI21_X4

* cell NOR2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 6 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 5 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X1

* cell OR2_X2
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X2 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 3 2 4 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 4 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR2_X2

* cell BUF_X16
* pin PWELL,VSS
* pin A
* pin Z
* pin NWELL,VDD
.SUBCKT BUF_X16 1 2 4 5
* net 1 PWELL,VSS
* net 2 A
* net 4 Z
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 3 2 5 5 PMOS_VTL L=0.05U W=5.04U AS=0.37485P AD=0.3528P PS=6.86U PD=6.16U
* device instance $9 r0 *1 1.705,0.995 PMOS_VTL
M$9 4 3 5 5 PMOS_VTL L=0.05U W=10.08U AS=0.7056P AD=0.72765P PS=12.32U PD=13.02U
* device instance $25 r0 *1 0.185,0.2975 NMOS_VTL
M$25 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.246925P AD=0.2324P PS=4.925U PD=4.44U
* device instance $33 r0 *1 1.705,0.2975 NMOS_VTL
M$33 4 3 1 1 NMOS_VTL L=0.05U W=6.64U AS=0.4648P AD=0.479325P PS=8.88U PD=9.365U
.ENDS BUF_X16

* cell BUF_X8
* pin PWELL,VSS
* pin Z
* pin NWELL,VDD
* pin A
.SUBCKT BUF_X8 1 3 4 5
* net 1 PWELL,VSS
* net 3 Z
* net 4 NWELL,VDD
* net 5 A
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 5 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 4 4 PMOS_VTL L=0.05U W=5.04U AS=0.3528P AD=0.37485P PS=6.16U PD=6.86U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.2324P AD=0.246925P PS=4.44U PD=4.925U
.ENDS BUF_X8

* cell OR2_X1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X1 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 7 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 4 1 3 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 3 2 4 3 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 4 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR2_X1

* cell OAI21_X2
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X2 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 3 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 5 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 6 1 4 6 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 7 2 4 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 4 3 7 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI21_X2

* cell AOI21_X1
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X1 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 2 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 7 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 8 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 6 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 4 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

* cell OR3_X1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 9 1 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 8 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 5 1 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 4 2 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 5 3 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR3_X1

* cell NOR3_X4
* pin PWELL,VSS
* pin A1
* pin A2
* pin A3
* pin ZN
* pin NWELL,VDD
.SUBCKT NOR3_X4 1 2 3 4 5 8
* net 1 PWELL,VSS
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 ZN
* net 8 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 5 2 7 8 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 6 3 7 8 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 1.875,0.995 PMOS_VTL
M$9 6 4 8 8 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $13 r0 *1 1.875,0.2975 NMOS_VTL
M$13 5 4 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $17 r0 *1 0.17,0.2975 NMOS_VTL
M$17 5 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 0.93,0.2975 NMOS_VTL
M$21 5 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NOR3_X4

* cell NOR2_X4
* pin A2
* pin A1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT NOR2_X4 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 ZN
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 9 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 3 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 8 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 1 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 3 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 6 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 1 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 3 1 4 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 4 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS NOR2_X4

* cell NAND4_X4
* pin PWELL,VSS
* pin A3
* pin A4
* pin A1
* pin A2
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND4_X4 1 2 3 7 8 9 10
* net 1 PWELL,VSS
* net 2 A3
* net 3 A4
* net 7 A1
* net 8 A2
* net 9 ZN
* net 10 NWELL,VDD
* device instance $1 r0 *1 0.215,0.995 PMOS_VTL
M$1 10 7 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.975,0.995 PMOS_VTL
M$5 10 8 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.22365P PS=3.08U PD=3.23U
* device instance $9 r0 *1 1.885,0.995 PMOS_VTL
M$9 10 2 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.22365P AD=0.1764P PS=3.23U PD=3.08U
* device instance $13 r0 *1 2.645,0.995 PMOS_VTL
M$13 10 3 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $17 r0 *1 1.885,0.2975 NMOS_VTL
M$17 5 2 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 2.645,0.2975 NMOS_VTL
M$21 1 3 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $25 r0 *1 0.215,0.2975 NMOS_VTL
M$25 9 7 4 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $29 r0 *1 0.975,0.2975 NMOS_VTL
M$29 5 8 4 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND4_X4

* cell XNOR2_X2
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT XNOR2_X2 2 3 4 5 7
* net 2 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 1.135,0.995 PMOS_VTL
M$1 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 1.325,0.995 PMOS_VTL
M$2 9 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 1.515,0.995 PMOS_VTL
M$3 5 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 1.705,0.995 PMOS_VTL
M$4 8 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.18,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $7 r0 *1 0.56,0.995 PMOS_VTL
M$7 1 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 0.75,0.995 PMOS_VTL
M$8 5 2 1 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.135,0.2975 NMOS_VTL
M$9 6 2 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $11 r0 *1 1.515,0.2975 NMOS_VTL
M$11 6 3 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $13 r0 *1 0.18,0.2975 NMOS_VTL
M$13 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $15 r0 *1 0.56,0.2975 NMOS_VTL
M$15 10 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.75,0.2975 NMOS_VTL
M$16 1 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X2

* cell HA_X1
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin CO
.SUBCKT HA_X1 1 2 4 5 6 9
* net 1 A
* net 2 B
* net 4 S
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 9 CO
* device instance $1 r0 *1 0.785,1.0275 PMOS_VTL
M$1 10 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $2 r0 *1 0.975,1.0275 PMOS_VTL
M$2 7 1 10 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $3 r0 *1 0.21,0.995 PMOS_VTL
M$3 4 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $4 r0 *1 0.4,0.995 PMOS_VTL
M$4 3 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.59,0.995 PMOS_VTL
M$5 5 7 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0338625P PS=0.77U PD=0.775U
* device instance $6 r0 *1 1.345,1.0275 PMOS_VTL
M$6 8 1 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $7 r0 *1 1.535,1.0275 PMOS_VTL
M$7 8 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $8 r0 *1 1.725,0.995 PMOS_VTL
M$8 9 8 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.785,0.195 NMOS_VTL
M$9 7 2 6 6 NMOS_VTL L=0.05U W=0.21U AS=0.0224P AD=0.0147P PS=0.56U PD=0.35U
* device instance $10 r0 *1 0.975,0.195 NMOS_VTL
M$10 6 1 7 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $11 r0 *1 0.21,0.2975 NMOS_VTL
M$11 11 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.4,0.2975 NMOS_VTL
M$12 4 1 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.59,0.2975 NMOS_VTL
M$13 6 7 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0224P PS=0.555U PD=0.56U
* device instance $14 r0 *1 1.345,0.195 NMOS_VTL
M$14 12 1 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $15 r0 *1 1.535,0.195 NMOS_VTL
M$15 6 2 12 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $16 r0 *1 1.725,0.2975 NMOS_VTL
M$16 9 8 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS HA_X1

* cell INV_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X1 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P PS=1.47U PD=1.47U
* device instance $2 r0 *1 0.17,0.2975 NMOS_VTL
M$2 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1

* cell CLKBUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.17,0.1875 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $5 r0 *1 0.36,0.1875 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.39U AS=0.0273P AD=0.034125P PS=0.67U PD=0.935U
.ENDS CLKBUF_X2

* cell BUF_X4
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT BUF_X4 1 3 4 5
* net 1 A
* net 3 NWELL,VDD
* net 4 Z
* net 5 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 2 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 4 2 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS BUF_X4

* cell CLKBUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT CLKBUF_X1 1 3 4
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.19,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.38,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.19,0.2075 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.095U AS=0.009975P AD=0.01015P PS=0.4U PD=0.335U
* device instance $4 r0 *1 0.38,0.2575 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01015P AD=0.020475P PS=0.335U PD=0.6U
.ENDS CLKBUF_X1

* cell AOI22_X1
* pin B2
* pin B1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AOI22_X1 1 2 3 4 5 7 8
* net 1 B2
* net 2 B1
* net 3 A1
* net 4 A2
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 7 1 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 6 2 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 8 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 6 4 8 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.185,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.375,0.2975 NMOS_VTL
M$6 8 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.565,0.2975 NMOS_VTL
M$7 9 3 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.755,0.2975 NMOS_VTL
M$8 5 4 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI22_X1

* cell BUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS BUF_X2

* cell AND2_X1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X1 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 7 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 5 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND2_X1

* cell NAND3_X4
* pin A2
* pin A1
* pin A3
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND3_X4 1 2 3 4 5 6
* net 1 A2
* net 2 A1
* net 3 A3
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 3 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 6 1 5 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $13 r0 *1 0.21,0.2975 NMOS_VTL
M$13 13 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $14 r0 *1 0.4,0.2975 NMOS_VTL
M$14 12 1 13 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.59,0.2975 NMOS_VTL
M$15 5 2 12 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.78,0.2975 NMOS_VTL
M$16 10 2 5 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 0.97,0.2975 NMOS_VTL
M$17 8 1 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.16,0.2975 NMOS_VTL
M$18 4 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.35,0.2975 NMOS_VTL
M$19 9 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.54,0.2975 NMOS_VTL
M$20 7 1 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.73,0.2975 NMOS_VTL
M$21 5 2 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.92,0.2975 NMOS_VTL
M$22 14 2 5 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.11,0.2975 NMOS_VTL
M$23 11 1 14 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.3,0.2975 NMOS_VTL
M$24 4 3 11 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X4

* cell INV_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X2 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 4 1 2 2 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
.ENDS INV_X2

* cell BUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.17,0.195 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U PD=0.555U
* device instance $4 r0 *1 0.36,0.2975 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X1

* cell DFF_X1
* pin PWELL,VSS
* pin QN
* pin Q
* pin D
* pin CK
* pin NWELL,VDD
.SUBCKT DFF_X1 1 8 9 14 15 16
* net 1 PWELL,VSS
* net 8 QN
* net 9 Q
* net 14 D
* net 15 CK
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.85,0.995 PMOS_VTL
M$1 16 6 8 16 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 3.04,0.995 PMOS_VTL
M$2 9 7 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.9425 PMOS_VTL
M$3 16 5 2 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $4 r0 *1 0.375,1.055 PMOS_VTL
M$4 17 3 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $5 r0 *1 0.565,1.055 PMOS_VTL
M$5 17 5 4 16 PMOS_VTL L=0.05U W=0.09U AS=0.018075P AD=0.0063P PS=0.565U
+ PD=0.23U
* device instance $6 r0 *1 0.76,0.975 PMOS_VTL
M$6 18 2 4 16 PMOS_VTL L=0.05U W=0.42U AS=0.018075P AD=0.0294P PS=0.565U
+ PD=0.56U
* device instance $7 r0 *1 0.95,0.975 PMOS_VTL
M$7 16 14 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $8 r0 *1 1.14,1.0275 PMOS_VTL
M$8 3 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $9 r0 *1 1.555,1.0275 PMOS_VTL
M$9 16 15 5 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $10 r0 *1 1.745,1.0275 PMOS_VTL
M$10 19 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $11 r0 *1 1.935,1.0275 PMOS_VTL
M$11 6 5 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $12 r0 *1 2.125,1.14 PMOS_VTL
M$12 20 2 6 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $13 r0 *1 2.32,1.14 PMOS_VTL
M$13 20 7 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $14 r0 *1 2.51,1.0275 PMOS_VTL
M$14 7 6 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.014175P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $15 r0 *1 2.85,0.2975 NMOS_VTL
M$15 1 6 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $16 r0 *1 3.04,0.2975 NMOS_VTL
M$16 9 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $17 r0 *1 0.185,0.285 NMOS_VTL
M$17 1 5 2 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $18 r0 *1 0.375,0.345 NMOS_VTL
M$18 10 3 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $19 r0 *1 0.565,0.345 NMOS_VTL
M$19 10 2 4 1 NMOS_VTL L=0.05U W=0.09U AS=0.013P AD=0.0063P PS=0.42U PD=0.23U
* device instance $20 r0 *1 1.14,0.285 NMOS_VTL
M$20 3 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $21 r0 *1 0.76,0.3175 NMOS_VTL
M$21 11 5 4 1 NMOS_VTL L=0.05U W=0.275U AS=0.013P AD=0.01925P PS=0.42U PD=0.415U
* device instance $22 r0 *1 0.95,0.3175 NMOS_VTL
M$22 1 14 11 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
* device instance $23 r0 *1 2.125,0.345 NMOS_VTL
M$23 12 5 6 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $24 r0 *1 2.32,0.345 NMOS_VTL
M$24 12 7 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $25 r0 *1 1.555,0.36 NMOS_VTL
M$25 1 15 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $26 r0 *1 1.745,0.36 NMOS_VTL
M$26 13 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 1.935,0.36 NMOS_VTL
M$27 6 2 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $28 r0 *1 2.51,0.36 NMOS_VTL
M$28 7 6 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0105P AD=0.02205P PS=0.35U PD=0.63U
.ENDS DFF_X1

* cell DFF_X2
* pin PWELL,VSS
* pin D
* pin CK
* pin QN
* pin Q
* pin NWELL,VDD
.SUBCKT DFF_X2 1 6 8 10 11 16
* net 1 PWELL,VSS
* net 6 D
* net 8 CK
* net 10 QN
* net 11 Q
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.855,0.995 PMOS_VTL
M$1 10 9 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 3.235,0.995 PMOS_VTL
M$3 11 2 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.2,0.9275 PMOS_VTL
M$5 16 7 3 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $6 r0 *1 0.39,1.04 PMOS_VTL
M$6 17 4 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $7 r0 *1 0.58,1.04 PMOS_VTL
M$7 17 7 5 16 PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P PS=0.56U PD=0.23U
* device instance $8 r0 *1 0.77,0.975 PMOS_VTL
M$8 18 3 5 16 PMOS_VTL L=0.05U W=0.42U AS=0.01785P AD=0.0294P PS=0.56U PD=0.56U
* device instance $9 r0 *1 0.96,0.975 PMOS_VTL
M$9 16 6 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $10 r0 *1 1.15,1.0275 PMOS_VTL
M$10 4 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $11 r0 *1 2.135,0.915 PMOS_VTL
M$11 20 3 9 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $12 r0 *1 2.325,0.915 PMOS_VTL
M$12 20 2 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.0252P AD=0.0063P PS=0.77U PD=0.23U
* device instance $13 r0 *1 1.565,1.0275 PMOS_VTL
M$13 16 8 7 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $14 r0 *1 1.755,1.0275 PMOS_VTL
M$14 19 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $15 r0 *1 1.945,1.0275 PMOS_VTL
M$15 9 7 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $16 r0 *1 2.515,0.995 PMOS_VTL
M$16 2 9 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0252P AD=0.06615P PS=0.77U PD=1.47U
* device instance $17 r0 *1 2.855,0.2975 NMOS_VTL
M$17 10 9 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U
+ PD=1.11U
* device instance $19 r0 *1 3.235,0.2975 NMOS_VTL
M$19 11 2 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U
+ PD=1.595U
* device instance $21 r0 *1 0.39,0.31 NMOS_VTL
M$21 12 4 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $22 r0 *1 0.58,0.31 NMOS_VTL
M$22 12 3 5 1 NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P PS=0.415U
+ PD=0.23U
* device instance $23 r0 *1 1.15,0.25 NMOS_VTL
M$23 4 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $24 r0 *1 0.77,0.2825 NMOS_VTL
M$24 13 7 5 1 NMOS_VTL L=0.05U W=0.275U AS=0.012775P AD=0.01925P PS=0.415U
+ PD=0.415U
* device instance $25 r0 *1 0.96,0.2825 NMOS_VTL
M$25 1 6 13 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
* device instance $26 r0 *1 0.2,0.37 NMOS_VTL
M$26 1 7 3 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $27 r0 *1 1.565,0.35 NMOS_VTL
M$27 1 8 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $28 r0 *1 1.755,0.35 NMOS_VTL
M$28 14 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $29 r0 *1 1.945,0.35 NMOS_VTL
M$29 9 3 14 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $30 r0 *1 2.135,0.41 NMOS_VTL
M$30 15 7 9 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $31 r0 *1 2.325,0.41 NMOS_VTL
M$31 15 2 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.017675P AD=0.0063P PS=0.555U
+ PD=0.23U
* device instance $32 r0 *1 2.515,0.2975 NMOS_VTL
M$32 2 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.017675P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS DFF_X2

* cell OAI21_X1
* pin B2
* pin B1
* pin A
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OAI21_X1 1 2 3 5 6 7
* net 1 B2
* net 2 B1
* net 3 A
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 6 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.195,0.2975 NMOS_VTL
M$4 6 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.385,0.2975 NMOS_VTL
M$5 4 2 6 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.575,0.2975 NMOS_VTL
M$6 7 3 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X1

* cell NAND3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 8 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X1

* cell MUX2_X1
* pin A
* pin S
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT MUX2_X1 1 2 3 5 6 8
* net 1 A
* net 2 S
* net 3 B
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 8 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 6 2 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 7 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 10 4 7 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $5 r0 *1 0.93,1.1525 PMOS_VTL
M$5 10 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 7 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.195 NMOS_VTL
M$7 5 2 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $8 r0 *1 0.36,0.195 NMOS_VTL
M$8 12 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.55,0.195 NMOS_VTL
M$9 7 4 12 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $10 r0 *1 0.74,0.195 NMOS_VTL
M$10 11 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $11 r0 *1 0.93,0.195 NMOS_VTL
M$11 5 3 11 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 7 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS MUX2_X1

* cell CLKBUF_X3
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X3 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.89U AS=0.1323P AD=0.15435P PS=2.31U PD=3.01U
* device instance $5 r0 *1 0.17,0.1875 NMOS_VTL
M$5 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $6 r0 *1 0.36,0.1875 NMOS_VTL
M$6 5 2 3 3 NMOS_VTL L=0.05U W=0.585U AS=0.04095P AD=0.047775P PS=1.005U
+ PD=1.27U
.ENDS CLKBUF_X3
