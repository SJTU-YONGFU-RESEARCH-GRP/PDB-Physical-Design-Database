module fixed_point_sqrt (clk,
    enable,
    reset,
    x,
    y);
 input clk;
 input enable;
 input reset;
 input [15:0] x;
 output [15:0] y;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _111_ (.A1(net7),
    .A2(net6),
    .A3(net8),
    .A4(net9),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _112_ (.A1(net20),
    .A2(net1),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _113_ (.A1(net1),
    .A2(_051_),
    .B(_052_),
    .C(net2),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _114_ (.I(net1),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _115_ (.I(net17),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _116_ (.A1(net11),
    .A2(net14),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _117_ (.A1(net3),
    .A2(net12),
    .A3(net13),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _118_ (.A1(net16),
    .A2(net15),
    .A3(net18),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _119_ (.A1(net10),
    .A2(_055_),
    .A3(_056_),
    .A4(_057_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _120_ (.A1(net4),
    .A2(net5),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _121_ (.A1(_051_),
    .A2(_059_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _122_ (.A1(_054_),
    .A2(_058_),
    .A3(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _123_ (.A1(net1),
    .A2(_061_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _124_ (.A1(net10),
    .A2(_055_),
    .A3(_056_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _125_ (.A1(_051_),
    .A2(_059_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _126_ (.A1(net16),
    .A2(net18),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _127_ (.A1(net15),
    .A2(net17),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _128_ (.A1(_063_),
    .A2(_064_),
    .A3(_065_),
    .A4(_066_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _129_ (.A1(net13),
    .A2(net6),
    .A3(net8),
    .A4(net9),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _130_ (.A1(net17),
    .A2(net4),
    .A3(net5),
    .A4(net7),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _131_ (.A1(net3),
    .A2(net10),
    .A3(net12),
    .A4(net15),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _132_ (.A1(net11),
    .A2(net14),
    .A3(_065_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _133_ (.A1(_068_),
    .A2(_069_),
    .A3(_070_),
    .A4(_071_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _134_ (.A1(_067_),
    .A2(_072_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _135_ (.I(_073_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _136_ (.A1(_053_),
    .A2(net22),
    .B1(_062_),
    .B2(_074_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _137_ (.A1(net2),
    .A2(_075_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _138_ (.A1(_053_),
    .A2(net21),
    .B1(_062_),
    .B2(_072_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _139_ (.A1(net2),
    .A2(_076_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _140_ (.A1(net3),
    .A2(net12),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _141_ (.I(net18),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _142_ (.A1(_078_),
    .A2(_054_),
    .A3(_051_),
    .A4(_059_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _143_ (.A1(net10),
    .A2(net16),
    .A3(net15),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _144_ (.A1(_055_),
    .A2(_077_),
    .A3(_079_),
    .A4(_080_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _145_ (.A1(_073_),
    .A2(_081_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _146_ (.A1(_053_),
    .A2(net25),
    .B1(_062_),
    .B2(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _147_ (.A1(net2),
    .A2(_083_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _148_ (.A1(net1),
    .A2(_061_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _149_ (.A1(net2),
    .A2(_084_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _150_ (.A1(net16),
    .A2(net15),
    .A3(_079_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _151_ (.A1(_054_),
    .A2(net6),
    .A3(_059_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _152_ (.I(net4),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _153_ (.A1(net17),
    .A2(_088_),
    .A3(net5),
    .A4(net6),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _154_ (.A1(_087_),
    .A2(_089_),
    .B(net7),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _155_ (.I(net5),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _156_ (.A1(net4),
    .A2(_091_),
    .A3(net7),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _157_ (.A1(net4),
    .A2(_091_),
    .A3(net7),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _158_ (.I(net6),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _159_ (.A1(net17),
    .A2(_094_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _160_ (.A1(_092_),
    .A2(_093_),
    .B(_095_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _161_ (.A1(net8),
    .A2(net9),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _162_ (.A1(_097_),
    .A2(_058_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _163_ (.A1(_090_),
    .A2(_096_),
    .B(_098_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _164_ (.A1(net3),
    .A2(net12),
    .Z(_100_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _165_ (.I(net13),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _166_ (.A1(net12),
    .A2(_101_),
    .B(net3),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _167_ (.A1(_100_),
    .A2(_102_),
    .B(_055_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _168_ (.I(net12),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _169_ (.A1(_104_),
    .A2(net11),
    .A3(net14),
    .A4(_101_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _170_ (.A1(net3),
    .A2(_105_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _171_ (.A1(net14),
    .A2(_056_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _172_ (.A1(_079_),
    .A2(_080_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _173_ (.A1(_103_),
    .A2(_106_),
    .A3(_107_),
    .B(_108_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _174_ (.A1(net11),
    .A2(net14),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _175_ (.A1(net10),
    .A2(net16),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _176_ (.A1(net15),
    .A2(_010_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _177_ (.A1(_056_),
    .A2(_079_),
    .A3(_009_),
    .A4(_011_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _178_ (.A1(_099_),
    .A2(_109_),
    .A3(_012_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _179_ (.I(_013_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _180_ (.A1(net1),
    .A2(net2),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _181_ (.A1(net2),
    .A2(_084_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _182_ (.A1(net3),
    .A2(net15),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _183_ (.A1(_105_),
    .A2(_010_),
    .A3(_017_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _184_ (.I0(_077_),
    .I1(_100_),
    .S(net11),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _185_ (.A1(net14),
    .A2(net13),
    .A3(_080_),
    .A4(_019_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _186_ (.A1(_018_),
    .A2(_020_),
    .B(_079_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _187_ (.A1(_072_),
    .A2(_021_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _188_ (.A1(net26),
    .A2(_015_),
    .B1(_016_),
    .B2(_022_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _189_ (.A1(_085_),
    .A2(_086_),
    .A3(_014_),
    .B(_023_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _190_ (.A1(_073_),
    .A2(_079_),
    .A3(_099_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _191_ (.I(_067_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _192_ (.A1(_104_),
    .A2(_101_),
    .A3(_055_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _193_ (.A1(_105_),
    .A2(_026_),
    .B(net3),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _194_ (.A1(_101_),
    .A2(_055_),
    .A3(_100_),
    .B(_027_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _195_ (.A1(_025_),
    .A2(_013_),
    .B1(_028_),
    .B2(_108_),
    .C(_072_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _196_ (.A1(net27),
    .A2(_015_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _197_ (.A1(_085_),
    .A2(_024_),
    .A3(_029_),
    .B(_030_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _198_ (.A1(net18),
    .A2(net17),
    .B(net4),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _199_ (.A1(_091_),
    .A2(_094_),
    .A3(_031_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _200_ (.A1(net7),
    .A2(_032_),
    .B(_097_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _201_ (.A1(_086_),
    .A2(_099_),
    .A3(_033_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _202_ (.A1(_073_),
    .A2(_012_),
    .A3(_034_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _203_ (.A1(net28),
    .A2(_015_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _204_ (.A1(_085_),
    .A2(_035_),
    .B(_036_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _205_ (.A1(net4),
    .A2(net7),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _206_ (.A1(_092_),
    .A2(_037_),
    .B(_095_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _207_ (.A1(_098_),
    .A2(_038_),
    .B(_053_),
    .C(_074_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _208_ (.A1(net4),
    .A2(_091_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _209_ (.A1(net18),
    .A2(net17),
    .A3(net4),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _210_ (.A1(_051_),
    .A2(_040_),
    .A3(_013_),
    .A4(_041_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _211_ (.A1(net1),
    .A2(net29),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _212_ (.A1(_039_),
    .A2(_042_),
    .B(_043_),
    .C(net2),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _213_ (.A1(net7),
    .A2(net6),
    .A3(_097_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _214_ (.A1(_044_),
    .A2(_033_),
    .B(_072_),
    .C(_064_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _215_ (.A1(_088_),
    .A2(net5),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _216_ (.I0(_040_),
    .I1(_046_),
    .S(net17),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _217_ (.A1(_044_),
    .A2(_058_),
    .A3(_047_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _218_ (.A1(_013_),
    .A2(_045_),
    .B(_048_),
    .C(_072_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _219_ (.A1(net30),
    .A2(_015_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _220_ (.A1(_085_),
    .A2(_049_),
    .B(_050_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _222_ (.I(net21),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _223_ (.I(net21),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _224_ (.I(net21),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _225_ (.I(net31),
    .Z(y[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _226_ (.I(net32),
    .Z(y[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _227_ (.I(net33),
    .Z(y[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _228_ (.I(net34),
    .Z(y[15]));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[10]$_SDFFE_PP0P_  (.D(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[1]$_SDFFE_PP0P_  (.D(_001_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[3]$_SDFFE_PP0P_  (.D(_002_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[4]$_SDFFE_PP0P_  (.D(_003_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[5]$_SDFFE_PP0P_  (.D(_004_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[6]$_SDFFE_PP0P_  (.D(_005_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[7]$_SDFFE_PP0P_  (.D(_006_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[8]$_SDFFE_PP0P_  (.D(_007_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \y[9]$_SDFFE_PP0P_  (.D(_008_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_70 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_72 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_73 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_74 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_75 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_76 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_77 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_78 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_79 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_80 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_81 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_82 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_83 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_84 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_87 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input1 (.I(enable),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input2 (.I(reset),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input3 (.I(x[0]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input4 (.I(x[10]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input5 (.I(x[11]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input6 (.I(x[12]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input7 (.I(x[13]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(x[14]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(x[15]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input10 (.I(x[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input11 (.I(x[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(x[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(x[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input14 (.I(x[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input15 (.I(x[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input16 (.I(x[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input17 (.I(x[8]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input18 (.I(x[9]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net19),
    .Z(y[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net20),
    .Z(y[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net21),
    .Z(y[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net22),
    .Z(y[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net23),
    .Z(y[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net24),
    .Z(y[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output25 (.I(net25),
    .Z(y[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output26 (.I(net26),
    .Z(y[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output27 (.I(net27),
    .Z(y[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output28 (.I(net28),
    .Z(y[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output29 (.I(net29),
    .Z(y[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output30 (.I(net30),
    .Z(y[9]));
 gf180mcu_fd_sc_mcu9t5v0__tiel _225__31 (.ZN(net31));
 gf180mcu_fd_sc_mcu9t5v0__tiel _226__32 (.ZN(net32));
 gf180mcu_fd_sc_mcu9t5v0__tiel _227__33 (.ZN(net33));
 gf180mcu_fd_sc_mcu9t5v0__tiel _228__34 (.ZN(net34));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_327 ();
endmodule
