module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire net3149;
 wire net3148;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire net3155;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire net3143;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire net3142;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire net3147;
 wire _02016_;
 wire _02017_;
 wire net3157;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire clknet_leaf_127_clk_i_regs;
 wire _02042_;
 wire _02043_;
 wire net3141;
 wire _02045_;
 wire _02046_;
 wire net3516;
 wire _02048_;
 wire net3139;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire net3160;
 wire net3138;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire clknet_leaf_128_clk_i_regs;
 wire _02156_;
 wire _02157_;
 wire clknet_leaf_129_clk_i_regs;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire clknet_leaf_134_clk_i_regs;
 wire clknet_leaf_136_clk_i_regs;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire clknet_leaf_137_clk_i_regs;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire clknet_leaf_138_clk_i_regs;
 wire clknet_leaf_139_clk_i_regs;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire clknet_leaf_141_clk_i_regs;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire clknet_leaf_142_clk_i_regs;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire clknet_leaf_143_clk_i_regs;
 wire _02410_;
 wire clknet_leaf_145_clk_i_regs;
 wire _02412_;
 wire net3554;
 wire net3515;
 wire _02415_;
 wire _02416_;
 wire clknet_leaf_147_clk_i_regs;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire net3128;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire net3553;
 wire _02446_;
 wire clknet_leaf_149_clk_i_regs;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire net3129;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire net3127;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire net3642;
 wire _02480_;
 wire net3126;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire net3131;
 wire _02517_;
 wire net3123;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire net3561;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire net3125;
 wire net3121;
 wire net3117;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire net3118;
 wire _02537_;
 wire _02538_;
 wire net3116;
 wire net3119;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire net3114;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire net3115;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire clknet_leaf_151_clk_i_regs;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire clknet_leaf_154_clk_i_regs;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire net3113;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire net3566;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire net3641;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire net3109;
 wire net3640;
 wire _02618_;
 wire _02619_;
 wire net3108;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire net3565;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire clknet_leaf_156_clk_i_regs;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire clknet_leaf_158_clk_i_regs;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire net3107;
 wire clknet_leaf_162_clk_i_regs;
 wire clknet_leaf_160_clk_i_regs;
 wire _02673_;
 wire clknet_leaf_165_clk_i_regs;
 wire clknet_leaf_166_clk_i_regs;
 wire net3106;
 wire net3105;
 wire _02678_;
 wire net3564;
 wire clknet_leaf_167_clk_i_regs;
 wire _02681_;
 wire clknet_leaf_169_clk_i_regs;
 wire clknet_leaf_171_clk_i_regs;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire clknet_leaf_174_clk_i_regs;
 wire clknet_leaf_177_clk_i_regs;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire clknet_leaf_178_clk_i_regs;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire clknet_leaf_179_clk_i_regs;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire clknet_leaf_180_clk_i_regs;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire net3103;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire clknet_leaf_182_clk_i_regs;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire clknet_leaf_185_clk_i_regs;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire clknet_leaf_183_clk_i_regs;
 wire clknet_leaf_186_clk_i_regs;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire clknet_leaf_187_clk_i_regs;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire clknet_leaf_188_clk_i_regs;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire clknet_leaf_191_clk_i_regs;
 wire net3563;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire clknet_leaf_193_clk_i_regs;
 wire _02872_;
 wire clknet_leaf_196_clk_i_regs;
 wire _02874_;
 wire _02875_;
 wire clknet_leaf_197_clk_i_regs;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire clknet_leaf_198_clk_i_regs;
 wire clknet_leaf_200_clk_i_regs;
 wire clknet_leaf_201_clk_i_regs;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire clknet_leaf_202_clk_i_regs;
 wire _02905_;
 wire _02906_;
 wire clknet_leaf_205_clk_i_regs;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire clknet_leaf_207_clk_i_regs;
 wire clknet_leaf_208_clk_i_regs;
 wire clknet_leaf_211_clk_i_regs;
 wire _02926_;
 wire _02927_;
 wire clknet_leaf_214_clk_i_regs;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire clknet_leaf_215_clk_i_regs;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire clknet_leaf_217_clk_i_regs;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire net3562;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire clknet_leaf_219_clk_i_regs;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire net3104;
 wire net3639;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire clknet_leaf_222_clk_i_regs;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire clknet_leaf_226_clk_i_regs;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire clknet_leaf_229_clk_i_regs;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire clknet_leaf_230_clk_i_regs;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire clknet_leaf_231_clk_i_regs;
 wire _03018_;
 wire _03019_;
 wire clknet_leaf_233_clk_i_regs;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire clknet_leaf_234_clk_i_regs;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire net3638;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire clknet_leaf_235_clk_i_regs;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire clknet_leaf_237_clk_i_regs;
 wire _03078_;
 wire _03079_;
 wire clknet_leaf_238_clk_i_regs;
 wire clknet_leaf_241_clk_i_regs;
 wire clknet_leaf_242_clk_i_regs;
 wire clknet_leaf_244_clk_i_regs;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire clknet_leaf_247_clk_i_regs;
 wire clknet_leaf_248_clk_i_regs;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire clknet_leaf_250_clk_i_regs;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire clknet_leaf_251_clk_i_regs;
 wire _03106_;
 wire _03107_;
 wire net3098;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire net3097;
 wire _03113_;
 wire _03114_;
 wire clknet_leaf_252_clk_i_regs;
 wire _03116_;
 wire clknet_leaf_254_clk_i_regs;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire clknet_leaf_255_clk_i_regs;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire clknet_leaf_256_clk_i_regs;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire clknet_leaf_258_clk_i_regs;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire clknet_leaf_260_clk_i_regs;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire clknet_leaf_262_clk_i_regs;
 wire _03154_;
 wire clknet_leaf_263_clk_i_regs;
 wire _03156_;
 wire clknet_leaf_264_clk_i_regs;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire clknet_leaf_265_clk_i_regs;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire clknet_leaf_266_clk_i_regs;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire clknet_leaf_269_clk_i_regs;
 wire net3096;
 wire _03221_;
 wire clknet_leaf_276_clk_i_regs;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire clknet_leaf_277_clk_i_regs;
 wire clknet_leaf_278_clk_i_regs;
 wire clknet_leaf_280_clk_i_regs;
 wire clknet_leaf_281_clk_i_regs;
 wire _03237_;
 wire clknet_leaf_283_clk_i_regs;
 wire _03239_;
 wire _03240_;
 wire clknet_leaf_282_clk_i_regs;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire clknet_leaf_284_clk_i_regs;
 wire clknet_leaf_285_clk_i_regs;
 wire _03248_;
 wire clknet_leaf_286_clk_i_regs;
 wire clknet_leaf_287_clk_i_regs;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire clknet_leaf_288_clk_i_regs;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire clknet_leaf_289_clk_i_regs;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire clknet_leaf_294_clk_i_regs;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire clknet_leaf_292_clk_i_regs;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire clknet_leaf_295_clk_i_regs;
 wire _03298_;
 wire clknet_leaf_296_clk_i_regs;
 wire _03300_;
 wire clknet_leaf_297_clk_i_regs;
 wire clknet_leaf_304_clk_i_regs;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire clknet_leaf_299_clk_i_regs;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire clknet_leaf_303_clk_i_regs;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire clknet_leaf_301_clk_i_regs;
 wire clknet_leaf_302_clk_i_regs;
 wire clknet_leaf_306_clk_i_regs;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire clknet_leaf_307_clk_i_regs;
 wire clknet_leaf_308_clk_i_regs;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire clknet_leaf_309_clk_i_regs;
 wire _03359_;
 wire _03360_;
 wire clknet_leaf_310_clk_i_regs;
 wire clknet_leaf_311_clk_i_regs;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire clknet_leaf_312_clk_i_regs;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire clknet_leaf_317_clk_i_regs;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire clknet_leaf_319_clk_i_regs;
 wire clknet_leaf_320_clk_i_regs;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire clknet_leaf_322_clk_i_regs;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire clknet_leaf_324_clk_i_regs;
 wire _03441_;
 wire _03442_;
 wire net3094;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire clknet_leaf_325_clk_i_regs;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire clknet_leaf_330_clk_i_regs;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire clknet_leaf_327_clk_i_regs;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire clknet_leaf_332_clk_i_regs;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire clknet_leaf_331_clk_i_regs;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire clknet_leaf_334_clk_i_regs;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire clknet_leaf_335_clk_i_regs;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire clknet_leaf_338_clk_i_regs;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire clknet_leaf_339_clk_i_regs;
 wire _03566_;
 wire _03567_;
 wire clknet_leaf_342_clk_i_regs;
 wire net3093;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire clknet_leaf_343_clk_i_regs;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire clknet_leaf_347_clk_i_regs;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire clknet_leaf_348_clk_i_regs;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire clknet_leaf_349_clk_i_regs;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire clknet_leaf_350_clk_i_regs;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire clknet_leaf_352_clk_i_regs;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire clknet_leaf_356_clk_i_regs;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire clknet_leaf_359_clk_i_regs;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire clknet_leaf_360_clk_i_regs;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire clknet_leaf_361_clk_i_regs;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire clknet_leaf_364_clk_i_regs;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire clknet_leaf_365_clk_i_regs;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire clknet_leaf_368_clk_i_regs;
 wire clknet_leaf_371_clk_i_regs;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire clknet_leaf_373_clk_i_regs;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire clknet_leaf_375_clk_i_regs;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire clknet_leaf_376_clk_i_regs;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire clknet_leaf_378_clk_i_regs;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire clknet_leaf_379_clk_i_regs;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire clknet_leaf_380_clk_i_regs;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire clknet_leaf_381_clk_i_regs;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire clknet_leaf_385_clk_i_regs;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire clknet_leaf_384_clk_i_regs;
 wire clknet_leaf_383_clk_i_regs;
 wire net3090;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire clknet_leaf_393_clk_i_regs;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire clknet_leaf_389_clk_i_regs;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire clknet_leaf_386_clk_i_regs;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire clknet_leaf_391_clk_i_regs;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire clknet_leaf_398_clk_i_regs;
 wire clknet_leaf_396_clk_i_regs;
 wire net3088;
 wire clknet_leaf_397_clk_i_regs;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire net3086;
 wire _04117_;
 wire net3085;
 wire net3084;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire net3082;
 wire _04124_;
 wire clknet_leaf_408_clk_i_regs;
 wire clknet_leaf_407_clk_i_regs;
 wire _04127_;
 wire clknet_leaf_405_clk_i_regs;
 wire _04129_;
 wire clknet_leaf_404_clk_i_regs;
 wire clknet_leaf_403_clk_i_regs;
 wire _04132_;
 wire _04133_;
 wire clknet_leaf_402_clk_i_regs;
 wire _04135_;
 wire clknet_leaf_400_clk_i_regs;
 wire clknet_leaf_399_clk_i_regs;
 wire _04138_;
 wire net3081;
 wire _04140_;
 wire clknet_leaf_412_clk_i_regs;
 wire clknet_leaf_409_clk_i_regs;
 wire _04143_;
 wire clknet_leaf_417_clk_i_regs;
 wire _04145_;
 wire clknet_leaf_416_clk_i_regs;
 wire _04147_;
 wire clknet_leaf_418_clk_i_regs;
 wire _04149_;
 wire net3637;
 wire _04151_;
 wire net3080;
 wire _04153_;
 wire net3079;
 wire clknet_leaf_419_clk_i_regs;
 wire _04156_;
 wire clknet_leaf_428_clk_i_regs;
 wire _04158_;
 wire clknet_leaf_427_clk_i_regs;
 wire clknet_leaf_426_clk_i_regs;
 wire clknet_leaf_424_clk_i_regs;
 wire clknet_leaf_423_clk_i_regs;
 wire clknet_leaf_422_clk_i_regs;
 wire clknet_leaf_420_clk_i_regs;
 wire net3074;
 wire clknet_leaf_430_clk_i_regs;
 wire clknet_leaf_433_clk_i_regs;
 wire clknet_leaf_431_clk_i_regs;
 wire net3076;
 wire clknet_leaf_453_clk_i_regs;
 wire clknet_leaf_450_clk_i_regs;
 wire clknet_leaf_449_clk_i_regs;
 wire clknet_leaf_447_clk_i_regs;
 wire clknet_leaf_446_clk_i_regs;
 wire clknet_leaf_443_clk_i_regs;
 wire clknet_leaf_442_clk_i_regs;
 wire clknet_leaf_440_clk_i_regs;
 wire clknet_leaf_436_clk_i_regs;
 wire clknet_leaf_435_clk_i_regs;
 wire net3101;
 wire clknet_leaf_456_clk_i_regs;
 wire net3102;
 wire net3077;
 wire net3071;
 wire clknet_leaf_462_clk_i_regs;
 wire net3067;
 wire net3066;
 wire clknet_leaf_465_clk_i_regs;
 wire _04189_;
 wire net3065;
 wire _04191_;
 wire net3062;
 wire clknet_leaf_466_clk_i_regs;
 wire net3060;
 wire net3058;
 wire net3057;
 wire net3056;
 wire net3055;
 wire _04199_;
 wire net3054;
 wire _04201_;
 wire net3053;
 wire clknet_leaf_467_clk_i_regs;
 wire _04204_;
 wire net3052;
 wire _04206_;
 wire net3670;
 wire net3653;
 wire _04209_;
 wire _04210_;
 wire net252;
 wire _04212_;
 wire net3652;
 wire net3651;
 wire net3089;
 wire _04216_;
 wire net3636;
 wire _04218_;
 wire net3444;
 wire clknet_leaf_15_clk_i_regs;
 wire _04221_;
 wire clknet_leaf_13_clk_i_regs;
 wire _04223_;
 wire clknet_leaf_39_clk_i_regs;
 wire net3443;
 wire _04226_;
 wire net3665;
 wire _04228_;
 wire net3584;
 wire net3442;
 wire _04231_;
 wire _04232_;
 wire clknet_leaf_90_clk_i_regs;
 wire _04234_;
 wire net3235;
 wire _04236_;
 wire clknet_leaf_38_clk_i_regs;
 wire _04238_;
 wire net3215;
 wire _04240_;
 wire net3612;
 wire _04242_;
 wire _04271_;
 wire _04273_;
 wire _04281_;
 wire _04283_;
 wire _04287_;
 wire _04288_;
 wire _04290_;
 wire _04293_;
 wire _04295_;
 wire _04298_;
 wire _04300_;
 wire _04304_;
 wire _04306_;
 wire _04309_;
 wire _04311_;
 wire _04314_;
 wire _04316_;
 wire _04319_;
 wire _04321_;
 wire _04323_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04406_;
 wire _04407_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04426_;
 wire _04427_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04457_;
 wire _04459_;
 wire _04460_;
 wire _04462_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04487_;
 wire _04488_;
 wire _04490_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04803_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire net149;
 wire _05087_;
 wire net148;
 wire net147;
 wire net146;
 wire net145;
 wire _05092_;
 wire net144;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire net143;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire net142;
 wire net141;
 wire net140;
 wire _05105_;
 wire net139;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire net138;
 wire net137;
 wire _05112_;
 wire net136;
 wire _05114_;
 wire _05115_;
 wire net135;
 wire net134;
 wire _05118_;
 wire net133;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire net132;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire net131;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire net130;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire net129;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire net128;
 wire net127;
 wire net126;
 wire _05266_;
 wire net125;
 wire net124;
 wire _05269_;
 wire _05270_;
 wire net123;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire net122;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire net121;
 wire _05324_;
 wire net120;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire net119;
 wire net118;
 wire _05333_;
 wire net117;
 wire net116;
 wire _05336_;
 wire net115;
 wire _05338_;
 wire _05339_;
 wire net114;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire net113;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire net112;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire net111;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire net110;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire net109;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire net108;
 wire _05468_;
 wire _05469_;
 wire net107;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire net106;
 wire _05488_;
 wire _05489_;
 wire net105;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire net104;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire net103;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire net102;
 wire _05546_;
 wire _05547_;
 wire net101;
 wire net100;
 wire net99;
 wire _05551_;
 wire net98;
 wire net97;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire net96;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire net95;
 wire net94;
 wire net93;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire net92;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire net91;
 wire net90;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire net89;
 wire _05611_;
 wire net88;
 wire net87;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire net86;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire net85;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire net84;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire net83;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire net82;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire net81;
 wire _05675_;
 wire _05676_;
 wire net80;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire net79;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire net78;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire net77;
 wire net76;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire net75;
 wire _05702_;
 wire net74;
 wire _05704_;
 wire _05705_;
 wire net73;
 wire _05707_;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire _05713_;
 wire _05714_;
 wire net67;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire net66;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire net65;
 wire _05730_;
 wire net64;
 wire _05732_;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire _05741_;
 wire _05742_;
 wire net55;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire net54;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire net53;
 wire _05762_;
 wire _05763_;
 wire net52;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire net51;
 wire _05772_;
 wire _05773_;
 wire net50;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire net49;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire net48;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire net47;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire net46;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire net45;
 wire net44;
 wire net43;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire net42;
 wire net41;
 wire _06096_;
 wire net40;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire net39;
 wire _06108_;
 wire _06109_;
 wire net38;
 wire net37;
 wire _06112_;
 wire _06113_;
 wire net36;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire net35;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire net34;
 wire _06133_;
 wire _06134_;
 wire net33;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire net32;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire net3473;
 wire net3480;
 wire net3528;
 wire _06202_;
 wire net3527;
 wire net3478;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire net3475;
 wire _06210_;
 wire net3555;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire net3559;
 wire _06217_;
 wire clknet_leaf_63_clk_i_regs;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire net3558;
 wire net3471;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire clknet_leaf_62_clk_i_regs;
 wire _06236_;
 wire _06237_;
 wire net3645;
 wire net3526;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire net3537;
 wire _06259_;
 wire net3577;
 wire clknet_leaf_57_clk_i_regs;
 wire clknet_leaf_56_clk_i_regs;
 wire net3587;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire net3608;
 wire _06268_;
 wire clknet_leaf_1_clk_i_regs;
 wire clknet_leaf_54_clk_i_regs;
 wire _06271_;
 wire net3525;
 wire net3513;
 wire _06274_;
 wire _06275_;
 wire net3502;
 wire _06277_;
 wire net3470;
 wire net3505;
 wire net3491;
 wire net3512;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire net3524;
 wire clknet_leaf_53_clk_i_regs;
 wire net3536;
 wire net3664;
 wire _06289_;
 wire _06290_;
 wire net3619;
 wire net3663;
 wire net3508;
 wire net3507;
 wire net3511;
 wire net3492;
 wire _06297_;
 wire _06298_;
 wire net3489;
 wire net3501;
 wire net3500;
 wire _06302_;
 wire _06303_;
 wire net3499;
 wire net3510;
 wire net3618;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire net3535;
 wire _06312_;
 wire _06313_;
 wire clknet_leaf_51_clk_i_regs;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire net3586;
 wire _06334_;
 wire net3465;
 wire net3479;
 wire _06337_;
 wire _06338_;
 wire net3557;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire net3477;
 wire net3469;
 wire net3644;
 wire clknet_leaf_67_clk_i_regs;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire clknet_leaf_65_clk_i_regs;
 wire net3523;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire net3495;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire net3522;
 wire _06381_;
 wire _06382_;
 wire clknet_leaf_0_clk_i_regs;
 wire _06384_;
 wire clknet_leaf_49_clk_i_regs;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire clknet_leaf_48_clk_i_regs;
 wire clknet_leaf_47_clk_i_regs;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire net3514;
 wire _06402_;
 wire clknet_leaf_8_clk_i_regs;
 wire _06404_;
 wire net3493;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire net3625;
 wire net3519;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire net3454;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire net3430;
 wire net3431;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire net3429;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire net3423;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire net3418;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire net3422;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire net3412;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire net3420;
 wire net3419;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire net3426;
 wire net3411;
 wire _06538_;
 wire _06539_;
 wire net3463;
 wire _06541_;
 wire _06542_;
 wire net3404;
 wire net3407;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire net3408;
 wire net3462;
 wire net3413;
 wire _06554_;
 wire _06555_;
 wire net3481;
 wire net3397;
 wire _06558_;
 wire _06559_;
 wire net3396;
 wire _06561_;
 wire _06562_;
 wire net3395;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire net3394;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire net3393;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire net3488;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire net3460;
 wire net3392;
 wire _06590_;
 wire _06591_;
 wire net3391;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire net3390;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire net3389;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire net3388;
 wire _06617_;
 wire net3387;
 wire net3386;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire net3406;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire net3384;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire net3383;
 wire net3382;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire net3381;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire net3380;
 wire _06722_;
 wire net3379;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire net3378;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire net3377;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire net3376;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire net3374;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire net3405;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire net3375;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire net3370;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire net3369;
 wire _06845_;
 wire net3368;
 wire net3367;
 wire net3366;
 wire _06849_;
 wire net3364;
 wire _06851_;
 wire net3363;
 wire _06853_;
 wire net3362;
 wire net3361;
 wire _06856_;
 wire _06857_;
 wire net3360;
 wire _06859_;
 wire _06860_;
 wire net3358;
 wire _06862_;
 wire _06863_;
 wire net3357;
 wire _06865_;
 wire net3353;
 wire net3354;
 wire net3352;
 wire net3351;
 wire _06870_;
 wire net3350;
 wire _06872_;
 wire net3349;
 wire net3348;
 wire _06875_;
 wire net3347;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire net3346;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire net3345;
 wire net3344;
 wire net3343;
 wire net3359;
 wire _06900_;
 wire _06901_;
 wire net3342;
 wire net3459;
 wire _06904_;
 wire _06905_;
 wire net3458;
 wire net3402;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire net3425;
 wire _06928_;
 wire _06929_;
 wire net3410;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire net3341;
 wire _06938_;
 wire net3409;
 wire net3356;
 wire net3355;
 wire _06942_;
 wire _06943_;
 wire net3400;
 wire net3398;
 wire _06946_;
 wire net3372;
 wire net3339;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire net3401;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire net3371;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire net3340;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire net3334;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire net3333;
 wire _07019_;
 wire _07020_;
 wire net3403;
 wire net3416;
 wire net3414;
 wire net3417;
 wire _07025_;
 wire net3336;
 wire _07027_;
 wire net3421;
 wire _07029_;
 wire net3329;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire net3330;
 wire net576;
 wire net3325;
 wire _07041_;
 wire _07042_;
 wire net3327;
 wire _07044_;
 wire _07045_;
 wire net3328;
 wire _07047_;
 wire _07048_;
 wire net3322;
 wire net3424;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire net3324;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire net3319;
 wire _07065_;
 wire _07066_;
 wire net3318;
 wire net3457;
 wire net3455;
 wire net3337;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire net3326;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire net3315;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire net3531;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire net3313;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire net3320;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire net3317;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire net3312;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire net3428;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire net3323;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire net3314;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire net3316;
 wire _07311_;
 wire net3427;
 wire net3309;
 wire net3310;
 wire net3321;
 wire net3311;
 wire net3303;
 wire net3307;
 wire net3306;
 wire _07320_;
 wire net3298;
 wire net3293;
 wire net3292;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire net3297;
 wire net3294;
 wire net3291;
 wire net3296;
 wire _07331_;
 wire _07332_;
 wire net3304;
 wire net3302;
 wire _07335_;
 wire net3290;
 wire net3289;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire net3287;
 wire net3301;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire net3456;
 wire _07355_;
 wire _07356_;
 wire net560;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire net3300;
 wire net3286;
 wire _07375_;
 wire _07376_;
 wire net3530;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire net3295;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire net3433;
 wire net3494;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire net3461;
 wire net3285;
 wire _07432_;
 wire _07433_;
 wire net3468;
 wire net3283;
 wire net3280;
 wire _07437_;
 wire _07438_;
 wire net3277;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire net3279;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire net3276;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire net3272;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire net3271;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire net3275;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire net3504;
 wire _07717_;
 wire _07718_;
 wire net3268;
 wire net3267;
 wire _07721_;
 wire net3509;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire net3266;
 wire _07734_;
 wire net3503;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire net3273;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire net3263;
 wire net3467;
 wire _07764_;
 wire _07765_;
 wire net3466;
 wire net3579;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire net3534;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire net3617;
 wire net3265;
 wire _07823_;
 wire net3274;
 wire net3258;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire net3578;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire net3474;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire net3472;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire net3264;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire net3270;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire net3533;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire net3261;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire net3482;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire net3483;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire net3484;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire net3616;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire net3255;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire net3254;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire net3445;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire net3498;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire net3669;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire net3615;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire clknet_leaf_44_clk_i_regs;
 wire net3253;
 wire _08414_;
 wire net3257;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire net3252;
 wire net3256;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire net3250;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire net3497;
 wire net3247;
 wire net3248;
 wire _08476_;
 wire net3244;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire net3259;
 wire _08483_;
 wire _08484_;
 wire net3240;
 wire _08486_;
 wire net3241;
 wire _08488_;
 wire net3655;
 wire net3243;
 wire _08491_;
 wire net3238;
 wire _08493_;
 wire net3614;
 wire net3236;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire net3496;
 wire _08500_;
 wire _08501_;
 wire net3234;
 wire _08503_;
 wire net3251;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire net3227;
 wire net3648;
 wire _08520_;
 wire net3532;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire net3230;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire net3232;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire net3225;
 wire _08535_;
 wire net3228;
 wire clknet_leaf_4_clk_i_regs;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire net3221;
 wire net3613;
 wire _08543_;
 wire _08544_;
 wire net3231;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire net3233;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire net3224;
 wire net3220;
 wire _08556_;
 wire net3226;
 wire _08558_;
 wire net3219;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire net3216;
 wire net3222;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire net3214;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire net3218;
 wire _08573_;
 wire net3223;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire net3210;
 wire net3208;
 wire _08581_;
 wire _08583_;
 wire net3212;
 wire _08585_;
 wire _08586_;
 wire net3207;
 wire clknet_leaf_43_clk_i_regs;
 wire _08589_;
 wire net3203;
 wire net3453;
 wire _08592_;
 wire net3202;
 wire clknet_leaf_101_clk_i_regs;
 wire _08595_;
 wire clknet_leaf_100_clk_i_regs;
 wire clknet_leaf_98_clk_i_regs;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire net3201;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire net3476;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08615_;
 wire _08616_;
 wire clknet_leaf_97_clk_i_regs;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire net3662;
 wire _08624_;
 wire clknet_leaf_95_clk_i_regs;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire net3199;
 wire net3091;
 wire net3194;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire net3195;
 wire net3191;
 wire net3092;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire net3643;
 wire net3100;
 wire net858;
 wire net3120;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire net3518;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire net3517;
 wire net3136;
 wire _08733_;
 wire _08734_;
 wire net3190;
 wire _08736_;
 wire net3137;
 wire _08738_;
 wire _08739_;
 wire net3134;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire net3452;
 wire net3145;
 wire net3146;
 wire net3151;
 wire net3161;
 wire net3162;
 wire net3165;
 wire net3166;
 wire _08756_;
 wire net3167;
 wire _08758_;
 wire _08759_;
 wire net3170;
 wire net3169;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire net3168;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire net3171;
 wire _08788_;
 wire _08789_;
 wire net3188;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire net3172;
 wire net3173;
 wire _08798_;
 wire _08799_;
 wire net3175;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire net3176;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire net3177;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire net3183;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire net3192;
 wire net3447;
 wire _08836_;
 wire _08837_;
 wire net3178;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire net3451;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire net3450;
 wire net3180;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire net3449;
 wire _08880_;
 wire _08881_;
 wire net3181;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire net3446;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire net3182;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire net3205;
 wire _08901_;
 wire net3184;
 wire net3200;
 wire net3189;
 wire _08905_;
 wire _08906_;
 wire net3197;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire net3186;
 wire _08912_;
 wire net3187;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire net3193;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire net3196;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire net3198;
 wire _08934_;
 wire _08935_;
 wire net3209;
 wire _08937_;
 wire _08938_;
 wire net3206;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire net3213;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire net3237;
 wire _08953_;
 wire net3239;
 wire _08955_;
 wire _08956_;
 wire net3448;
 wire net3249;
 wire _08959_;
 wire net3262;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire net3281;
 wire _08965_;
 wire _08966_;
 wire net3432;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire net3278;
 wire _08975_;
 wire net3288;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire net3299;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire net3284;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire net3305;
 wire _08992_;
 wire net3332;
 wire net3335;
 wire _08995_;
 wire net3338;
 wire _08997_;
 wire net3385;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire net3373;
 wire net3399;
 wire clknet_leaf_7_clk_i_regs;
 wire clknet_leaf_42_clk_i_regs;
 wire clknet_leaf_40_clk_i_regs;
 wire net3590;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire net3589;
 wire net3576;
 wire _09016_;
 wire net3588;
 wire _09018_;
 wire net3596;
 wire _09020_;
 wire net3580;
 wire _09022_;
 wire _09023_;
 wire net3595;
 wire net3594;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire net3593;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire net3592;
 wire net3591;
 wire _09046_;
 wire net3624;
 wire net3623;
 wire net3605;
 wire net3602;
 wire net3604;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire net3601;
 wire _09060_;
 wire net3599;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire net3164;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire net3163;
 wire clknet_0_clk_i;
 wire net3174;
 wire _09079_;
 wire _09080_;
 wire net3158;
 wire _09082_;
 wire _09083_;
 wire net255;
 wire net3539;
 wire _09086_;
 wire clknet_leaf_104_clk_i_regs;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire clknet_leaf_108_clk_i_regs;
 wire clknet_leaf_106_clk_i_regs;
 wire _09104_;
 wire _09105_;
 wire clknet_leaf_109_clk_i_regs;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire clknet_leaf_110_clk_i_regs;
 wire _09121_;
 wire _09122_;
 wire clknet_leaf_111_clk_i_regs;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire clknet_leaf_112_clk_i_regs;
 wire clknet_leaf_113_clk_i_regs;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire clknet_leaf_119_clk_i_regs;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire clknet_leaf_122_clk_i_regs;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire clknet_leaf_124_clk_i_regs;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire clknet_leaf_125_clk_i_regs;
 wire net3159;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire clknet_leaf_126_clk_i_regs;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire net3156;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire net3204;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire net3154;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire net3185;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire net3153;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire net3152;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire net3211;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire net3150;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire net3365;
 wire net3520;
 wire net3521;
 wire net3464;
 wire net3415;
 wire net3179;
 wire net31;
 wire clk_i_regs;
 wire \alu_adder_result_ex[0] ;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire \alu_adder_result_ex[1] ;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net30;
 wire net2;
 wire net1;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire clk;
 wire core_busy_d;
 wire core_busy_q;
 wire \core_clock_gate_i.en_latch ;
 wire net150;
 wire \cs_registers_i.csr_depc_o[10] ;
 wire \cs_registers_i.csr_depc_o[11] ;
 wire \cs_registers_i.csr_depc_o[12] ;
 wire \cs_registers_i.csr_depc_o[13] ;
 wire \cs_registers_i.csr_depc_o[14] ;
 wire \cs_registers_i.csr_depc_o[15] ;
 wire \cs_registers_i.csr_depc_o[16] ;
 wire \cs_registers_i.csr_depc_o[17] ;
 wire \cs_registers_i.csr_depc_o[18] ;
 wire \cs_registers_i.csr_depc_o[19] ;
 wire \cs_registers_i.csr_depc_o[1] ;
 wire \cs_registers_i.csr_depc_o[20] ;
 wire \cs_registers_i.csr_depc_o[21] ;
 wire \cs_registers_i.csr_depc_o[22] ;
 wire \cs_registers_i.csr_depc_o[23] ;
 wire \cs_registers_i.csr_depc_o[24] ;
 wire \cs_registers_i.csr_depc_o[25] ;
 wire \cs_registers_i.csr_depc_o[26] ;
 wire \cs_registers_i.csr_depc_o[27] ;
 wire \cs_registers_i.csr_depc_o[28] ;
 wire \cs_registers_i.csr_depc_o[29] ;
 wire \cs_registers_i.csr_depc_o[2] ;
 wire \cs_registers_i.csr_depc_o[30] ;
 wire \cs_registers_i.csr_depc_o[31] ;
 wire \cs_registers_i.csr_depc_o[3] ;
 wire \cs_registers_i.csr_depc_o[4] ;
 wire \cs_registers_i.csr_depc_o[5] ;
 wire \cs_registers_i.csr_depc_o[6] ;
 wire \cs_registers_i.csr_depc_o[7] ;
 wire \cs_registers_i.csr_depc_o[8] ;
 wire \cs_registers_i.csr_depc_o[9] ;
 wire \cs_registers_i.csr_mepc_o[0] ;
 wire \cs_registers_i.csr_mepc_o[10] ;
 wire \cs_registers_i.csr_mepc_o[11] ;
 wire \cs_registers_i.csr_mepc_o[12] ;
 wire \cs_registers_i.csr_mepc_o[13] ;
 wire \cs_registers_i.csr_mepc_o[14] ;
 wire \cs_registers_i.csr_mepc_o[15] ;
 wire \cs_registers_i.csr_mepc_o[16] ;
 wire \cs_registers_i.csr_mepc_o[17] ;
 wire \cs_registers_i.csr_mepc_o[18] ;
 wire \cs_registers_i.csr_mepc_o[19] ;
 wire \cs_registers_i.csr_mepc_o[1] ;
 wire \cs_registers_i.csr_mepc_o[20] ;
 wire \cs_registers_i.csr_mepc_o[21] ;
 wire \cs_registers_i.csr_mepc_o[22] ;
 wire \cs_registers_i.csr_mepc_o[23] ;
 wire \cs_registers_i.csr_mepc_o[24] ;
 wire \cs_registers_i.csr_mepc_o[25] ;
 wire \cs_registers_i.csr_mepc_o[26] ;
 wire \cs_registers_i.csr_mepc_o[27] ;
 wire \cs_registers_i.csr_mepc_o[28] ;
 wire \cs_registers_i.csr_mepc_o[29] ;
 wire \cs_registers_i.csr_mepc_o[2] ;
 wire \cs_registers_i.csr_mepc_o[30] ;
 wire \cs_registers_i.csr_mepc_o[31] ;
 wire \cs_registers_i.csr_mepc_o[3] ;
 wire \cs_registers_i.csr_mepc_o[4] ;
 wire \cs_registers_i.csr_mepc_o[5] ;
 wire \cs_registers_i.csr_mepc_o[6] ;
 wire \cs_registers_i.csr_mepc_o[7] ;
 wire \cs_registers_i.csr_mepc_o[8] ;
 wire \cs_registers_i.csr_mepc_o[9] ;
 wire \cs_registers_i.csr_mstatus_mie_o ;
 wire \cs_registers_i.csr_mstatus_tw_o ;
 wire \cs_registers_i.csr_mtvec_o[10] ;
 wire \cs_registers_i.csr_mtvec_o[11] ;
 wire \cs_registers_i.csr_mtvec_o[12] ;
 wire \cs_registers_i.csr_mtvec_o[13] ;
 wire \cs_registers_i.csr_mtvec_o[14] ;
 wire \cs_registers_i.csr_mtvec_o[15] ;
 wire \cs_registers_i.csr_mtvec_o[16] ;
 wire \cs_registers_i.csr_mtvec_o[17] ;
 wire \cs_registers_i.csr_mtvec_o[18] ;
 wire \cs_registers_i.csr_mtvec_o[19] ;
 wire \cs_registers_i.csr_mtvec_o[20] ;
 wire \cs_registers_i.csr_mtvec_o[21] ;
 wire \cs_registers_i.csr_mtvec_o[22] ;
 wire \cs_registers_i.csr_mtvec_o[23] ;
 wire \cs_registers_i.csr_mtvec_o[24] ;
 wire \cs_registers_i.csr_mtvec_o[25] ;
 wire \cs_registers_i.csr_mtvec_o[26] ;
 wire \cs_registers_i.csr_mtvec_o[27] ;
 wire \cs_registers_i.csr_mtvec_o[28] ;
 wire \cs_registers_i.csr_mtvec_o[29] ;
 wire \cs_registers_i.csr_mtvec_o[30] ;
 wire \cs_registers_i.csr_mtvec_o[31] ;
 wire \cs_registers_i.csr_mtvec_o[8] ;
 wire \cs_registers_i.csr_mtvec_o[9] ;
 wire \cs_registers_i.dcsr_q[0] ;
 wire \cs_registers_i.dcsr_q[11] ;
 wire \cs_registers_i.dcsr_q[12] ;
 wire \cs_registers_i.dcsr_q[13] ;
 wire \cs_registers_i.dcsr_q[15] ;
 wire \cs_registers_i.dcsr_q[1] ;
 wire \cs_registers_i.dcsr_q[2] ;
 wire \cs_registers_i.dcsr_q[6] ;
 wire \cs_registers_i.dcsr_q[7] ;
 wire \cs_registers_i.dcsr_q[8] ;
 wire \cs_registers_i.debug_mode_i ;
 wire \cs_registers_i.dscratch0_q[0] ;
 wire \cs_registers_i.dscratch0_q[10] ;
 wire \cs_registers_i.dscratch0_q[11] ;
 wire \cs_registers_i.dscratch0_q[12] ;
 wire \cs_registers_i.dscratch0_q[13] ;
 wire \cs_registers_i.dscratch0_q[14] ;
 wire \cs_registers_i.dscratch0_q[15] ;
 wire \cs_registers_i.dscratch0_q[16] ;
 wire \cs_registers_i.dscratch0_q[17] ;
 wire \cs_registers_i.dscratch0_q[18] ;
 wire \cs_registers_i.dscratch0_q[19] ;
 wire \cs_registers_i.dscratch0_q[1] ;
 wire \cs_registers_i.dscratch0_q[20] ;
 wire \cs_registers_i.dscratch0_q[21] ;
 wire \cs_registers_i.dscratch0_q[22] ;
 wire \cs_registers_i.dscratch0_q[23] ;
 wire \cs_registers_i.dscratch0_q[24] ;
 wire \cs_registers_i.dscratch0_q[25] ;
 wire \cs_registers_i.dscratch0_q[26] ;
 wire \cs_registers_i.dscratch0_q[27] ;
 wire \cs_registers_i.dscratch0_q[28] ;
 wire \cs_registers_i.dscratch0_q[29] ;
 wire \cs_registers_i.dscratch0_q[2] ;
 wire \cs_registers_i.dscratch0_q[30] ;
 wire \cs_registers_i.dscratch0_q[31] ;
 wire \cs_registers_i.dscratch0_q[3] ;
 wire \cs_registers_i.dscratch0_q[4] ;
 wire \cs_registers_i.dscratch0_q[5] ;
 wire \cs_registers_i.dscratch0_q[6] ;
 wire \cs_registers_i.dscratch0_q[7] ;
 wire \cs_registers_i.dscratch0_q[8] ;
 wire \cs_registers_i.dscratch0_q[9] ;
 wire \cs_registers_i.dscratch1_q[0] ;
 wire \cs_registers_i.dscratch1_q[10] ;
 wire \cs_registers_i.dscratch1_q[11] ;
 wire \cs_registers_i.dscratch1_q[12] ;
 wire \cs_registers_i.dscratch1_q[13] ;
 wire \cs_registers_i.dscratch1_q[14] ;
 wire \cs_registers_i.dscratch1_q[15] ;
 wire \cs_registers_i.dscratch1_q[16] ;
 wire \cs_registers_i.dscratch1_q[17] ;
 wire \cs_registers_i.dscratch1_q[18] ;
 wire \cs_registers_i.dscratch1_q[19] ;
 wire \cs_registers_i.dscratch1_q[1] ;
 wire \cs_registers_i.dscratch1_q[20] ;
 wire \cs_registers_i.dscratch1_q[21] ;
 wire \cs_registers_i.dscratch1_q[22] ;
 wire \cs_registers_i.dscratch1_q[23] ;
 wire \cs_registers_i.dscratch1_q[24] ;
 wire \cs_registers_i.dscratch1_q[25] ;
 wire \cs_registers_i.dscratch1_q[26] ;
 wire \cs_registers_i.dscratch1_q[27] ;
 wire \cs_registers_i.dscratch1_q[28] ;
 wire \cs_registers_i.dscratch1_q[29] ;
 wire \cs_registers_i.dscratch1_q[2] ;
 wire \cs_registers_i.dscratch1_q[30] ;
 wire \cs_registers_i.dscratch1_q[31] ;
 wire \cs_registers_i.dscratch1_q[3] ;
 wire \cs_registers_i.dscratch1_q[4] ;
 wire \cs_registers_i.dscratch1_q[5] ;
 wire \cs_registers_i.dscratch1_q[6] ;
 wire \cs_registers_i.dscratch1_q[7] ;
 wire \cs_registers_i.dscratch1_q[8] ;
 wire \cs_registers_i.dscratch1_q[9] ;
 wire \cs_registers_i.mcause_q[0] ;
 wire \cs_registers_i.mcause_q[1] ;
 wire \cs_registers_i.mcause_q[2] ;
 wire \cs_registers_i.mcause_q[3] ;
 wire \cs_registers_i.mcause_q[4] ;
 wire \cs_registers_i.mcause_q[5] ;
 wire \cs_registers_i.mcountinhibit_q[0] ;
 wire \cs_registers_i.mcountinhibit_q[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[10] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[11] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[12] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[13] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[14] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[15] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[16] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[17] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[18] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[19] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[1] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[20] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[21] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[22] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[23] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[24] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[25] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[26] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[27] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[28] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[29] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[30] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[31] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[32] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[33] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[34] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[35] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[36] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[37] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[38] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[39] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[3] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[40] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[41] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[42] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[43] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[44] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[45] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[46] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[47] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[48] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[49] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[4] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[50] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[51] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[52] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[53] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[54] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[55] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[56] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[57] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[58] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[59] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[5] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[60] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[61] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[62] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[63] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[6] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[7] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[8] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[9] ;
 wire \cs_registers_i.mhpmcounter[1856] ;
 wire \cs_registers_i.mhpmcounter[1857] ;
 wire \cs_registers_i.mhpmcounter[1858] ;
 wire \cs_registers_i.mhpmcounter[1859] ;
 wire \cs_registers_i.mhpmcounter[1860] ;
 wire \cs_registers_i.mhpmcounter[1861] ;
 wire \cs_registers_i.mhpmcounter[1862] ;
 wire \cs_registers_i.mhpmcounter[1863] ;
 wire \cs_registers_i.mhpmcounter[1864] ;
 wire \cs_registers_i.mhpmcounter[1865] ;
 wire \cs_registers_i.mhpmcounter[1866] ;
 wire \cs_registers_i.mhpmcounter[1867] ;
 wire \cs_registers_i.mhpmcounter[1868] ;
 wire \cs_registers_i.mhpmcounter[1869] ;
 wire \cs_registers_i.mhpmcounter[1870] ;
 wire \cs_registers_i.mhpmcounter[1871] ;
 wire \cs_registers_i.mhpmcounter[1872] ;
 wire \cs_registers_i.mhpmcounter[1873] ;
 wire \cs_registers_i.mhpmcounter[1874] ;
 wire \cs_registers_i.mhpmcounter[1875] ;
 wire \cs_registers_i.mhpmcounter[1876] ;
 wire \cs_registers_i.mhpmcounter[1877] ;
 wire \cs_registers_i.mhpmcounter[1878] ;
 wire \cs_registers_i.mhpmcounter[1879] ;
 wire \cs_registers_i.mhpmcounter[1880] ;
 wire \cs_registers_i.mhpmcounter[1881] ;
 wire \cs_registers_i.mhpmcounter[1882] ;
 wire \cs_registers_i.mhpmcounter[1883] ;
 wire \cs_registers_i.mhpmcounter[1884] ;
 wire \cs_registers_i.mhpmcounter[1885] ;
 wire \cs_registers_i.mhpmcounter[1886] ;
 wire \cs_registers_i.mhpmcounter[1887] ;
 wire \cs_registers_i.mhpmcounter[1888] ;
 wire \cs_registers_i.mhpmcounter[1889] ;
 wire \cs_registers_i.mhpmcounter[1890] ;
 wire \cs_registers_i.mhpmcounter[1891] ;
 wire \cs_registers_i.mhpmcounter[1892] ;
 wire \cs_registers_i.mhpmcounter[1893] ;
 wire \cs_registers_i.mhpmcounter[1894] ;
 wire \cs_registers_i.mhpmcounter[1895] ;
 wire \cs_registers_i.mhpmcounter[1896] ;
 wire \cs_registers_i.mhpmcounter[1897] ;
 wire \cs_registers_i.mhpmcounter[1898] ;
 wire \cs_registers_i.mhpmcounter[1899] ;
 wire \cs_registers_i.mhpmcounter[1900] ;
 wire \cs_registers_i.mhpmcounter[1901] ;
 wire \cs_registers_i.mhpmcounter[1902] ;
 wire \cs_registers_i.mhpmcounter[1903] ;
 wire \cs_registers_i.mhpmcounter[1904] ;
 wire \cs_registers_i.mhpmcounter[1905] ;
 wire \cs_registers_i.mhpmcounter[1906] ;
 wire \cs_registers_i.mhpmcounter[1907] ;
 wire \cs_registers_i.mhpmcounter[1908] ;
 wire \cs_registers_i.mhpmcounter[1909] ;
 wire \cs_registers_i.mhpmcounter[1910] ;
 wire \cs_registers_i.mhpmcounter[1911] ;
 wire \cs_registers_i.mhpmcounter[1912] ;
 wire \cs_registers_i.mhpmcounter[1913] ;
 wire \cs_registers_i.mhpmcounter[1914] ;
 wire \cs_registers_i.mhpmcounter[1915] ;
 wire \cs_registers_i.mhpmcounter[1916] ;
 wire \cs_registers_i.mhpmcounter[1917] ;
 wire \cs_registers_i.mhpmcounter[1918] ;
 wire \cs_registers_i.mhpmcounter[1919] ;
 wire \cs_registers_i.mie_q[0] ;
 wire \cs_registers_i.mie_q[10] ;
 wire \cs_registers_i.mie_q[11] ;
 wire \cs_registers_i.mie_q[12] ;
 wire \cs_registers_i.mie_q[13] ;
 wire \cs_registers_i.mie_q[14] ;
 wire \cs_registers_i.mie_q[15] ;
 wire \cs_registers_i.mie_q[16] ;
 wire \cs_registers_i.mie_q[17] ;
 wire \cs_registers_i.mie_q[1] ;
 wire \cs_registers_i.mie_q[2] ;
 wire \cs_registers_i.mie_q[3] ;
 wire \cs_registers_i.mie_q[4] ;
 wire \cs_registers_i.mie_q[5] ;
 wire \cs_registers_i.mie_q[6] ;
 wire \cs_registers_i.mie_q[7] ;
 wire \cs_registers_i.mie_q[8] ;
 wire \cs_registers_i.mie_q[9] ;
 wire \cs_registers_i.mscratch_q[0] ;
 wire \cs_registers_i.mscratch_q[10] ;
 wire \cs_registers_i.mscratch_q[11] ;
 wire \cs_registers_i.mscratch_q[12] ;
 wire \cs_registers_i.mscratch_q[13] ;
 wire \cs_registers_i.mscratch_q[14] ;
 wire \cs_registers_i.mscratch_q[15] ;
 wire \cs_registers_i.mscratch_q[16] ;
 wire \cs_registers_i.mscratch_q[17] ;
 wire \cs_registers_i.mscratch_q[18] ;
 wire \cs_registers_i.mscratch_q[19] ;
 wire \cs_registers_i.mscratch_q[1] ;
 wire \cs_registers_i.mscratch_q[20] ;
 wire \cs_registers_i.mscratch_q[21] ;
 wire \cs_registers_i.mscratch_q[22] ;
 wire \cs_registers_i.mscratch_q[23] ;
 wire \cs_registers_i.mscratch_q[24] ;
 wire \cs_registers_i.mscratch_q[25] ;
 wire \cs_registers_i.mscratch_q[26] ;
 wire \cs_registers_i.mscratch_q[27] ;
 wire \cs_registers_i.mscratch_q[28] ;
 wire \cs_registers_i.mscratch_q[29] ;
 wire \cs_registers_i.mscratch_q[2] ;
 wire \cs_registers_i.mscratch_q[30] ;
 wire \cs_registers_i.mscratch_q[31] ;
 wire \cs_registers_i.mscratch_q[3] ;
 wire \cs_registers_i.mscratch_q[4] ;
 wire \cs_registers_i.mscratch_q[5] ;
 wire \cs_registers_i.mscratch_q[6] ;
 wire \cs_registers_i.mscratch_q[7] ;
 wire \cs_registers_i.mscratch_q[8] ;
 wire \cs_registers_i.mscratch_q[9] ;
 wire \cs_registers_i.mstack_cause_q[0] ;
 wire \cs_registers_i.mstack_cause_q[1] ;
 wire \cs_registers_i.mstack_cause_q[2] ;
 wire \cs_registers_i.mstack_cause_q[3] ;
 wire \cs_registers_i.mstack_cause_q[4] ;
 wire \cs_registers_i.mstack_cause_q[5] ;
 wire \cs_registers_i.mstack_epc_q[0] ;
 wire \cs_registers_i.mstack_epc_q[10] ;
 wire \cs_registers_i.mstack_epc_q[11] ;
 wire \cs_registers_i.mstack_epc_q[12] ;
 wire \cs_registers_i.mstack_epc_q[13] ;
 wire \cs_registers_i.mstack_epc_q[14] ;
 wire \cs_registers_i.mstack_epc_q[15] ;
 wire \cs_registers_i.mstack_epc_q[16] ;
 wire \cs_registers_i.mstack_epc_q[17] ;
 wire \cs_registers_i.mstack_epc_q[18] ;
 wire \cs_registers_i.mstack_epc_q[19] ;
 wire \cs_registers_i.mstack_epc_q[1] ;
 wire \cs_registers_i.mstack_epc_q[20] ;
 wire \cs_registers_i.mstack_epc_q[21] ;
 wire \cs_registers_i.mstack_epc_q[22] ;
 wire \cs_registers_i.mstack_epc_q[23] ;
 wire \cs_registers_i.mstack_epc_q[24] ;
 wire \cs_registers_i.mstack_epc_q[25] ;
 wire \cs_registers_i.mstack_epc_q[26] ;
 wire \cs_registers_i.mstack_epc_q[27] ;
 wire \cs_registers_i.mstack_epc_q[28] ;
 wire \cs_registers_i.mstack_epc_q[29] ;
 wire \cs_registers_i.mstack_epc_q[2] ;
 wire \cs_registers_i.mstack_epc_q[30] ;
 wire \cs_registers_i.mstack_epc_q[31] ;
 wire \cs_registers_i.mstack_epc_q[3] ;
 wire \cs_registers_i.mstack_epc_q[4] ;
 wire \cs_registers_i.mstack_epc_q[5] ;
 wire \cs_registers_i.mstack_epc_q[6] ;
 wire \cs_registers_i.mstack_epc_q[7] ;
 wire \cs_registers_i.mstack_epc_q[8] ;
 wire \cs_registers_i.mstack_epc_q[9] ;
 wire \cs_registers_i.mstack_q[0] ;
 wire \cs_registers_i.mstack_q[1] ;
 wire \cs_registers_i.mstack_q[2] ;
 wire \cs_registers_i.mstatus_q[1] ;
 wire \cs_registers_i.mstatus_q[2] ;
 wire \cs_registers_i.mstatus_q[3] ;
 wire \cs_registers_i.mstatus_q[4] ;
 wire \cs_registers_i.mtval_q[0] ;
 wire \cs_registers_i.mtval_q[10] ;
 wire \cs_registers_i.mtval_q[11] ;
 wire \cs_registers_i.mtval_q[12] ;
 wire \cs_registers_i.mtval_q[13] ;
 wire \cs_registers_i.mtval_q[14] ;
 wire \cs_registers_i.mtval_q[15] ;
 wire \cs_registers_i.mtval_q[16] ;
 wire \cs_registers_i.mtval_q[17] ;
 wire \cs_registers_i.mtval_q[18] ;
 wire \cs_registers_i.mtval_q[19] ;
 wire \cs_registers_i.mtval_q[1] ;
 wire \cs_registers_i.mtval_q[20] ;
 wire \cs_registers_i.mtval_q[21] ;
 wire \cs_registers_i.mtval_q[22] ;
 wire \cs_registers_i.mtval_q[23] ;
 wire \cs_registers_i.mtval_q[24] ;
 wire \cs_registers_i.mtval_q[25] ;
 wire \cs_registers_i.mtval_q[26] ;
 wire \cs_registers_i.mtval_q[27] ;
 wire \cs_registers_i.mtval_q[28] ;
 wire \cs_registers_i.mtval_q[29] ;
 wire \cs_registers_i.mtval_q[2] ;
 wire \cs_registers_i.mtval_q[30] ;
 wire \cs_registers_i.mtval_q[31] ;
 wire \cs_registers_i.mtval_q[3] ;
 wire \cs_registers_i.mtval_q[4] ;
 wire \cs_registers_i.mtval_q[5] ;
 wire \cs_registers_i.mtval_q[6] ;
 wire \cs_registers_i.mtval_q[7] ;
 wire \cs_registers_i.mtval_q[8] ;
 wire \cs_registers_i.mtval_q[9] ;
 wire \cs_registers_i.nmi_mode_i ;
 wire \cs_registers_i.pc_id_i[10] ;
 wire \cs_registers_i.pc_id_i[11] ;
 wire \cs_registers_i.pc_id_i[12] ;
 wire \cs_registers_i.pc_id_i[13] ;
 wire \cs_registers_i.pc_id_i[14] ;
 wire \cs_registers_i.pc_id_i[15] ;
 wire \cs_registers_i.pc_id_i[16] ;
 wire \cs_registers_i.pc_id_i[17] ;
 wire \cs_registers_i.pc_id_i[18] ;
 wire \cs_registers_i.pc_id_i[19] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[20] ;
 wire \cs_registers_i.pc_id_i[21] ;
 wire \cs_registers_i.pc_id_i[22] ;
 wire \cs_registers_i.pc_id_i[23] ;
 wire \cs_registers_i.pc_id_i[24] ;
 wire \cs_registers_i.pc_id_i[25] ;
 wire \cs_registers_i.pc_id_i[26] ;
 wire \cs_registers_i.pc_id_i[27] ;
 wire \cs_registers_i.pc_id_i[28] ;
 wire \cs_registers_i.pc_id_i[29] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_id_i[30] ;
 wire \cs_registers_i.pc_id_i[31] ;
 wire \cs_registers_i.pc_id_i[3] ;
 wire \cs_registers_i.pc_id_i[4] ;
 wire \cs_registers_i.pc_id_i[5] ;
 wire \cs_registers_i.pc_id_i[6] ;
 wire \cs_registers_i.pc_id_i[7] ;
 wire \cs_registers_i.pc_id_i[8] ;
 wire \cs_registers_i.pc_id_i[9] ;
 wire \cs_registers_i.pc_if_i[10] ;
 wire \cs_registers_i.pc_if_i[11] ;
 wire \cs_registers_i.pc_if_i[12] ;
 wire \cs_registers_i.pc_if_i[13] ;
 wire \cs_registers_i.pc_if_i[14] ;
 wire \cs_registers_i.pc_if_i[15] ;
 wire \cs_registers_i.pc_if_i[16] ;
 wire \cs_registers_i.pc_if_i[17] ;
 wire \cs_registers_i.pc_if_i[18] ;
 wire \cs_registers_i.pc_if_i[19] ;
 wire \cs_registers_i.pc_if_i[1] ;
 wire \cs_registers_i.pc_if_i[20] ;
 wire \cs_registers_i.pc_if_i[21] ;
 wire \cs_registers_i.pc_if_i[22] ;
 wire \cs_registers_i.pc_if_i[23] ;
 wire \cs_registers_i.pc_if_i[24] ;
 wire \cs_registers_i.pc_if_i[25] ;
 wire \cs_registers_i.pc_if_i[26] ;
 wire \cs_registers_i.pc_if_i[27] ;
 wire \cs_registers_i.pc_if_i[28] ;
 wire \cs_registers_i.pc_if_i[29] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.pc_if_i[30] ;
 wire \cs_registers_i.pc_if_i[31] ;
 wire \cs_registers_i.pc_if_i[3] ;
 wire \cs_registers_i.pc_if_i[4] ;
 wire \cs_registers_i.pc_if_i[5] ;
 wire \cs_registers_i.pc_if_i[6] ;
 wire \cs_registers_i.pc_if_i[7] ;
 wire \cs_registers_i.pc_if_i[8] ;
 wire \cs_registers_i.pc_if_i[9] ;
 wire \cs_registers_i.priv_mode_id_o[0] ;
 wire \cs_registers_i.priv_mode_id_o[1] ;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire \ex_block_i.alu_i.imd_val_q_i[0] ;
 wire \ex_block_i.alu_i.imd_val_q_i[10] ;
 wire \ex_block_i.alu_i.imd_val_q_i[11] ;
 wire \ex_block_i.alu_i.imd_val_q_i[12] ;
 wire \ex_block_i.alu_i.imd_val_q_i[13] ;
 wire \ex_block_i.alu_i.imd_val_q_i[14] ;
 wire \ex_block_i.alu_i.imd_val_q_i[15] ;
 wire \ex_block_i.alu_i.imd_val_q_i[16] ;
 wire \ex_block_i.alu_i.imd_val_q_i[17] ;
 wire \ex_block_i.alu_i.imd_val_q_i[18] ;
 wire \ex_block_i.alu_i.imd_val_q_i[19] ;
 wire \ex_block_i.alu_i.imd_val_q_i[1] ;
 wire \ex_block_i.alu_i.imd_val_q_i[20] ;
 wire \ex_block_i.alu_i.imd_val_q_i[21] ;
 wire \ex_block_i.alu_i.imd_val_q_i[22] ;
 wire \ex_block_i.alu_i.imd_val_q_i[23] ;
 wire \ex_block_i.alu_i.imd_val_q_i[24] ;
 wire \ex_block_i.alu_i.imd_val_q_i[25] ;
 wire \ex_block_i.alu_i.imd_val_q_i[26] ;
 wire \ex_block_i.alu_i.imd_val_q_i[27] ;
 wire \ex_block_i.alu_i.imd_val_q_i[28] ;
 wire \ex_block_i.alu_i.imd_val_q_i[29] ;
 wire \ex_block_i.alu_i.imd_val_q_i[2] ;
 wire \ex_block_i.alu_i.imd_val_q_i[30] ;
 wire \ex_block_i.alu_i.imd_val_q_i[31] ;
 wire \ex_block_i.alu_i.imd_val_q_i[32] ;
 wire \ex_block_i.alu_i.imd_val_q_i[33] ;
 wire \ex_block_i.alu_i.imd_val_q_i[34] ;
 wire \ex_block_i.alu_i.imd_val_q_i[35] ;
 wire \ex_block_i.alu_i.imd_val_q_i[36] ;
 wire \ex_block_i.alu_i.imd_val_q_i[37] ;
 wire \ex_block_i.alu_i.imd_val_q_i[38] ;
 wire \ex_block_i.alu_i.imd_val_q_i[39] ;
 wire \ex_block_i.alu_i.imd_val_q_i[3] ;
 wire \ex_block_i.alu_i.imd_val_q_i[40] ;
 wire \ex_block_i.alu_i.imd_val_q_i[41] ;
 wire \ex_block_i.alu_i.imd_val_q_i[42] ;
 wire \ex_block_i.alu_i.imd_val_q_i[43] ;
 wire \ex_block_i.alu_i.imd_val_q_i[44] ;
 wire \ex_block_i.alu_i.imd_val_q_i[45] ;
 wire \ex_block_i.alu_i.imd_val_q_i[46] ;
 wire \ex_block_i.alu_i.imd_val_q_i[47] ;
 wire \ex_block_i.alu_i.imd_val_q_i[48] ;
 wire \ex_block_i.alu_i.imd_val_q_i[49] ;
 wire \ex_block_i.alu_i.imd_val_q_i[4] ;
 wire \ex_block_i.alu_i.imd_val_q_i[50] ;
 wire \ex_block_i.alu_i.imd_val_q_i[51] ;
 wire \ex_block_i.alu_i.imd_val_q_i[52] ;
 wire \ex_block_i.alu_i.imd_val_q_i[53] ;
 wire \ex_block_i.alu_i.imd_val_q_i[54] ;
 wire \ex_block_i.alu_i.imd_val_q_i[55] ;
 wire \ex_block_i.alu_i.imd_val_q_i[56] ;
 wire \ex_block_i.alu_i.imd_val_q_i[57] ;
 wire \ex_block_i.alu_i.imd_val_q_i[58] ;
 wire \ex_block_i.alu_i.imd_val_q_i[59] ;
 wire \ex_block_i.alu_i.imd_val_q_i[5] ;
 wire \ex_block_i.alu_i.imd_val_q_i[60] ;
 wire \ex_block_i.alu_i.imd_val_q_i[61] ;
 wire \ex_block_i.alu_i.imd_val_q_i[62] ;
 wire \ex_block_i.alu_i.imd_val_q_i[63] ;
 wire \ex_block_i.alu_i.imd_val_q_i[6] ;
 wire \ex_block_i.alu_i.imd_val_q_i[7] ;
 wire \ex_block_i.alu_i.imd_val_q_i[8] ;
 wire \ex_block_i.alu_i.imd_val_q_i[9] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ;
 wire fetch_enable_q;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[4] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[4] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1000] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1001] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1002] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1003] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1004] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1005] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1006] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1007] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1008] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1009] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[100] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1010] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1011] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1012] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1013] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1014] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1015] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1016] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1017] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1018] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1019] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[101] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1020] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1021] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1022] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1023] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[102] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[103] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[104] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[105] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[106] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[107] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[108] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[109] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[110] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[111] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[112] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[113] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[114] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[115] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[116] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[117] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[118] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[119] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[120] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[121] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[122] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[123] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[124] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[125] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[126] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[127] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[128] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[129] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[130] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[131] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[132] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[133] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[134] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[135] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[136] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[137] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[138] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[139] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[140] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[141] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[142] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[143] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[144] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[145] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[146] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[147] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[148] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[149] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[150] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[151] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[152] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[153] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[154] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[155] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[156] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[157] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[158] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[159] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[160] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[161] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[162] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[163] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[164] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[165] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[166] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[167] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[168] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[169] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[170] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[171] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[172] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[173] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[174] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[175] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[176] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[177] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[178] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[179] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[180] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[181] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[182] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[183] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[184] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[185] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[186] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[187] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[188] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[189] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[190] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[191] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[192] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[193] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[194] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[195] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[196] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[197] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[198] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[199] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[200] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[201] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[202] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[203] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[204] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[205] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[206] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[207] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[208] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[209] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[210] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[211] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[212] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[213] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[214] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[215] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[216] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[217] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[218] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[219] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[220] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[221] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[222] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[223] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[224] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[225] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[226] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[227] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[228] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[229] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[230] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[231] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[232] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[233] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[234] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[235] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[236] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[237] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[238] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[239] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[240] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[241] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[242] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[243] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[244] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[245] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[246] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[247] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[248] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[249] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[250] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[251] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[252] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[253] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[254] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[255] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[256] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[257] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[258] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[259] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[260] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[261] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[262] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[263] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[264] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[265] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[266] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[267] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[268] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[269] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[270] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[271] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[272] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[273] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[274] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[275] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[276] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[277] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[278] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[279] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[280] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[281] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[282] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[283] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[284] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[285] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[286] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[287] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[288] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[289] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[290] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[291] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[292] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[293] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[294] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[295] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[296] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[297] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[298] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[299] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[300] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[301] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[302] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[303] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[304] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[305] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[306] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[307] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[308] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[309] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[310] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[311] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[312] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[313] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[314] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[315] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[316] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[317] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[318] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[319] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[320] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[321] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[322] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[323] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[324] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[325] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[326] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[327] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[328] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[329] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[32] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[330] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[331] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[332] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[333] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[334] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[335] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[336] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[337] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[338] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[339] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[33] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[340] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[341] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[342] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[343] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[344] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[345] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[346] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[347] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[348] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[349] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[34] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[350] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[351] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[352] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[353] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[354] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[355] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[356] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[357] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[358] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[359] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[35] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[360] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[361] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[362] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[363] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[364] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[365] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[366] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[367] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[368] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[369] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[36] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[370] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[371] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[372] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[373] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[374] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[375] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[376] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[377] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[378] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[379] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[37] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[380] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[381] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[382] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[383] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[384] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[385] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[386] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[387] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[388] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[389] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[38] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[390] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[391] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[392] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[393] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[394] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[395] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[396] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[397] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[398] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[399] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[39] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[400] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[401] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[402] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[403] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[404] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[405] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[406] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[407] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[408] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[409] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[40] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[410] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[411] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[412] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[413] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[414] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[415] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[416] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[417] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[418] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[419] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[41] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[420] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[421] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[422] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[423] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[424] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[425] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[426] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[427] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[428] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[429] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[42] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[430] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[431] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[432] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[433] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[434] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[435] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[436] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[437] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[438] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[439] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[43] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[440] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[441] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[442] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[443] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[444] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[445] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[446] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[447] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[448] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[449] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[44] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[450] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[451] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[452] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[453] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[454] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[455] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[456] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[457] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[458] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[459] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[45] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[460] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[461] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[462] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[463] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[464] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[465] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[466] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[467] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[468] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[469] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[46] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[470] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[471] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[472] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[473] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[474] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[475] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[476] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[477] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[478] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[479] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[47] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[480] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[481] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[482] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[483] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[484] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[485] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[486] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[487] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[488] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[489] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[48] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[490] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[491] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[492] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[493] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[494] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[495] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[496] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[497] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[498] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[499] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[49] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[500] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[501] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[502] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[503] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[504] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[505] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[506] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[507] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[508] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[509] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[50] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[510] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[511] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[512] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[513] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[514] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[515] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[516] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[517] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[518] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[519] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[51] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[520] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[521] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[522] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[523] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[524] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[525] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[526] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[527] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[528] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[529] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[52] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[530] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[531] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[532] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[533] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[534] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[535] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[536] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[537] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[538] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[539] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[53] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[540] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[541] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[542] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[543] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[544] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[545] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[546] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[547] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[548] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[549] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[54] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[550] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[551] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[552] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[553] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[554] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[555] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[556] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[557] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[558] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[559] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[55] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[560] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[561] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[562] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[563] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[564] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[565] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[566] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[567] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[568] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[569] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[56] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[570] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[571] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[572] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[573] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[574] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[575] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[576] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[577] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[578] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[579] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[57] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[580] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[581] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[582] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[583] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[584] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[585] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[586] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[587] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[588] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[589] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[58] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[590] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[591] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[592] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[593] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[594] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[595] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[596] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[597] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[598] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[599] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[59] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[600] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[601] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[602] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[603] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[604] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[605] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[606] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[607] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[608] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[609] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[60] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[610] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[611] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[612] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[613] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[614] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[615] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[616] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[617] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[618] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[619] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[61] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[620] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[621] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[622] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[623] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[624] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[625] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[626] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[627] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[628] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[629] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[62] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[630] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[631] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[632] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[633] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[634] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[635] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[636] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[637] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[638] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[639] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[63] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[640] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[641] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[642] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[643] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[644] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[645] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[646] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[647] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[648] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[649] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[64] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[650] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[651] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[652] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[653] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[654] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[655] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[656] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[657] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[658] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[659] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[65] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[660] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[661] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[662] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[663] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[664] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[665] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[666] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[667] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[668] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[669] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[66] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[670] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[671] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[672] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[673] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[674] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[675] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[676] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[677] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[678] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[679] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[67] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[680] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[681] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[682] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[683] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[684] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[685] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[686] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[687] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[688] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[689] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[68] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[690] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[691] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[692] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[693] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[694] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[695] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[696] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[697] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[698] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[699] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[69] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[700] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[701] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[702] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[703] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[704] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[705] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[706] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[707] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[708] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[709] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[70] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[710] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[711] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[712] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[713] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[714] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[715] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[716] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[717] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[718] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[719] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[71] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[720] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[721] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[722] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[723] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[724] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[725] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[726] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[727] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[728] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[729] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[72] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[730] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[731] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[732] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[733] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[734] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[735] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[736] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[737] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[738] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[739] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[73] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[740] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[741] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[742] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[743] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[744] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[745] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[746] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[747] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[748] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[749] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[74] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[750] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[751] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[752] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[753] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[754] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[755] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[756] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[757] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[758] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[759] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[75] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[760] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[761] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[762] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[763] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[764] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[765] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[766] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[767] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[768] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[769] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[76] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[770] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[771] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[772] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[773] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[774] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[775] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[776] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[777] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[778] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[779] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[77] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[780] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[781] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[782] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[783] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[784] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[785] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[786] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[787] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[788] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[789] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[78] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[790] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[791] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[792] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[793] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[794] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[795] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[796] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[797] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[798] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[799] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[79] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[800] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[801] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[802] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[803] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[804] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[805] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[806] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[807] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[808] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[809] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[80] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[810] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[811] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[812] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[813] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[814] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[815] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[816] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[817] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[818] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[819] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[81] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[820] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[821] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[822] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[823] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[824] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[825] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[826] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[827] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[828] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[829] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[82] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[830] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[831] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[832] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[833] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[834] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[835] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[836] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[837] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[838] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[839] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[83] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[840] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[841] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[842] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[843] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[844] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[845] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[846] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[847] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[848] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[849] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[84] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[850] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[851] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[852] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[853] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[854] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[855] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[856] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[857] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[858] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[859] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[85] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[860] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[861] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[862] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[863] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[864] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[865] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[866] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[867] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[868] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[869] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[86] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[870] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[871] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[872] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[873] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[874] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[875] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[876] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[877] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[878] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[879] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[87] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[880] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[881] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[882] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[883] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[884] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[885] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[886] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[887] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[888] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[889] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[88] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[890] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[891] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[892] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[893] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[894] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[895] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[896] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[897] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[898] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[899] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[89] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[900] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[901] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[902] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[903] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[904] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[905] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[906] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[907] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[908] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[909] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[90] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[910] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[911] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[912] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[913] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[914] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[915] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[916] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[917] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[918] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[919] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[91] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[920] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[921] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[922] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[923] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[924] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[925] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[926] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[927] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[928] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[929] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[92] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[930] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[931] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[932] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[933] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[934] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[935] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[936] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[937] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[938] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[939] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[93] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[940] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[941] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[942] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[943] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[944] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[945] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[946] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[947] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[948] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[949] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[94] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[950] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[951] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[952] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[953] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[954] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[955] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[956] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[957] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[958] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[959] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[95] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[960] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[961] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[962] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[963] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[964] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[965] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[966] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[967] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[968] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[969] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[96] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[970] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[971] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[972] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[973] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[974] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[975] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[976] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[977] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[978] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[979] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[97] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[980] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[981] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[982] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[983] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[984] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[985] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[986] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[987] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[988] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[989] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[98] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[990] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[991] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[992] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[993] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[994] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[995] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[996] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[997] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[998] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[999] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[99] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[4] ;
 wire \id_stage_i.branch_set ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[0] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[1] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[2] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[3] ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.exc_req_q ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.illegal_insn_q ;
 wire \id_stage_i.controller_i.instr_compressed_i[0] ;
 wire \id_stage_i.controller_i.instr_compressed_i[10] ;
 wire \id_stage_i.controller_i.instr_compressed_i[11] ;
 wire \id_stage_i.controller_i.instr_compressed_i[12] ;
 wire \id_stage_i.controller_i.instr_compressed_i[13] ;
 wire \id_stage_i.controller_i.instr_compressed_i[14] ;
 wire \id_stage_i.controller_i.instr_compressed_i[15] ;
 wire \id_stage_i.controller_i.instr_compressed_i[1] ;
 wire \id_stage_i.controller_i.instr_compressed_i[2] ;
 wire \id_stage_i.controller_i.instr_compressed_i[3] ;
 wire \id_stage_i.controller_i.instr_compressed_i[4] ;
 wire \id_stage_i.controller_i.instr_compressed_i[5] ;
 wire \id_stage_i.controller_i.instr_compressed_i[6] ;
 wire \id_stage_i.controller_i.instr_compressed_i[7] ;
 wire \id_stage_i.controller_i.instr_compressed_i[8] ;
 wire \id_stage_i.controller_i.instr_compressed_i[9] ;
 wire \id_stage_i.controller_i.instr_fetch_err_i ;
 wire \id_stage_i.controller_i.instr_fetch_err_plus2_i ;
 wire \id_stage_i.controller_i.instr_i[0] ;
 wire \id_stage_i.controller_i.instr_i[12] ;
 wire \id_stage_i.controller_i.instr_i[13] ;
 wire \id_stage_i.controller_i.instr_i[14] ;
 wire \id_stage_i.controller_i.instr_i[1] ;
 wire \id_stage_i.controller_i.instr_i[25] ;
 wire \id_stage_i.controller_i.instr_i[26] ;
 wire \id_stage_i.controller_i.instr_i[27] ;
 wire \id_stage_i.controller_i.instr_i[28] ;
 wire \id_stage_i.controller_i.instr_i[29] ;
 wire \id_stage_i.controller_i.instr_i[2] ;
 wire \id_stage_i.controller_i.instr_i[30] ;
 wire \id_stage_i.controller_i.instr_i[31] ;
 wire \id_stage_i.controller_i.instr_i[3] ;
 wire \id_stage_i.controller_i.instr_i[4] ;
 wire \id_stage_i.controller_i.instr_i[5] ;
 wire \id_stage_i.controller_i.instr_i[6] ;
 wire \id_stage_i.controller_i.instr_is_compressed_i ;
 wire \id_stage_i.controller_i.instr_valid_i ;
 wire \id_stage_i.controller_i.load_err_i ;
 wire \id_stage_i.controller_i.load_err_q ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[0] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[10] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[11] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[12] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[13] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[14] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[15] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[16] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[17] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[18] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[19] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[1] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[20] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[21] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[22] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[23] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[24] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[25] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[26] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[27] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[28] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[29] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[2] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[30] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[31] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[3] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[4] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[5] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[6] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[7] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[8] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[9] ;
 wire \id_stage_i.controller_i.store_err_i ;
 wire \id_stage_i.controller_i.store_err_q ;
 wire \id_stage_i.decoder_i.illegal_c_insn_i ;
 wire \id_stage_i.id_fsm_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire \load_store_unit_i.data_sign_ext_q ;
 wire \load_store_unit_i.data_type_q[1] ;
 wire \load_store_unit_i.data_type_q[2] ;
 wire \load_store_unit_i.data_we_q ;
 wire \load_store_unit_i.handle_misaligned_q ;
 wire \load_store_unit_i.ls_fsm_cs[0] ;
 wire \load_store_unit_i.ls_fsm_cs[1] ;
 wire \load_store_unit_i.ls_fsm_cs[2] ;
 wire \load_store_unit_i.lsu_err_q ;
 wire \load_store_unit_i.rdata_offset_q[0] ;
 wire \load_store_unit_i.rdata_offset_q[1] ;
 wire \load_store_unit_i.rdata_q[0] ;
 wire \load_store_unit_i.rdata_q[10] ;
 wire \load_store_unit_i.rdata_q[11] ;
 wire \load_store_unit_i.rdata_q[12] ;
 wire \load_store_unit_i.rdata_q[13] ;
 wire \load_store_unit_i.rdata_q[14] ;
 wire \load_store_unit_i.rdata_q[15] ;
 wire \load_store_unit_i.rdata_q[16] ;
 wire \load_store_unit_i.rdata_q[17] ;
 wire \load_store_unit_i.rdata_q[18] ;
 wire \load_store_unit_i.rdata_q[19] ;
 wire \load_store_unit_i.rdata_q[1] ;
 wire \load_store_unit_i.rdata_q[20] ;
 wire \load_store_unit_i.rdata_q[21] ;
 wire \load_store_unit_i.rdata_q[22] ;
 wire \load_store_unit_i.rdata_q[23] ;
 wire \load_store_unit_i.rdata_q[2] ;
 wire \load_store_unit_i.rdata_q[3] ;
 wire \load_store_unit_i.rdata_q[4] ;
 wire \load_store_unit_i.rdata_q[5] ;
 wire \load_store_unit_i.rdata_q[6] ;
 wire \load_store_unit_i.rdata_q[7] ;
 wire \load_store_unit_i.rdata_q[8] ;
 wire \load_store_unit_i.rdata_q[9] ;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3490;
 wire net3506;
 wire net3529;
 wire net3560;
 wire net3556;
 wire net3600;
 wire net3603;
 wire net3598;
 wire net3597;
 wire net3607;
 wire net251;
 wire net3611;
 wire net3606;
 wire net3610;
 wire net3441;
 wire net3649;
 wire net3440;
 wire net3571;
 wire clknet_leaf_89_clk_i_regs;
 wire clknet_leaf_87_clk_i_regs;
 wire clknet_leaf_84_clk_i_regs;
 wire clknet_leaf_80_clk_i_regs;
 wire clknet_leaf_79_clk_i_regs;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_60_clk_i_regs;
 wire net3568;
 wire net3609;
 wire net3583;
 wire net3635;
 wire net3585;
 wire net3582;
 wire net3242;
 wire net3581;
 wire net3439;
 wire clknet_leaf_36_clk_i_regs;
 wire net3229;
 wire net3438;
 wire clknet_leaf_35_clk_i_regs;
 wire net254;
 wire net3437;
 wire clknet_leaf_34_clk_i_regs;
 wire clknet_leaf_12_clk_i_regs;
 wire net3124;
 wire net3122;
 wire net3436;
 wire net3133;
 wire clknet_leaf_31_clk_i_regs;
 wire clknet_leaf_29_clk_i_regs;
 wire net3132;
 wire net3435;
 wire clknet_leaf_11_clk_i_regs;
 wire net3217;
 wire net3538;
 wire clknet_leaf_26_clk_i_regs;
 wire net3434;
 wire net3622;
 wire net3130;
 wire net3140;
 wire clknet_leaf_28_clk_i_regs;
 wire net3620;
 wire clknet_leaf_24_clk_i_regs;
 wire clknet_leaf_18_clk_i_regs;
 wire net3621;
 wire clknet_leaf_17_clk_i_regs;
 wire clknet_leaf_23_clk_i_regs;
 wire clknet_leaf_22_clk_i_regs;
 wire clknet_leaf_27_clk_i_regs;
 wire net3135;
 wire net3282;
 wire net3144;
 wire net3269;
 wire net3260;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_leaf_10_clk_i_regs;
 wire clknet_leaf_20_clk_i_regs;
 wire net3246;
 wire net3245;
 wire clknet_leaf_77_clk_i_regs;
 wire clknet_leaf_75_clk_i_regs;
 wire clknet_leaf_74_clk_i_regs;
 wire net3634;
 wire net3633;
 wire clknet_leaf_71_clk_i_regs;
 wire clknet_leaf_68_clk_i_regs;
 wire net3632;
 wire net3552;
 wire net3551;
 wire net3550;
 wire clknet_leaf_102_clk_i_regs;
 wire net3547;
 wire clknet_leaf_58_clk_i_regs;
 wire net3546;
 wire net3540;
 wire net3647;
 wire net3646;
 wire net3549;
 wire net3569;
 wire net3545;
 wire net3544;
 wire net3543;
 wire net3548;
 wire net3541;
 wire net3542;
 wire net3659;
 wire net3567;
 wire net3631;
 wire net3087;
 wire net3630;
 wire net3650;
 wire net3629;
 wire net3657;
 wire net3628;
 wire net3570;
 wire net3627;
 wire net253;
 wire net3083;
 wire net3099;
 wire net3075;
 wire net3073;
 wire net3626;
 wire net3072;
 wire net3112;
 wire net3575;
 wire net3574;
 wire net3069;
 wire net3111;
 wire net3061;
 wire net3667;
 wire net250;
 wire net3064;
 wire net3078;
 wire net3068;
 wire net3110;
 wire net3063;
 wire net3666;
 wire net3070;
 wire net3051;
 wire net3059;
 wire net3050;
 wire net3677;
 wire net3675;
 wire net3674;
 wire net3654;
 wire net3661;
 wire net3656;
 wire net3658;
 wire net3660;
 wire net3573;
 wire net3572;
 wire net3673;
 wire net3668;
 wire net3672;
 wire net3671;
 wire net3676;
 wire clknet_leaf_468_clk_i_regs;
 wire clknet_leaf_469_clk_i_regs;
 wire clknet_leaf_470_clk_i_regs;
 wire clknet_leaf_473_clk_i_regs;
 wire clknet_leaf_476_clk_i_regs;
 wire clknet_leaf_478_clk_i_regs;
 wire clknet_leaf_480_clk_i_regs;
 wire clknet_leaf_483_clk_i_regs;
 wire clknet_leaf_484_clk_i_regs;
 wire clknet_leaf_486_clk_i_regs;
 wire clknet_leaf_488_clk_i_regs;
 wire clknet_leaf_492_clk_i_regs;
 wire clknet_leaf_493_clk_i_regs;
 wire clknet_leaf_494_clk_i_regs;
 wire clknet_leaf_495_clk_i_regs;
 wire clknet_leaf_497_clk_i_regs;
 wire clknet_leaf_498_clk_i_regs;
 wire clknet_leaf_501_clk_i_regs;
 wire clknet_leaf_503_clk_i_regs;
 wire clknet_leaf_507_clk_i_regs;
 wire clknet_leaf_510_clk_i_regs;
 wire clknet_leaf_512_clk_i_regs;
 wire clknet_leaf_513_clk_i_regs;
 wire clknet_leaf_514_clk_i_regs;
 wire clknet_leaf_516_clk_i_regs;
 wire clknet_leaf_517_clk_i_regs;
 wire clknet_leaf_518_clk_i_regs;
 wire clknet_leaf_522_clk_i_regs;
 wire clknet_leaf_523_clk_i_regs;
 wire clknet_leaf_525_clk_i_regs;
 wire clknet_leaf_526_clk_i_regs;
 wire clknet_leaf_528_clk_i_regs;
 wire clknet_leaf_531_clk_i_regs;
 wire clknet_leaf_532_clk_i_regs;
 wire clknet_leaf_533_clk_i_regs;
 wire clknet_leaf_535_clk_i_regs;
 wire clknet_leaf_536_clk_i_regs;
 wire clknet_leaf_537_clk_i_regs;
 wire clknet_leaf_540_clk_i_regs;
 wire clknet_leaf_543_clk_i_regs;
 wire clknet_leaf_544_clk_i_regs;
 wire clknet_leaf_546_clk_i_regs;
 wire clknet_leaf_547_clk_i_regs;
 wire clknet_leaf_548_clk_i_regs;
 wire clknet_leaf_549_clk_i_regs;
 wire clknet_leaf_550_clk_i_regs;
 wire clknet_leaf_551_clk_i_regs;
 wire clknet_leaf_556_clk_i_regs;
 wire clknet_leaf_557_clk_i_regs;
 wire clknet_leaf_558_clk_i_regs;
 wire clknet_leaf_559_clk_i_regs;
 wire clknet_leaf_560_clk_i_regs;
 wire clknet_leaf_561_clk_i_regs;
 wire clknet_leaf_563_clk_i_regs;
 wire clknet_leaf_565_clk_i_regs;
 wire clknet_leaf_566_clk_i_regs;
 wire clknet_leaf_571_clk_i_regs;
 wire clknet_0_clk_i_regs;
 wire clknet_3_0_0_clk_i_regs;
 wire clknet_3_1_0_clk_i_regs;
 wire clknet_3_2_0_clk_i_regs;
 wire clknet_3_3_0_clk_i_regs;
 wire clknet_3_4_0_clk_i_regs;
 wire clknet_3_5_0_clk_i_regs;
 wire clknet_3_6_0_clk_i_regs;
 wire clknet_3_7_0_clk_i_regs;
 wire clknet_6_0__leaf_clk_i_regs;
 wire clknet_6_1__leaf_clk_i_regs;
 wire clknet_6_2__leaf_clk_i_regs;
 wire clknet_6_3__leaf_clk_i_regs;
 wire clknet_6_4__leaf_clk_i_regs;
 wire clknet_6_5__leaf_clk_i_regs;
 wire clknet_6_6__leaf_clk_i_regs;
 wire clknet_6_7__leaf_clk_i_regs;
 wire clknet_6_8__leaf_clk_i_regs;
 wire clknet_6_9__leaf_clk_i_regs;
 wire clknet_6_10__leaf_clk_i_regs;
 wire clknet_6_11__leaf_clk_i_regs;
 wire clknet_6_12__leaf_clk_i_regs;
 wire clknet_6_13__leaf_clk_i_regs;
 wire clknet_6_14__leaf_clk_i_regs;
 wire clknet_6_15__leaf_clk_i_regs;
 wire clknet_6_16__leaf_clk_i_regs;
 wire clknet_6_17__leaf_clk_i_regs;
 wire clknet_6_18__leaf_clk_i_regs;
 wire clknet_6_19__leaf_clk_i_regs;
 wire clknet_6_20__leaf_clk_i_regs;
 wire clknet_6_21__leaf_clk_i_regs;
 wire clknet_6_22__leaf_clk_i_regs;
 wire clknet_6_23__leaf_clk_i_regs;
 wire clknet_6_24__leaf_clk_i_regs;
 wire clknet_6_25__leaf_clk_i_regs;
 wire clknet_6_26__leaf_clk_i_regs;
 wire clknet_6_27__leaf_clk_i_regs;
 wire clknet_6_28__leaf_clk_i_regs;
 wire clknet_6_29__leaf_clk_i_regs;
 wire clknet_6_30__leaf_clk_i_regs;
 wire clknet_6_31__leaf_clk_i_regs;
 wire clknet_6_32__leaf_clk_i_regs;
 wire clknet_6_33__leaf_clk_i_regs;
 wire clknet_6_34__leaf_clk_i_regs;
 wire clknet_6_35__leaf_clk_i_regs;
 wire clknet_6_36__leaf_clk_i_regs;
 wire clknet_6_37__leaf_clk_i_regs;
 wire clknet_6_38__leaf_clk_i_regs;
 wire clknet_6_39__leaf_clk_i_regs;
 wire clknet_6_40__leaf_clk_i_regs;
 wire clknet_6_41__leaf_clk_i_regs;
 wire clknet_6_42__leaf_clk_i_regs;
 wire clknet_6_43__leaf_clk_i_regs;
 wire clknet_6_44__leaf_clk_i_regs;
 wire clknet_6_45__leaf_clk_i_regs;
 wire clknet_6_46__leaf_clk_i_regs;
 wire clknet_6_47__leaf_clk_i_regs;
 wire clknet_6_48__leaf_clk_i_regs;
 wire clknet_6_49__leaf_clk_i_regs;
 wire clknet_6_50__leaf_clk_i_regs;
 wire clknet_6_51__leaf_clk_i_regs;
 wire clknet_6_52__leaf_clk_i_regs;
 wire clknet_6_53__leaf_clk_i_regs;
 wire clknet_6_54__leaf_clk_i_regs;
 wire clknet_6_55__leaf_clk_i_regs;
 wire clknet_6_56__leaf_clk_i_regs;
 wire clknet_6_57__leaf_clk_i_regs;
 wire clknet_6_58__leaf_clk_i_regs;
 wire clknet_6_59__leaf_clk_i_regs;
 wire clknet_6_60__leaf_clk_i_regs;
 wire clknet_6_61__leaf_clk_i_regs;
 wire clknet_6_62__leaf_clk_i_regs;
 wire clknet_6_63__leaf_clk_i_regs;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_328_clk;
 wire clknet_leaf_331_clk;
 wire clknet_leaf_332_clk;
 wire clknet_leaf_335_clk;
 wire clknet_leaf_336_clk;
 wire clknet_leaf_344_clk;
 wire clknet_leaf_345_clk;
 wire clknet_leaf_351_clk;
 wire clknet_leaf_352_clk;
 wire clknet_leaf_353_clk;
 wire clknet_leaf_354_clk;
 wire clknet_leaf_358_clk;
 wire clknet_leaf_360_clk;
 wire clknet_leaf_361_clk;
 wire clknet_leaf_363_clk;
 wire clknet_leaf_364_clk;
 wire clknet_leaf_365_clk;
 wire clknet_leaf_366_clk;
 wire clknet_leaf_372_clk;
 wire clknet_leaf_375_clk;
 wire clknet_leaf_376_clk;
 wire clknet_leaf_377_clk;
 wire clknet_leaf_378_clk;
 wire clknet_leaf_382_clk;
 wire clknet_leaf_383_clk;
 wire clknet_leaf_384_clk;
 wire clknet_leaf_385_clk;
 wire clknet_leaf_390_clk;
 wire clknet_leaf_398_clk;
 wire clknet_leaf_401_clk;
 wire clknet_leaf_403_clk;
 wire clknet_leaf_406_clk;
 wire clknet_leaf_407_clk;
 wire clknet_leaf_408_clk;
 wire clknet_leaf_409_clk;
 wire clknet_leaf_410_clk;
 wire clknet_leaf_413_clk;
 wire clknet_leaf_420_clk;
 wire clknet_leaf_423_clk;
 wire clknet_leaf_425_clk;
 wire clknet_leaf_426_clk;
 wire clknet_leaf_427_clk;
 wire clknet_leaf_428_clk;
 wire clknet_leaf_436_clk;
 wire clknet_leaf_437_clk;
 wire clknet_leaf_440_clk;
 wire clknet_leaf_452_clk;
 wire clknet_leaf_455_clk;
 wire clknet_leaf_459_clk;
 wire clknet_leaf_468_clk;
 wire clknet_leaf_475_clk;
 wire clknet_leaf_476_clk;
 wire clknet_leaf_479_clk;
 wire clknet_leaf_485_clk;
 wire clknet_leaf_486_clk;
 wire clknet_leaf_489_clk;
 wire clknet_leaf_494_clk;
 wire clknet_leaf_495_clk;
 wire clknet_leaf_497_clk;
 wire clknet_leaf_498_clk;
 wire clknet_leaf_499_clk;
 wire clknet_leaf_501_clk;
 wire clknet_leaf_502_clk;
 wire clknet_leaf_503_clk;
 wire clknet_leaf_504_clk;
 wire clknet_leaf_511_clk;
 wire clknet_leaf_514_clk;
 wire clknet_leaf_515_clk;
 wire clknet_leaf_520_clk;
 wire clknet_leaf_521_clk;
 wire clknet_leaf_522_clk;
 wire clknet_leaf_528_clk;
 wire clknet_leaf_530_clk;
 wire clknet_leaf_531_clk;
 wire clknet_leaf_532_clk;
 wire clknet_leaf_533_clk;
 wire clknet_leaf_534_clk;
 wire clknet_leaf_537_clk;
 wire clknet_leaf_539_clk;
 wire clknet_leaf_540_clk;
 wire clknet_leaf_543_clk;
 wire clknet_leaf_544_clk;
 wire clknet_leaf_546_clk;
 wire clknet_leaf_549_clk;
 wire clknet_leaf_550_clk;
 wire clknet_leaf_552_clk;
 wire clknet_leaf_553_clk;
 wire clknet_leaf_555_clk;
 wire clknet_leaf_559_clk;
 wire clknet_leaf_560_clk;
 wire clknet_leaf_564_clk;
 wire clknet_leaf_567_clk;
 wire clknet_leaf_569_clk;
 wire clknet_leaf_570_clk;
 wire clknet_leaf_571_clk;
 wire clknet_leaf_572_clk;
 wire clknet_leaf_573_clk;
 wire clknet_leaf_575_clk;
 wire clknet_leaf_580_clk;
 wire clknet_leaf_583_clk;
 wire clknet_leaf_584_clk;
 wire clknet_leaf_587_clk;
 wire clknet_leaf_588_clk;
 wire clknet_leaf_589_clk;
 wire clknet_leaf_590_clk;
 wire clknet_leaf_592_clk;
 wire clknet_leaf_593_clk;
 wire clknet_leaf_594_clk;
 wire clknet_leaf_601_clk;
 wire clknet_leaf_608_clk;
 wire clknet_leaf_609_clk;
 wire clknet_leaf_610_clk;
 wire clknet_leaf_611_clk;
 wire clknet_leaf_612_clk;
 wire clknet_leaf_620_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire delaynet_0_core_clock;
 wire delaynet_1_core_clock;
 wire delaynet_2_core_clock;
 wire delaynet_3_core_clock;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net484;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net386;
 wire net387;
 wire net391;
 wire net392;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net459;
 wire net460;
 wire net464;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net528;
 wire net529;
 wire net530;
 wire net547;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net575;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net737;
 wire net584;
 wire net585;
 wire net625;
 wire net627;
 wire net632;
 wire net633;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net335;
 wire net343;
 wire net344;
 wire net345;
 wire net385;
 wire net388;
 wire net389;
 wire net390;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net455;
 wire net458;
 wire net461;
 wire net462;
 wire net463;
 wire net465;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net485;
 wire net486;
 wire net487;
 wire net738;
 wire [0:0] _09744_;
 wire [0:0] _09745_;
 wire [0:0] _09746_;
 wire [0:0] _09747_;
 wire [0:0] _09748_;
 wire [0:0] _09749_;
 wire [0:0] _09750_;
 wire [0:0] _09751_;
 wire [0:0] _09752_;
 wire [0:0] _09753_;
 wire [0:0] _09754_;
 wire [0:0] _09755_;
 wire [0:0] _09756_;
 wire [0:0] _09757_;
 wire [0:0] _09758_;
 wire [0:0] _09759_;
 wire [0:0] _09760_;
 wire [0:0] _09761_;
 wire [0:0] _09762_;
 wire [0:0] _09763_;
 wire [0:0] _09764_;
 wire [0:0] _09765_;
 wire [0:0] _09766_;
 wire [0:0] _09767_;
 wire [0:0] _09768_;
 wire [0:0] _09769_;
 wire [0:0] _09770_;
 wire [0:0] _09771_;
 wire [0:0] _09772_;
 wire [0:0] _09773_;
 wire [0:0] _09774_;
 wire [0:0] _09775_;
 wire [0:0] _09776_;
 wire [0:0] _09777_;
 wire [0:0] _09778_;
 wire [0:0] _09779_;
 wire [0:0] _09780_;
 wire [0:0] _09781_;
 wire [0:0] _09782_;
 wire [0:0] _09783_;
 wire [0:0] _09784_;
 wire [0:0] _09785_;
 wire [0:0] _09786_;
 wire [0:0] _09787_;
 wire [0:0] _09788_;
 wire [0:0] _09789_;
 wire [0:0] _09790_;
 wire [0:0] _09791_;
 wire [0:0] _09792_;
 wire [0:0] _09793_;
 wire [0:0] _09794_;
 wire [0:0] _09795_;
 wire [0:0] _09796_;
 wire [0:0] _09797_;
 wire [0:0] _09798_;
 wire [0:0] _09799_;
 wire [0:0] _09800_;
 wire [0:0] _09801_;
 wire [0:0] _09802_;
 wire [0:0] _09803_;
 wire [0:0] _09804_;
 wire [0:0] _09805_;
 wire [0:0] _09806_;
 wire [0:0] _09807_;
 wire [0:0] _09808_;
 wire [0:0] _09809_;
 wire [0:0] _09810_;
 wire [0:0] _09811_;
 wire [0:0] _09812_;
 wire [0:0] _09813_;
 wire [0:0] _09814_;
 wire [0:0] _09815_;
 wire [0:0] _09816_;
 wire [0:0] _09817_;
 wire [0:0] _09818_;
 wire [0:0] _09819_;
 wire [0:0] _09820_;
 wire [0:0] _09821_;
 wire [0:0] _09822_;
 wire [0:0] _09823_;
 wire [0:0] _09824_;
 wire [0:0] _09825_;
 wire [0:0] _09826_;
 wire [0:0] _09827_;
 wire [0:0] _09828_;
 wire [0:0] _09829_;
 wire [0:0] _09830_;
 wire [0:0] _09831_;
 wire [0:0] _09832_;
 wire [0:0] _09833_;
 wire [0:0] _09834_;
 wire [0:0] _09835_;
 wire [0:0] _09836_;
 wire [0:0] _09837_;
 wire [0:0] _09838_;
 wire [0:0] _09839_;
 wire [0:0] _09840_;
 wire [0:0] _09841_;
 wire [0:0] _09842_;
 wire [0:0] _09843_;
 wire [0:0] _09844_;
 wire [0:0] _09845_;
 wire [0:0] _09846_;
 wire [0:0] _09847_;
 wire [0:0] _09848_;
 wire [0:0] _09849_;
 wire [0:0] _09850_;
 wire [0:0] _09851_;
 wire [0:0] _09852_;
 wire [0:0] _09853_;
 wire [0:0] _09854_;
 wire [0:0] _09855_;
 wire [0:0] _09856_;
 wire [0:0] _09857_;
 wire [0:0] _09858_;
 wire [0:0] _09859_;
 wire [0:0] _09860_;
 wire [0:0] _09861_;
 wire [0:0] _09862_;
 wire [0:0] _09863_;
 wire [0:0] _09864_;
 wire [0:0] _09865_;
 wire [0:0] _09866_;
 wire [0:0] _09867_;
 wire [0:0] _09868_;
 wire [0:0] _09869_;
 wire [0:0] _09870_;
 wire [0:0] _09871_;
 wire [0:0] _09872_;
 wire [0:0] _09873_;
 wire [0:0] _09874_;
 wire [0:0] _09875_;
 wire [0:0] _09876_;
 wire [0:0] _09877_;
 wire [0:0] _09878_;
 wire [0:0] _09879_;
 wire [0:0] _09880_;
 wire [0:0] _09881_;
 wire [0:0] _09882_;
 wire [0:0] _09883_;
 wire [0:0] _09884_;
 wire [0:0] _09885_;
 wire [0:0] _09886_;
 wire [0:0] _09887_;
 wire [0:0] _09888_;
 wire [0:0] _09889_;
 wire [0:0] _09890_;
 wire [0:0] _09891_;
 wire [0:0] _09892_;
 wire [0:0] _09893_;
 wire [0:0] _09894_;
 wire [0:0] _09895_;
 wire [0:0] _09896_;
 wire [0:0] _09897_;
 wire [0:0] _09898_;
 wire [0:0] _09899_;
 wire [0:0] _09900_;
 wire [0:0] _09901_;
 wire [0:0] _09902_;
 wire [0:0] _09903_;
 wire [0:0] _09904_;
 wire [0:0] _09905_;
 wire [0:0] _09906_;
 wire [0:0] _09907_;
 wire [0:0] _09908_;
 wire [0:0] _09909_;
 wire [0:0] _09910_;
 wire [0:0] _09911_;
 wire [0:0] _09912_;
 wire [0:0] _09913_;
 wire [0:0] _09914_;
 wire [0:0] _09915_;
 wire [0:0] _09916_;
 wire [0:0] _09917_;
 wire [0:0] _09918_;
 wire [0:0] _09919_;
 wire [0:0] _09920_;
 wire [0:0] _09921_;
 wire [0:0] _09922_;
 wire [0:0] _09923_;
 wire [0:0] _09924_;
 wire [0:0] _09925_;
 wire [0:0] _09926_;
 wire [0:0] _09927_;
 wire [0:0] _09928_;
 wire [0:0] _09929_;
 wire [0:0] _09930_;
 wire [0:0] _09931_;
 wire [0:0] _09932_;
 wire [0:0] _09933_;
 wire [0:0] _09934_;
 wire [0:0] _09935_;
 wire [0:0] _09936_;
 wire [0:0] _09937_;
 wire [0:0] _09938_;
 wire [0:0] _09939_;
 wire [0:0] _09940_;
 wire [0:0] _09941_;
 wire [0:0] _09942_;
 wire [0:0] _09943_;
 wire [0:0] _09944_;
 wire [0:0] _09945_;
 wire [0:0] _09946_;
 wire [0:0] _09947_;
 wire [0:0] _09948_;
 wire [0:0] _09949_;
 wire [0:0] _09950_;
 wire [0:0] _09951_;
 wire [0:0] _09952_;
 wire [0:0] _09953_;
 wire [0:0] _09954_;
 wire [0:0] _09955_;
 wire [0:0] _09956_;
 wire [0:0] _09957_;
 wire [0:0] _09958_;
 wire [0:0] _09959_;
 wire [0:0] _09960_;
 wire [0:0] _09961_;
 wire [0:0] _09962_;
 wire [0:0] _09963_;
 wire [0:0] _09964_;
 wire [0:0] _09965_;
 wire [0:0] _09966_;
 wire [0:0] _09967_;
 wire [0:0] _09968_;
 wire [0:0] _09969_;
 wire [0:0] _09970_;
 wire [0:0] _09971_;
 wire [0:0] _09972_;
 wire [0:0] _09973_;
 wire [0:0] _09974_;
 wire [0:0] _09975_;
 wire [0:0] _09976_;
 wire [0:0] _09977_;
 wire [0:0] _09978_;
 wire [0:0] _09979_;
 wire [0:0] _09980_;
 wire [0:0] _09981_;
 wire [0:0] _09982_;
 wire [0:0] _09983_;
 wire [0:0] _09984_;
 wire [0:0] _09985_;
 wire [0:0] _09986_;
 wire [0:0] _09987_;
 wire [0:0] _09988_;
 wire [0:0] _09989_;
 wire [0:0] _09990_;
 wire [0:0] _09991_;
 wire [0:0] _09992_;
 wire [0:0] _09993_;
 wire [0:0] _09994_;
 wire [0:0] _09995_;
 wire [0:0] _09996_;
 wire [0:0] _09997_;
 wire [0:0] _09998_;
 wire [0:0] _09999_;
 wire [0:0] _10000_;
 wire [0:0] _10001_;
 wire [0:0] _10002_;
 wire [0:0] _10003_;
 wire [0:0] _10004_;
 wire [0:0] _10005_;
 wire [0:0] _10006_;
 wire [0:0] _10007_;
 wire [0:0] _10008_;
 wire [0:0] _10009_;
 wire [0:0] _10010_;
 wire [0:0] _10011_;
 wire [0:0] _10012_;
 wire [0:0] _10013_;
 wire [0:0] _10014_;
 wire [0:0] _10015_;
 wire [0:0] _10016_;
 wire [0:0] _10017_;
 wire [0:0] _10018_;
 wire [0:0] _10019_;
 wire [0:0] _10020_;
 wire [0:0] _10021_;
 wire [0:0] _10022_;
 wire [0:0] _10023_;
 wire [0:0] _10024_;
 wire [0:0] _10025_;
 wire [0:0] _10026_;
 wire [0:0] _10027_;
 wire [0:0] _10028_;
 wire [0:0] _10029_;
 wire [0:0] _10030_;
 wire [0:0] _10031_;
 wire [0:0] _10032_;
 wire [0:0] _10033_;
 wire [0:0] _10034_;
 wire [0:0] _10035_;
 wire [0:0] _10036_;
 wire [0:0] _10037_;
 wire [0:0] _10038_;
 wire [0:0] _10039_;
 wire [0:0] _10040_;
 wire [0:0] _10041_;
 wire [0:0] _10042_;
 wire [0:0] _10043_;
 wire [0:0] _10044_;
 wire [0:0] _10045_;
 wire [0:0] _10046_;
 wire [0:0] _10047_;
 wire [0:0] _10048_;
 wire [0:0] _10049_;
 wire [0:0] _10050_;
 wire [0:0] _10051_;
 wire [0:0] _10052_;
 wire [0:0] _10053_;
 wire [0:0] _10054_;
 wire [0:0] _10055_;
 wire [0:0] _10056_;
 wire [0:0] _10057_;
 wire [0:0] _10058_;
 wire [0:0] _10059_;
 wire [0:0] _10060_;
 wire [0:0] _10061_;
 wire [0:0] _10062_;
 wire [0:0] _10063_;
 wire [0:0] _10064_;
 wire [0:0] _10065_;
 wire [0:0] _10066_;
 wire [0:0] _10067_;
 wire [0:0] _10068_;
 wire [0:0] _10069_;
 wire [0:0] _10070_;
 wire [0:0] _10071_;
 wire [0:0] _10072_;
 wire [0:0] _10073_;
 wire [0:0] _10074_;
 wire [0:0] _10075_;
 wire [0:0] _10076_;
 wire [0:0] _10077_;
 wire [0:0] _10078_;
 wire [0:0] _10079_;
 wire [0:0] _10080_;
 wire [0:0] _10081_;
 wire [0:0] _10082_;
 wire [0:0] _10083_;
 wire [0:0] _10084_;
 wire [0:0] _10085_;
 wire [0:0] _10086_;
 wire [0:0] _10087_;
 wire [0:0] _10088_;
 wire [0:0] _10089_;
 wire [0:0] _10090_;
 wire [0:0] _10091_;
 wire [0:0] _10092_;
 wire [0:0] _10093_;
 wire [0:0] _10094_;
 wire [0:0] _10095_;
 wire [0:0] _10096_;
 wire [0:0] _10097_;
 wire [0:0] _10098_;
 wire [0:0] _10099_;
 wire [0:0] _10100_;
 wire [0:0] _10101_;
 wire [0:0] _10102_;
 wire [0:0] _10103_;
 wire [0:0] _10104_;
 wire [0:0] _10105_;
 wire [0:0] _10106_;
 wire [0:0] _10107_;
 wire [0:0] _10108_;
 wire [0:0] _10109_;
 wire [0:0] _10110_;
 wire [0:0] _10111_;
 wire [0:0] _10112_;
 wire [0:0] _10113_;
 wire [0:0] _10114_;
 wire [0:0] _10115_;
 wire [0:0] _10116_;
 wire [0:0] _10117_;
 wire [0:0] _10118_;
 wire [0:0] _10119_;
 wire [0:0] _10120_;
 wire [0:0] _10121_;
 wire [0:0] _10122_;
 wire [0:0] _10123_;
 wire [0:0] _10124_;
 wire [0:0] _10125_;
 wire [0:0] _10126_;
 wire [0:0] _10127_;
 wire [0:0] _10128_;
 wire [0:0] _10129_;
 wire [0:0] _10130_;
 wire [0:0] _10131_;
 wire [0:0] _10132_;
 wire [0:0] _10133_;
 wire [0:0] _10134_;
 wire [0:0] _10135_;
 wire [0:0] _10136_;
 wire [0:0] _10137_;
 wire [0:0] _10138_;
 wire [0:0] _10139_;
 wire [0:0] _10140_;
 wire [0:0] _10141_;
 wire [0:0] _10142_;
 wire [0:0] _10143_;
 wire [0:0] _10144_;
 wire [0:0] _10145_;
 wire [0:0] _10146_;
 wire [0:0] _10147_;
 wire [0:0] _10148_;
 wire [0:0] _10149_;
 wire [0:0] _10150_;
 wire [0:0] _10151_;
 wire [0:0] _10152_;
 wire [0:0] _10153_;
 wire [0:0] _10154_;
 wire [0:0] _10155_;
 wire [0:0] _10156_;
 wire [0:0] _10157_;
 wire [0:0] _10158_;
 wire [0:0] _10159_;
 wire [0:0] _10160_;
 wire [0:0] _10161_;
 wire [0:0] _10162_;
 wire [0:0] _10163_;
 wire [0:0] _10164_;
 wire [0:0] _10165_;
 wire [0:0] _10166_;
 wire [0:0] _10167_;
 wire [0:0] _10168_;
 wire [0:0] _10169_;
 wire [0:0] _10170_;
 wire [0:0] _10171_;
 wire [0:0] _10172_;
 wire [0:0] _10173_;
 wire [0:0] _10174_;
 wire [0:0] _10175_;
 wire [0:0] _10176_;
 wire [0:0] _10177_;
 wire [0:0] _10178_;
 wire [0:0] _10179_;
 wire [0:0] _10180_;
 wire [0:0] _10181_;
 wire [0:0] _10182_;
 wire [0:0] _10183_;
 wire [0:0] _10184_;
 wire [0:0] _10185_;
 wire [0:0] _10186_;
 wire [0:0] _10187_;
 wire [0:0] _10188_;
 wire [0:0] _10189_;
 wire [0:0] _10190_;
 wire [0:0] _10191_;
 wire [0:0] _10192_;
 wire [0:0] _10193_;
 wire [0:0] _10194_;
 wire [0:0] _10195_;
 wire [0:0] _10196_;
 wire [0:0] _10197_;
 wire [0:0] _10198_;
 wire [0:0] _10199_;
 wire [0:0] _10200_;
 wire [0:0] _10201_;
 wire [0:0] _10202_;
 wire [0:0] _10203_;
 wire [0:0] _10204_;
 wire [0:0] _10205_;
 wire [0:0] _10206_;
 wire [0:0] _10207_;
 wire [0:0] _10208_;
 wire [0:0] _10209_;
 wire [0:0] _10210_;
 wire [0:0] _10211_;
 wire [0:0] _10212_;
 wire [0:0] _10213_;
 wire [0:0] _10214_;
 wire [0:0] _10215_;
 wire [0:0] _10216_;
 wire [0:0] _10217_;
 wire [0:0] _10218_;
 wire [0:0] _10219_;
 wire [0:0] _10220_;
 wire [0:0] _10221_;
 wire [0:0] _10222_;
 wire [0:0] _10223_;
 wire [0:0] _10224_;
 wire [0:0] _10225_;
 wire [0:0] _10226_;
 wire [0:0] _10227_;
 wire [0:0] _10228_;
 wire [0:0] _10229_;
 wire [0:0] _10230_;
 wire [0:0] _10231_;
 wire [0:0] _10232_;
 wire [0:0] _10233_;
 wire [0:0] _10234_;
 wire [0:0] _10235_;
 wire [0:0] _10236_;
 wire [0:0] _10237_;
 wire [0:0] _10238_;
 wire [0:0] _10239_;
 wire [0:0] _10240_;
 wire [0:0] _10241_;
 wire [0:0] _10242_;
 wire [0:0] _10243_;
 wire [0:0] _10244_;
 wire [0:0] _10245_;
 wire [0:0] _10246_;
 wire [0:0] _10247_;
 wire [0:0] _10248_;
 wire [0:0] _10249_;
 wire [0:0] _10250_;
 wire [0:0] _10251_;
 wire [0:0] _10252_;
 wire [0:0] _10253_;
 wire [0:0] _10254_;
 wire [0:0] _10255_;
 wire [0:0] _10256_;
 wire [0:0] _10257_;
 wire [0:0] _10258_;
 wire [0:0] _10259_;
 wire [0:0] _10260_;
 wire [0:0] _10261_;
 wire [0:0] _10262_;
 wire [0:0] _10263_;
 wire [0:0] _10264_;
 wire [0:0] _10265_;
 wire [0:0] _10266_;
 wire [0:0] _10267_;
 wire [0:0] _10268_;
 wire [0:0] _10269_;
 wire [0:0] _10270_;
 wire [0:0] _10271_;
 wire [0:0] _10272_;
 wire [0:0] _10273_;
 wire [0:0] _10274_;
 wire [0:0] _10275_;
 wire [0:0] _10276_;
 wire [0:0] _10277_;
 wire [0:0] _10278_;
 wire [0:0] _10279_;
 wire [0:0] _10280_;
 wire [0:0] _10281_;
 wire [0:0] _10282_;
 wire [0:0] _10283_;
 wire [0:0] _10284_;
 wire [0:0] _10285_;
 wire [0:0] _10286_;
 wire [0:0] _10287_;
 wire [0:0] _10288_;
 wire [0:0] _10289_;
 wire [0:0] _10290_;
 wire [0:0] _10291_;
 wire [0:0] _10292_;
 wire [0:0] _10293_;
 wire [0:0] _10294_;
 wire [0:0] _10295_;
 wire [0:0] _10296_;
 wire [0:0] _10297_;
 wire [0:0] _10298_;
 wire [0:0] _10299_;
 wire [0:0] _10300_;
 wire [0:0] _10301_;
 wire [0:0] _10302_;
 wire [0:0] _10303_;
 wire [0:0] _10304_;
 wire [0:0] _10305_;
 wire [0:0] _10306_;
 wire [0:0] _10307_;
 wire [0:0] _10308_;
 wire [0:0] _10309_;
 wire [0:0] _10310_;
 wire [0:0] _10311_;
 wire [0:0] _10312_;
 wire [0:0] _10313_;
 wire [0:0] _10314_;
 wire [0:0] _10315_;
 wire [0:0] _10316_;
 wire [0:0] _10317_;
 wire [0:0] _10318_;
 wire [0:0] _10319_;
 wire [0:0] _10320_;
 wire [0:0] _10321_;
 wire [0:0] _10322_;
 wire [0:0] _10323_;
 wire [0:0] _10324_;
 wire [0:0] _10325_;
 wire [0:0] _10326_;
 wire [0:0] _10327_;
 wire [0:0] _10328_;
 wire [0:0] _10329_;
 wire [0:0] _10330_;
 wire [0:0] _10331_;
 wire [0:0] _10332_;
 wire [0:0] _10333_;
 wire [0:0] _10334_;
 wire [0:0] _10335_;
 wire [0:0] _10336_;
 wire [0:0] _10337_;
 wire [0:0] _10338_;
 wire [0:0] _10339_;
 wire [0:0] _10340_;
 wire [0:0] _10341_;
 wire [0:0] _10342_;
 wire [0:0] _10343_;
 wire [0:0] _10344_;
 wire [0:0] _10345_;
 wire [0:0] _10346_;
 wire [0:0] _10347_;
 wire [0:0] _10348_;
 wire [0:0] _10349_;
 wire [0:0] _10350_;
 wire [0:0] _10351_;
 wire [0:0] _10352_;
 wire [0:0] _10353_;
 wire [0:0] _10354_;
 wire [0:0] _10355_;
 wire [0:0] _10356_;
 wire [0:0] _10357_;
 wire [0:0] _10358_;
 wire [0:0] _10359_;
 wire [0:0] _10360_;
 wire [0:0] _10361_;
 wire [0:0] _10362_;
 wire [0:0] _10363_;
 wire [0:0] _10364_;
 wire [0:0] _10365_;
 wire [0:0] _10366_;
 wire [0:0] _10367_;
 wire [0:0] _10368_;
 wire [0:0] _10369_;
 wire [0:0] _10370_;
 wire [0:0] _10371_;
 wire [0:0] _10372_;
 wire [0:0] _10373_;
 wire [0:0] _10374_;
 wire [0:0] _10375_;
 wire [0:0] _10376_;
 wire [0:0] _10377_;
 wire [0:0] _10378_;
 wire [0:0] _10379_;
 wire [0:0] _10380_;
 wire [0:0] _10381_;
 wire [0:0] _10382_;
 wire [0:0] _10383_;
 wire [0:0] _10384_;
 wire [0:0] _10385_;
 wire [0:0] _10386_;
 wire [0:0] _10387_;
 wire [0:0] _10388_;
 wire [0:0] _10389_;
 wire [0:0] _10390_;
 wire [0:0] _10391_;
 wire [0:0] _10392_;
 wire [0:0] _10393_;
 wire [0:0] _10394_;
 wire [0:0] _10395_;
 wire [0:0] _10396_;
 wire [0:0] _10397_;
 wire [0:0] _10398_;
 wire [0:0] _10399_;
 wire [0:0] _10400_;
 wire [0:0] _10401_;
 wire [0:0] _10402_;
 wire [0:0] _10403_;
 wire [0:0] _10404_;
 wire [0:0] _10405_;
 wire [0:0] _10406_;
 wire [0:0] _10407_;
 wire [0:0] _10408_;
 wire [0:0] _10409_;
 wire [0:0] _10410_;
 wire [0:0] _10411_;
 wire [0:0] _10412_;
 wire [0:0] _10413_;
 wire [0:0] _10414_;
 wire [0:0] _10415_;
 wire [0:0] _10416_;
 wire [0:0] _10417_;
 wire [0:0] _10418_;
 wire [0:0] _10419_;
 wire [0:0] _10420_;
 wire [0:0] _10421_;
 wire [0:0] _10422_;
 wire [0:0] _10423_;
 wire [0:0] _10424_;
 wire [0:0] _10425_;
 wire [0:0] _10426_;
 wire [0:0] _10427_;
 wire [0:0] _10428_;
 wire [0:0] _10429_;
 wire [0:0] _10430_;
 wire [0:0] _10431_;
 wire [0:0] _10432_;
 wire [0:0] _10433_;
 wire [0:0] _10434_;
 wire [0:0] _10435_;
 wire [0:0] _10436_;
 wire [0:0] _10437_;
 wire [0:0] _10438_;
 wire [0:0] _10439_;
 wire [0:0] _10440_;
 wire [0:0] _10441_;
 wire [0:0] _10442_;
 wire [0:0] _10443_;
 wire [0:0] _10444_;
 wire [0:0] _10445_;
 wire [0:0] _10446_;
 wire [0:0] _10447_;
 wire [0:0] _10448_;
 wire [0:0] _10449_;
 wire [0:0] _10450_;
 wire [0:0] _10451_;
 wire [0:0] _10452_;
 wire [0:0] _10453_;
 wire [0:0] _10454_;
 wire [0:0] _10455_;
 wire [0:0] _10456_;
 wire [0:0] _10457_;
 wire [0:0] _10458_;
 wire [0:0] _10459_;
 wire [0:0] _10460_;
 wire [0:0] _10461_;
 wire [0:0] _10462_;
 wire [0:0] _10463_;
 wire [0:0] _10464_;
 wire [0:0] _10465_;
 wire [0:0] _10466_;
 wire [0:0] _10467_;
 wire [0:0] _10468_;
 wire [0:0] _10469_;
 wire [0:0] _10470_;
 wire [0:0] _10471_;
 wire [0:0] _10472_;
 wire [0:0] _10473_;
 wire [0:0] _10474_;
 wire [0:0] _10475_;
 wire [0:0] _10476_;
 wire [0:0] _10477_;
 wire [0:0] _10478_;
 wire [0:0] _10479_;
 wire [0:0] _10480_;
 wire [0:0] _10481_;
 wire [0:0] _10482_;
 wire [0:0] _10483_;
 wire [0:0] _10484_;
 wire [0:0] _10485_;
 wire [0:0] _10486_;
 wire [0:0] _10487_;
 wire [0:0] _10488_;
 wire [0:0] _10489_;
 wire [0:0] _10490_;
 wire [0:0] _10491_;
 wire [0:0] _10492_;
 wire [0:0] _10493_;
 wire [0:0] _10494_;
 wire [0:0] _10495_;
 wire [0:0] _10496_;
 wire [0:0] _10497_;
 wire [0:0] _10498_;
 wire [0:0] _10499_;
 wire [0:0] _10500_;
 wire [0:0] _10501_;
 wire [0:0] _10502_;
 wire [0:0] _10503_;
 wire [0:0] _10504_;
 wire [0:0] _10505_;
 wire [0:0] _10506_;
 wire [0:0] _10507_;
 wire [0:0] _10508_;
 wire [0:0] _10509_;
 wire [0:0] _10510_;
 wire [0:0] _10511_;
 wire [0:0] _10512_;
 wire [0:0] _10513_;
 wire [0:0] _10514_;
 wire [0:0] _10515_;
 wire [0:0] _10516_;
 wire [0:0] _10517_;
 wire [0:0] _10518_;
 wire [0:0] _10519_;
 wire [0:0] _10520_;
 wire [0:0] _10521_;
 wire [0:0] _10522_;
 wire [0:0] _10523_;
 wire [0:0] _10524_;
 wire [0:0] _10525_;
 wire [0:0] _10526_;
 wire [0:0] _10527_;
 wire [0:0] _10528_;
 wire [0:0] _10529_;
 wire [0:0] _10530_;
 wire [0:0] _10531_;
 wire [0:0] _10532_;
 wire [0:0] _10533_;
 wire [0:0] _10534_;
 wire [0:0] _10535_;
 wire [0:0] _10536_;
 wire [0:0] _10537_;
 wire [0:0] _10538_;
 wire [0:0] _10539_;
 wire [0:0] _10540_;
 wire [0:0] _10541_;
 wire [0:0] _10542_;
 wire [0:0] _10543_;
 wire [0:0] _10544_;
 wire [0:0] _10545_;
 wire [0:0] _10546_;
 wire [0:0] _10547_;
 wire [0:0] _10548_;
 wire [0:0] _10549_;
 wire [0:0] _10550_;
 wire [0:0] _10551_;
 wire [0:0] _10552_;
 wire [0:0] _10553_;
 wire [0:0] _10554_;
 wire [0:0] _10555_;
 wire [0:0] _10556_;
 wire [0:0] _10557_;
 wire [0:0] _10558_;
 wire [0:0] _10559_;
 wire [0:0] _10560_;
 wire [0:0] _10561_;
 wire [0:0] _10562_;
 wire [0:0] _10563_;
 wire [0:0] _10564_;
 wire [0:0] _10565_;
 wire [0:0] _10566_;
 wire [0:0] _10567_;
 wire [0:0] _10568_;
 wire [0:0] _10569_;
 wire [0:0] _10570_;
 wire [0:0] _10571_;
 wire [0:0] _10572_;
 wire [0:0] _10573_;
 wire [0:0] _10574_;
 wire [0:0] _10575_;
 wire [0:0] _10576_;
 wire [0:0] _10577_;
 wire [0:0] _10578_;
 wire [0:0] _10579_;
 wire [0:0] _10580_;
 wire [0:0] _10581_;
 wire [0:0] _10582_;
 wire [0:0] _10583_;
 wire [0:0] _10584_;
 wire [0:0] _10585_;
 wire [0:0] _10586_;
 wire [0:0] _10587_;
 wire [0:0] _10588_;
 wire [0:0] _10589_;
 wire [0:0] _10590_;
 wire [0:0] _10591_;
 wire [0:0] _10592_;
 wire [0:0] _10593_;
 wire [0:0] _10594_;
 wire [0:0] _10595_;
 wire [0:0] _10596_;
 wire [0:0] _10597_;
 wire [0:0] _10598_;
 wire [0:0] _10599_;
 wire [0:0] _10600_;
 wire [0:0] _10601_;
 wire [0:0] _10602_;
 wire [0:0] _10603_;
 wire [0:0] _10604_;
 wire [0:0] _10605_;
 wire [0:0] _10606_;
 wire [0:0] _10607_;
 wire [0:0] _10608_;
 wire [0:0] _10609_;
 wire [0:0] _10610_;
 wire [0:0] _10611_;
 wire [0:0] _10612_;
 wire [0:0] _10613_;
 wire [0:0] _10614_;
 wire [0:0] _10615_;
 wire [0:0] _10616_;
 wire [0:0] _10617_;
 wire [0:0] _10618_;
 wire [0:0] _10619_;
 wire [0:0] _10620_;
 wire [0:0] _10621_;
 wire [0:0] _10622_;
 wire [0:0] _10623_;
 wire [0:0] _10624_;
 wire [0:0] _10625_;
 wire [0:0] _10626_;
 wire [0:0] _10627_;
 wire [0:0] _10628_;
 wire [0:0] _10629_;
 wire [0:0] _10630_;
 wire [0:0] _10631_;
 wire [0:0] _10632_;
 wire [0:0] _10633_;
 wire [0:0] _10634_;
 wire [0:0] _10635_;
 wire [0:0] _10636_;
 wire [0:0] _10637_;
 wire [0:0] _10638_;
 wire [0:0] _10639_;
 wire [0:0] _10640_;
 wire [0:0] _10641_;
 wire [0:0] _10642_;
 wire [0:0] _10643_;
 wire [0:0] _10644_;
 wire [0:0] _10645_;
 wire [0:0] _10646_;
 wire [0:0] _10647_;
 wire [0:0] _10648_;
 wire [0:0] _10649_;
 wire [0:0] _10650_;
 wire [0:0] _10651_;
 wire [0:0] _10652_;
 wire [0:0] _10653_;
 wire [0:0] _10654_;
 wire [0:0] _10655_;
 wire [0:0] _10656_;
 wire [0:0] _10657_;
 wire [0:0] _10658_;
 wire [0:0] _10659_;
 wire [0:0] _10660_;
 wire [0:0] _10661_;
 wire [0:0] _10662_;
 wire [0:0] _10663_;
 wire [0:0] _10664_;
 wire [0:0] _10665_;
 wire [0:0] _10666_;
 wire [0:0] _10667_;
 wire [0:0] _10668_;
 wire [0:0] _10669_;
 wire [0:0] _10670_;
 wire [0:0] _10671_;
 wire [0:0] _10672_;
 wire [0:0] _10673_;
 wire [0:0] _10674_;
 wire [0:0] _10675_;
 wire [0:0] _10676_;
 wire [0:0] _10677_;
 wire [0:0] _10678_;
 wire [0:0] _10679_;
 wire [0:0] _10680_;
 wire [0:0] _10681_;
 wire [0:0] _10682_;
 wire [0:0] _10683_;
 wire [0:0] _10684_;
 wire [0:0] _10685_;
 wire [0:0] _10686_;
 wire [0:0] _10687_;
 wire [0:0] _10688_;
 wire [0:0] _10689_;
 wire [0:0] _10690_;
 wire [0:0] _10691_;
 wire [0:0] _10692_;
 wire [0:0] _10693_;
 wire [0:0] _10694_;
 wire [0:0] _10695_;
 wire [0:0] _10696_;
 wire [0:0] _10697_;
 wire [0:0] _10698_;
 wire [0:0] _10699_;
 wire [0:0] _10700_;
 wire [0:0] _10701_;
 wire [0:0] _10702_;
 wire [0:0] _10703_;
 wire [0:0] _10704_;
 wire [0:0] _10705_;
 wire [0:0] _10706_;
 wire [0:0] _10707_;
 wire [0:0] _10708_;
 wire [0:0] _10709_;
 wire [0:0] _10710_;
 wire [0:0] _10711_;
 wire [0:0] _10712_;
 wire [0:0] _10713_;
 wire [0:0] _10714_;
 wire [0:0] _10715_;
 wire [0:0] _10716_;
 wire [0:0] _10717_;
 wire [0:0] _10718_;
 wire [0:0] _10719_;
 wire [0:0] _10720_;
 wire [0:0] _10721_;
 wire [0:0] _10722_;
 wire [0:0] _10723_;
 wire [0:0] _10724_;
 wire [0:0] _10725_;
 wire [0:0] _10726_;
 wire [0:0] _10727_;
 wire [0:0] _10728_;
 wire [0:0] _10729_;
 wire [0:0] _10730_;
 wire [0:0] _10731_;
 wire [0:0] _10732_;
 wire [0:0] _10733_;
 wire [0:0] _10734_;
 wire [0:0] _10735_;
 wire [0:0] _10736_;
 wire [0:0] _10737_;
 wire [0:0] _10738_;
 wire [0:0] _10739_;
 wire [0:0] _10740_;
 wire [0:0] _10741_;
 wire [0:0] _10742_;
 wire [0:0] _10743_;
 wire [0:0] _10744_;
 wire [0:0] _10745_;
 wire [0:0] _10746_;
 wire [0:0] _10747_;
 wire [0:0] _10748_;
 wire [0:0] _10749_;
 wire [0:0] _10750_;
 wire [0:0] _10751_;
 wire [0:0] _10752_;
 wire [0:0] _10753_;
 wire [0:0] _10754_;
 wire [0:0] _10755_;
 wire [0:0] _10756_;
 wire [0:0] _10757_;
 wire [0:0] _10758_;
 wire [0:0] _10759_;
 wire [0:0] _10760_;
 wire [0:0] _10761_;
 wire [0:0] _10762_;
 wire [0:0] _10763_;
 wire [0:0] _10764_;
 wire [0:0] _10765_;
 wire [0:0] _10766_;
 wire [0:0] _10767_;
 wire [0:0] _10768_;
 wire [0:0] _10769_;
 wire [0:0] _10770_;
 wire [0:0] _10771_;
 wire [0:0] _10772_;
 wire [0:0] _10773_;
 wire [0:0] _10774_;
 wire [0:0] _10775_;
 wire [0:0] _10776_;
 wire [0:0] _10777_;
 wire [0:0] _10778_;
 wire [0:0] _10779_;
 wire [0:0] _10780_;
 wire [0:0] _10781_;
 wire [0:0] _10782_;
 wire [0:0] _10783_;
 wire [0:0] _10784_;
 wire [0:0] _10785_;
 wire [0:0] _10786_;
 wire [0:0] _10787_;
 wire [0:0] _10788_;
 wire [0:0] _10789_;
 wire [0:0] _10790_;
 wire [0:0] _10791_;
 wire [0:0] _10792_;
 wire [0:0] _10793_;
 wire [0:0] _10794_;
 wire [0:0] _10795_;
 wire [0:0] _10796_;
 wire [0:0] _10797_;
 wire [0:0] _10798_;
 wire [0:0] _10799_;
 wire [0:0] _10800_;
 wire [0:0] _10801_;
 wire [0:0] _10802_;
 wire [0:0] _10803_;
 wire [0:0] _10804_;
 wire [0:0] _10805_;
 wire [0:0] _10806_;
 wire [0:0] _10807_;
 wire [0:0] _10808_;
 wire [0:0] _10809_;
 wire [0:0] _10810_;
 wire [0:0] _10811_;
 wire [0:0] _10812_;
 wire [0:0] _10813_;
 wire [0:0] _10814_;
 wire [0:0] _10815_;
 wire [0:0] _10816_;
 wire [0:0] _10817_;
 wire [0:0] _10818_;
 wire [0:0] _10819_;
 wire [0:0] _10820_;
 wire [0:0] _10821_;
 wire [0:0] _10822_;
 wire [0:0] _10823_;
 wire [0:0] _10824_;
 wire [0:0] _10825_;
 wire [0:0] _10826_;
 wire [0:0] _10827_;
 wire [0:0] _10828_;
 wire [0:0] _10829_;
 wire [0:0] _10830_;
 wire [0:0] _10831_;
 wire [0:0] _10832_;
 wire [0:0] _10833_;
 wire [0:0] _10834_;
 wire [0:0] _10835_;
 wire [0:0] _10836_;
 wire [0:0] _10837_;
 wire [0:0] _10838_;
 wire [0:0] _10839_;
 wire [0:0] _10840_;
 wire [0:0] _10841_;
 wire [0:0] _10842_;
 wire [0:0] _10843_;
 wire [0:0] _10844_;
 wire [0:0] _10845_;
 wire [0:0] _10846_;
 wire [0:0] _10847_;
 wire [0:0] _10848_;
 wire [0:0] _10849_;
 wire [0:0] _10850_;
 wire [0:0] _10851_;
 wire [0:0] _10852_;
 wire [0:0] _10853_;
 wire [0:0] _10854_;
 wire [0:0] _10855_;
 wire [0:0] _10856_;
 wire [0:0] _10857_;
 wire [0:0] _10858_;
 wire [0:0] _10859_;
 wire [0:0] _10860_;
 wire [0:0] _10861_;
 wire [0:0] _10862_;
 wire [0:0] _10863_;
 wire [0:0] _10864_;
 wire [0:0] _10865_;
 wire [0:0] _10866_;
 wire [0:0] _10867_;
 wire [0:0] _10868_;
 wire [0:0] _10869_;
 wire [0:0] _10870_;
 wire [0:0] _10871_;
 wire [0:0] _10872_;
 wire [0:0] _10873_;
 wire [0:0] _10874_;
 wire [0:0] _10875_;
 wire [0:0] _10876_;
 wire [0:0] _10877_;
 wire [0:0] _10878_;
 wire [0:0] _10879_;
 wire [0:0] _10880_;
 wire [0:0] _10881_;
 wire [0:0] _10882_;
 wire [0:0] _10883_;
 wire [0:0] _10884_;
 wire [0:0] _10885_;
 wire [0:0] _10886_;
 wire [0:0] _10887_;
 wire [0:0] _10888_;
 wire [0:0] _10889_;
 wire [0:0] _10890_;
 wire [0:0] _10891_;
 wire [0:0] _10892_;
 wire [0:0] _10893_;
 wire [0:0] _10894_;
 wire [0:0] _10895_;
 wire [0:0] _10896_;
 wire [0:0] _10897_;
 wire [0:0] _10898_;
 wire [0:0] _10899_;
 wire [0:0] _10900_;
 wire [0:0] _10901_;
 wire [0:0] _10902_;
 wire [0:0] _10903_;
 wire [0:0] _10904_;
 wire [0:0] _10905_;
 wire [0:0] _10906_;
 wire [0:0] _10907_;
 wire [0:0] _10908_;
 wire [0:0] _10909_;
 wire [0:0] _10910_;
 wire [0:0] _10911_;
 wire [0:0] _10912_;
 wire [0:0] _10913_;
 wire [0:0] _10914_;
 wire [0:0] _10915_;
 wire [0:0] _10916_;
 wire [0:0] _10917_;
 wire [0:0] _10918_;
 wire [0:0] _10919_;
 wire [0:0] _10920_;
 wire [0:0] _10921_;
 wire [0:0] _10922_;
 wire [0:0] _10923_;
 wire [0:0] _10924_;
 wire [0:0] _10925_;
 wire [0:0] _10926_;
 wire [0:0] _10927_;
 wire [0:0] _10928_;
 wire [0:0] _10929_;
 wire [0:0] _10930_;
 wire [0:0] _10931_;
 wire [0:0] _10932_;
 wire [0:0] _10933_;
 wire [0:0] _10934_;
 wire [0:0] _10935_;
 wire [0:0] _10936_;
 wire [0:0] _10937_;
 wire [0:0] _10938_;
 wire [0:0] _10939_;
 wire [0:0] _10940_;
 wire [0:0] _10941_;
 wire [0:0] _10942_;
 wire [0:0] _10943_;
 wire [0:0] _10944_;
 wire [0:0] _10945_;
 wire [0:0] _10946_;
 wire [0:0] _10947_;
 wire [0:0] _10948_;
 wire [0:0] _10949_;
 wire [0:0] _10950_;
 wire [0:0] _10951_;
 wire [0:0] _10952_;
 wire [0:0] _10953_;
 wire [0:0] _10954_;
 wire [0:0] _10955_;
 wire [0:0] _10956_;
 wire [0:0] _10957_;
 wire [0:0] _10958_;
 wire [0:0] _10959_;
 wire [0:0] _10960_;
 wire [0:0] _10961_;
 wire [0:0] _10962_;
 wire [0:0] _10963_;
 wire [0:0] _10964_;
 wire [0:0] _10965_;
 wire [0:0] _10966_;
 wire [0:0] _10967_;
 wire [0:0] _10968_;
 wire [0:0] _10969_;
 wire [0:0] _10970_;
 wire [0:0] _10971_;
 wire [0:0] _10972_;
 wire [0:0] _10973_;
 wire [0:0] _10974_;
 wire [0:0] _10975_;
 wire [0:0] _10976_;
 wire [0:0] _10977_;
 wire [0:0] _10978_;
 wire [0:0] _10979_;
 wire [0:0] _10980_;
 wire [0:0] _10981_;
 wire [0:0] _10982_;
 wire [0:0] _10983_;
 wire [0:0] _10984_;
 wire [0:0] _10985_;
 wire [0:0] _10986_;
 wire [0:0] _10987_;
 wire [0:0] _10988_;
 wire [0:0] _10989_;
 wire [0:0] _10990_;
 wire [0:0] _10991_;
 wire [0:0] _10992_;
 wire [0:0] _10993_;
 wire [0:0] _10994_;
 wire [0:0] _10995_;
 wire [0:0] _10996_;
 wire [0:0] _10997_;
 wire [0:0] _10998_;
 wire [0:0] _10999_;
 wire [0:0] _11000_;
 wire [0:0] _11001_;
 wire [0:0] _11002_;
 wire [0:0] _11003_;
 wire [0:0] _11004_;
 wire [0:0] _11005_;
 wire [0:0] _11006_;
 wire [0:0] _11007_;
 wire [0:0] _11008_;
 wire [0:0] _11009_;
 wire [0:0] _11010_;
 wire [0:0] _11011_;
 wire [0:0] _11012_;
 wire [0:0] _11013_;
 wire [0:0] _11014_;
 wire [0:0] _11015_;
 wire [0:0] _11016_;
 wire [0:0] _11017_;
 wire [0:0] _11018_;
 wire [0:0] _11019_;
 wire [0:0] _11020_;
 wire [0:0] _11021_;
 wire [0:0] _11022_;
 wire [0:0] _11023_;
 wire [0:0] _11024_;
 wire [0:0] _11025_;
 wire [0:0] _11026_;
 wire [0:0] _11027_;
 wire [0:0] _11028_;
 wire [0:0] _11029_;
 wire [0:0] _11030_;
 wire [0:0] _11031_;
 wire [0:0] _11032_;
 wire [0:0] _11033_;
 wire [0:0] _11034_;
 wire [0:0] _11035_;
 wire [0:0] _11036_;
 wire [0:0] _11037_;
 wire [0:0] _11038_;
 wire [0:0] _11039_;
 wire [0:0] _11040_;
 wire [0:0] _11041_;
 wire [0:0] _11042_;
 wire [0:0] _11043_;
 wire [0:0] _11044_;
 wire [0:0] _11045_;
 wire [0:0] _11046_;
 wire [0:0] _11047_;
 wire [0:0] _11048_;
 wire [0:0] _11049_;
 wire [0:0] _11050_;
 wire [0:0] _11051_;
 wire [0:0] _11052_;
 wire [0:0] _11053_;
 wire [0:0] _11054_;
 wire [0:0] _11055_;
 wire [0:0] _11056_;
 wire [0:0] _11057_;
 wire [0:0] _11058_;
 wire [0:0] _11059_;
 wire [0:0] _11060_;
 wire [0:0] _11061_;
 wire [0:0] _11062_;
 wire [0:0] _11063_;
 wire [0:0] _11064_;
 wire [0:0] _11065_;
 wire [0:0] _11066_;
 wire [0:0] _11067_;
 wire [0:0] _11068_;
 wire [0:0] _11069_;
 wire [0:0] _11070_;
 wire [0:0] _11071_;
 wire [0:0] _11072_;
 wire [0:0] _11073_;
 wire [0:0] _11074_;
 wire [0:0] _11075_;
 wire [0:0] _11076_;
 wire [0:0] _11077_;
 wire [0:0] _11078_;
 wire [0:0] _11079_;
 wire [0:0] _11080_;
 wire [0:0] _11081_;
 wire [0:0] _11082_;
 wire [0:0] _11083_;
 wire [0:0] _11084_;
 wire [0:0] _11085_;
 wire [0:0] _11086_;
 wire [0:0] _11087_;
 wire [0:0] _11088_;
 wire [0:0] _11089_;
 wire [0:0] _11090_;
 wire [0:0] _11091_;
 wire [0:0] _11092_;
 wire [0:0] _11093_;
 wire [0:0] _11094_;
 wire [0:0] _11095_;
 wire [0:0] _11096_;
 wire [0:0] _11097_;
 wire [0:0] _11098_;
 wire [0:0] _11099_;
 wire [0:0] _11100_;
 wire [0:0] _11101_;
 wire [0:0] _11102_;
 wire [0:0] _11103_;
 wire [0:0] _11104_;
 wire [0:0] _11105_;
 wire [0:0] _11106_;
 wire [0:0] _11107_;
 wire [0:0] _11108_;
 wire [0:0] _11109_;
 wire [0:0] _11110_;
 wire [0:0] _11111_;
 wire [0:0] _11112_;
 wire [0:0] _11113_;
 wire [0:0] _11114_;
 wire [0:0] _11115_;
 wire [0:0] _11116_;
 wire [0:0] _11117_;
 wire [0:0] _11118_;
 wire [0:0] _11119_;
 wire [0:0] _11120_;
 wire [0:0] _11121_;
 wire [0:0] _11122_;
 wire [0:0] _11123_;
 wire [0:0] _11124_;
 wire [0:0] _11125_;
 wire [0:0] _11126_;
 wire [0:0] _11127_;
 wire [0:0] _11128_;
 wire [0:0] _11129_;
 wire [0:0] _11130_;
 wire [0:0] _11131_;
 wire [0:0] _11132_;
 wire [0:0] _11133_;
 wire [0:0] _11134_;
 wire [0:0] _11135_;
 wire [0:0] _11136_;
 wire [0:0] _11137_;
 wire [0:0] _11138_;
 wire [0:0] _11139_;
 wire [0:0] _11140_;
 wire [0:0] _11141_;
 wire [0:0] _11142_;
 wire [0:0] _11143_;
 wire [0:0] _11144_;
 wire [0:0] _11145_;
 wire [0:0] _11146_;
 wire [0:0] _11147_;
 wire [0:0] _11148_;
 wire [0:0] _11149_;
 wire [0:0] _11150_;
 wire [0:0] _11151_;
 wire [0:0] _11152_;
 wire [0:0] _11154_;
 wire [0:0] _11155_;
 wire [0:0] _11156_;
 wire [0:0] _11157_;
 wire [0:0] _11158_;
 wire [0:0] _11159_;
 wire [0:0] _11160_;
 wire [0:0] _11161_;
 wire [0:0] _11162_;
 wire [0:0] _11163_;
 wire [0:0] _11164_;
 wire [0:0] _11165_;
 wire [0:0] _11166_;
 wire [0:0] _11167_;
 wire [0:0] _11168_;
 wire [0:0] _11169_;
 wire [0:0] _11170_;
 wire [0:0] _11171_;
 wire [0:0] _11172_;
 wire [0:0] _11173_;
 wire [0:0] _11174_;
 wire [0:0] _11175_;
 wire [0:0] _11176_;
 wire [0:0] _11177_;
 wire [0:0] _11178_;
 wire [0:0] _11179_;
 wire [0:0] _11180_;
 wire [0:0] _11181_;
 wire [0:0] _11182_;
 wire [0:0] _11183_;
 wire [0:0] _11184_;
 wire [0:0] _11185_;
 wire [0:0] _11186_;
 wire [0:0] _11187_;
 wire [0:0] _11188_;
 wire [0:0] _11189_;
 wire [0:0] _11190_;
 wire [0:0] _11191_;
 wire [0:0] _11192_;
 wire [0:0] _11193_;
 wire [0:0] _11194_;
 wire [0:0] _11195_;
 wire [0:0] _11196_;
 wire [0:0] _11197_;
 wire [0:0] _11198_;
 wire [0:0] _11199_;
 wire [0:0] _11200_;
 wire [0:0] _11201_;
 wire [0:0] _11202_;
 wire [0:0] _11203_;
 wire [0:0] _11204_;
 wire [0:0] _11205_;
 wire [0:0] _11206_;
 wire [0:0] _11207_;
 wire [0:0] _11208_;
 wire [0:0] _11209_;
 wire [0:0] _11210_;
 wire [0:0] _11211_;
 wire [0:0] _11212_;
 wire [0:0] _11213_;
 wire [0:0] _11214_;
 wire [0:0] _11215_;
 wire [0:0] _11216_;
 wire [0:0] _11217_;
 wire [0:0] _11218_;
 wire [0:0] _11219_;
 wire [0:0] _11220_;
 wire [0:0] _11221_;
 wire [0:0] _11222_;
 wire [0:0] _11223_;
 wire [0:0] _11224_;
 wire [0:0] _11225_;
 wire [0:0] _11226_;
 wire [0:0] _11227_;
 wire [0:0] _11228_;
 wire [0:0] _11229_;
 wire [0:0] _11230_;
 wire [0:0] _11231_;
 wire [0:0] _11232_;
 wire [0:0] _11233_;
 wire [0:0] _11234_;
 wire [0:0] _11235_;
 wire [0:0] _11236_;
 wire [0:0] _11237_;
 wire [0:0] _11238_;
 wire [0:0] _11239_;
 wire [0:0] _11240_;
 wire [0:0] _11241_;
 wire [0:0] _11242_;
 wire [0:0] _11243_;
 wire [0:0] _11244_;
 wire [0:0] _11245_;
 wire [0:0] _11246_;
 wire [0:0] _11247_;
 wire [0:0] _11248_;
 wire [0:0] _11249_;
 wire [0:0] _11250_;
 wire [0:0] _11251_;
 wire [0:0] _11252_;
 wire [0:0] _11253_;
 wire [0:0] _11254_;
 wire [0:0] _11255_;
 wire [0:0] _11256_;
 wire [0:0] _11257_;
 wire [0:0] _11258_;
 wire [0:0] _11259_;
 wire [0:0] _11260_;
 wire [0:0] _11261_;
 wire [0:0] _11262_;
 wire [0:0] _11263_;
 wire [0:0] _11264_;
 wire [0:0] _11265_;
 wire [0:0] _11266_;
 wire [0:0] _11267_;
 wire [0:0] _11268_;
 wire [0:0] _11269_;
 wire [0:0] _11270_;
 wire [0:0] _11271_;
 wire [0:0] _11272_;
 wire [0:0] _11273_;
 wire [0:0] _11274_;
 wire [0:0] _11275_;
 wire [0:0] _11276_;
 wire [0:0] _11277_;
 wire [0:0] _11278_;
 wire [0:0] _11279_;
 wire [0:0] _11280_;
 wire [0:0] _11281_;
 wire [0:0] _11282_;
 wire [0:0] _11283_;
 wire [0:0] _11284_;
 wire [0:0] _11285_;
 wire [0:0] _11286_;
 wire [0:0] _11287_;
 wire [0:0] _11288_;
 wire [0:0] _11289_;
 wire [0:0] _11290_;
 wire [0:0] _11291_;
 wire [0:0] _11292_;
 wire [0:0] _11293_;
 wire [0:0] _11294_;
 wire [0:0] _11295_;
 wire [0:0] _11296_;
 wire [0:0] _11297_;
 wire [0:0] _11298_;
 wire [0:0] _11299_;
 wire [0:0] _11300_;
 wire [0:0] _11301_;
 wire [0:0] _11302_;
 wire [0:0] _11303_;
 wire [0:0] _11304_;
 wire [0:0] _11305_;
 wire [0:0] _11306_;
 wire [0:0] _11307_;
 wire [0:0] _11308_;
 wire [0:0] _11309_;
 wire [0:0] _11310_;
 wire [0:0] _11311_;
 wire [0:0] _11312_;
 wire [0:0] _11313_;
 wire [0:0] _11314_;
 wire [0:0] _11315_;
 wire [0:0] _11316_;
 wire [0:0] _11317_;
 wire [0:0] _11318_;
 wire [0:0] _11319_;
 wire [0:0] _11320_;
 wire [0:0] _11321_;
 wire [0:0] _11322_;
 wire [0:0] _11323_;
 wire [0:0] _11324_;
 wire [0:0] _11325_;
 wire [0:0] _11326_;
 wire [0:0] _11327_;
 wire [0:0] _11328_;
 wire [0:0] _11329_;
 wire [0:0] _11330_;
 wire [0:0] _11331_;
 wire [0:0] _11332_;
 wire [0:0] _11333_;
 wire [0:0] _11334_;
 wire [0:0] _11335_;
 wire [0:0] _11336_;
 wire [0:0] _11337_;
 wire [0:0] _11338_;
 wire [0:0] _11339_;
 wire [0:0] _11340_;
 wire [0:0] _11341_;
 wire [0:0] _11342_;
 wire [0:0] _11343_;
 wire [0:0] _11344_;
 wire [0:0] _11345_;
 wire [0:0] _11346_;
 wire [0:0] _11347_;
 wire [0:0] _11348_;
 wire [0:0] _11349_;
 wire [0:0] _11350_;
 wire [0:0] _11351_;
 wire [0:0] _11352_;
 wire [0:0] _11353_;
 wire [0:0] _11354_;
 wire [0:0] _11355_;
 wire [0:0] _11356_;
 wire [0:0] _11357_;
 wire [0:0] _11358_;
 wire [0:0] _11359_;
 wire [0:0] _11360_;
 wire [0:0] _11361_;
 wire [0:0] _11362_;
 wire [0:0] _11363_;
 wire [0:0] _11364_;
 wire [0:0] _11365_;
 wire [0:0] _11366_;
 wire [0:0] _11367_;
 wire [0:0] _11368_;
 wire [0:0] _11369_;
 wire [0:0] _11370_;
 wire [0:0] _11371_;
 wire [0:0] _11372_;
 wire [0:0] _11373_;
 wire [0:0] _11374_;
 wire [0:0] _11375_;
 wire [0:0] _11376_;
 wire [0:0] _11377_;
 wire [0:0] _11378_;
 wire [0:0] _11379_;
 wire [0:0] _11380_;
 wire [0:0] _11381_;
 wire [0:0] _11382_;
 wire [0:0] _11383_;
 wire [0:0] _11384_;
 wire [0:0] _11385_;
 wire [0:0] _11386_;
 wire [0:0] _11387_;
 wire [0:0] _11388_;
 wire [0:0] _11389_;
 wire [0:0] _11390_;
 wire [0:0] _11391_;
 wire [0:0] _11393_;
 wire [0:0] _11394_;
 wire [0:0] _11395_;
 wire [0:0] _11397_;
 wire [0:0] _11398_;
 wire [0:0] _11399_;
 wire [0:0] _11400_;
 wire [0:0] _11401_;
 wire [0:0] _11402_;
 wire [0:0] _11404_;
 wire [0:0] _11405_;
 wire [0:0] _11406_;
 wire [0:0] _11407_;
 wire [0:0] _11408_;
 wire [0:0] _11409_;
 wire [0:0] _11410_;
 wire [0:0] _11411_;
 wire [0:0] _11412_;
 wire [0:0] _11413_;
 wire [0:0] _11414_;
 wire [0:0] _11415_;
 wire [0:0] _11416_;
 wire [0:0] _11417_;
 wire [0:0] _11418_;
 wire [0:0] _11419_;
 wire [0:0] _11420_;
 wire [0:0] _11421_;
 wire [0:0] _11422_;
 wire [0:0] _11423_;
 wire [0:0] _11424_;
 wire [0:0] _11425_;
 wire [0:0] _11427_;
 wire [0:0] _11428_;
 wire [0:0] _11429_;
 wire [0:0] _11430_;
 wire [0:0] _11431_;
 wire [0:0] _11432_;
 wire [0:0] _11433_;
 wire [0:0] _11434_;
 wire [0:0] _11435_;
 wire [0:0] _11436_;
 wire [0:0] _11437_;
 wire [0:0] _11438_;
 wire [0:0] _11439_;
 wire [0:0] _11440_;
 wire [0:0] _11441_;
 wire [0:0] _11442_;
 wire [0:0] _11443_;
 wire [0:0] _11444_;
 wire [0:0] _11445_;
 wire [0:0] _11446_;
 wire [0:0] _11447_;
 wire [0:0] _11448_;
 wire [0:0] _11449_;
 wire [0:0] _11450_;
 wire [0:0] _11451_;
 wire [0:0] _11452_;
 wire [0:0] _11453_;
 wire [0:0] _11454_;
 wire [0:0] _11455_;
 wire [0:0] _11456_;
 wire [0:0] _11457_;
 wire [0:0] _11458_;
 wire [0:0] _11459_;
 wire [0:0] _11460_;
 wire [0:0] _11461_;
 wire [0:0] _11462_;
 wire [0:0] _11463_;
 wire [0:0] _11464_;
 wire [0:0] _11465_;
 wire [0:0] _11466_;
 wire [0:0] _11467_;
 wire [0:0] _11468_;
 wire [0:0] _11469_;
 wire [0:0] _11470_;
 wire [0:0] _11471_;
 wire [0:0] _11472_;
 wire [0:0] _11473_;
 wire [0:0] _11474_;
 wire [0:0] _11475_;
 wire [0:0] _11476_;
 wire [0:0] _11477_;
 wire [0:0] _11478_;
 wire [0:0] _11479_;
 wire [0:0] _11480_;
 wire [0:0] _11481_;
 wire [0:0] _11482_;
 wire [0:0] _11483_;
 wire [0:0] _11484_;
 wire [0:0] _11485_;
 wire [0:0] _11486_;
 wire [0:0] _11487_;
 wire [0:0] _11488_;
 wire [0:0] _11489_;
 wire [0:0] _11490_;
 wire [0:0] _11491_;
 wire [0:0] _11492_;
 wire [0:0] _11493_;
 wire [0:0] _11494_;
 wire [0:0] _11495_;
 wire [0:0] _11496_;
 wire [0:0] _11497_;
 wire [0:0] _11498_;
 wire [0:0] _11499_;
 wire [0:0] _11500_;
 wire [0:0] _11501_;
 wire [0:0] _11502_;
 wire [0:0] _11503_;
 wire [0:0] _11504_;
 wire [0:0] _11505_;
 wire [0:0] _11506_;
 wire [0:0] _11507_;
 wire [0:0] _11508_;
 wire [0:0] _11509_;
 wire [0:0] _11510_;
 wire [0:0] _11511_;
 wire [0:0] _11512_;
 wire [0:0] _11513_;
 wire [0:0] _11514_;
 wire [0:0] _11515_;
 wire [0:0] _11516_;
 wire [0:0] _11517_;
 wire [0:0] _11518_;
 wire [0:0] _11519_;
 wire [0:0] _11520_;
 wire [0:0] _11521_;
 wire [0:0] _11522_;
 wire [0:0] _11523_;
 wire [0:0] _11524_;
 wire [0:0] _11525_;
 wire [0:0] _11526_;
 wire [0:0] _11527_;
 wire [0:0] _11528_;
 wire [0:0] _11529_;
 wire [0:0] _11530_;
 wire [0:0] _11531_;
 wire [0:0] _11532_;
 wire [0:0] _11533_;
 wire [0:0] _11534_;
 wire [0:0] _11535_;
 wire [0:0] _11536_;
 wire [0:0] _11537_;
 wire [0:0] _11538_;
 wire [0:0] _11539_;
 wire [0:0] _11540_;
 wire [0:0] _11541_;
 wire [0:0] _11542_;
 wire [0:0] _11543_;
 wire [0:0] _11544_;
 wire [0:0] _11545_;
 wire [0:0] _11546_;
 wire [0:0] _11547_;
 wire [0:0] _11548_;
 wire [0:0] _11549_;
 wire [0:0] _11550_;
 wire [0:0] _11551_;
 wire [0:0] _11552_;
 wire [0:0] _11553_;
 wire [0:0] _11554_;
 wire [0:0] _11555_;
 wire [0:0] _11556_;
 wire [0:0] _11557_;
 wire [0:0] _11558_;
 wire [0:0] _11559_;
 wire [0:0] _11560_;
 wire [0:0] _11561_;
 wire [0:0] _11562_;
 wire [0:0] _11563_;
 wire [0:0] _11564_;
 wire [0:0] _11565_;
 wire [0:0] _11566_;
 wire [0:0] _11567_;
 wire [0:0] _11568_;
 wire [0:0] _11569_;
 wire [0:0] _11570_;
 wire [0:0] _11571_;
 wire [0:0] _11572_;
 wire [0:0] _11573_;
 wire [0:0] _11574_;
 wire [0:0] _11575_;
 wire [0:0] _11576_;
 wire [0:0] _11577_;
 wire [0:0] _11578_;
 wire [0:0] _11579_;
 wire [0:0] _11580_;
 wire [0:0] _11581_;
 wire [0:0] _11582_;
 wire [0:0] _11583_;
 wire [0:0] _11584_;
 wire [0:0] _11585_;
 wire [0:0] _11586_;
 wire [0:0] _11587_;
 wire [0:0] _11588_;
 wire [0:0] _11589_;
 wire [0:0] _11590_;
 wire [0:0] _11591_;
 wire [0:0] _11592_;
 wire [0:0] _11593_;
 wire [0:0] _11594_;
 wire [0:0] _11595_;
 wire [0:0] _11596_;
 wire [0:0] _11597_;
 wire [0:0] _11598_;
 wire [0:0] _11599_;
 wire [0:0] _11600_;
 wire [0:0] _11601_;
 wire [0:0] _11602_;
 wire [0:0] _11603_;
 wire [0:0] _11604_;
 wire [0:0] _11605_;
 wire [0:0] _11606_;
 wire [0:0] _11607_;
 wire [0:0] _11608_;
 wire [0:0] _11609_;
 wire [0:0] _11610_;
 wire [0:0] _11611_;
 wire [0:0] _11612_;
 wire [0:0] _11613_;
 wire [0:0] _11614_;
 wire [0:0] _11615_;
 wire [0:0] _11616_;
 wire [0:0] _11617_;
 wire [0:0] _11618_;
 wire [0:0] _11619_;
 wire [0:0] _11620_;
 wire [0:0] _11621_;
 wire [0:0] _11622_;
 wire [0:0] _11623_;
 wire [0:0] _11624_;
 wire [0:0] _11625_;
 wire [0:0] _11626_;
 wire [0:0] _11627_;
 wire [0:0] _11628_;
 wire [0:0] _11629_;
 wire [0:0] _11630_;
 wire [0:0] _11631_;
 wire [0:0] _11632_;
 wire [0:0] _11633_;
 wire [0:0] _11634_;
 wire [0:0] _11635_;
 wire [0:0] _11636_;
 wire [0:0] _11637_;
 wire [0:0] _11638_;
 wire [0:0] _11639_;
 wire [0:0] _11640_;
 wire [0:0] _11641_;
 wire [0:0] _11643_;
 wire [0:0] _11644_;
 wire [0:0] _11645_;
 wire [0:0] _11646_;
 wire [0:0] _11647_;
 wire [0:0] _11648_;
 wire [0:0] _11649_;
 wire [0:0] _11650_;
 wire [0:0] _11651_;
 wire [0:0] _11652_;
 wire [0:0] _11653_;
 wire [0:0] _11654_;
 wire [0:0] _11655_;
 wire [0:0] _11656_;
 wire [0:0] _11657_;
 wire [0:0] _11658_;
 wire [0:0] _11659_;
 wire [0:0] _11660_;
 wire [0:0] _11661_;
 wire [0:0] _11662_;
 wire [0:0] _11663_;
 wire [0:0] _11664_;

 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11666_ (.I(\load_store_unit_i.handle_misaligned_q ),
    .ZN(_11641_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11667_ (.A1(\id_stage_i.controller_i.instr_i[0] ),
    .A2(\id_stage_i.controller_i.instr_i[1] ),
    .Z(_06198_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3473 (.I(\id_stage_i.controller_i.instr_valid_i ),
    .Z(net3473));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3480 (.I(\id_stage_i.controller_i.instr_i[30] ),
    .Z(net3480));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3528 (.I(net3526),
    .Z(net3528));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11671_ (.A1(\id_stage_i.controller_i.instr_i[3] ),
    .A2(\id_stage_i.controller_i.instr_i[2] ),
    .ZN(_06202_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3527 (.I(net3526),
    .Z(net3527));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3478 (.I(\id_stage_i.controller_i.instr_i[3] ),
    .Z(net3478));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11674_ (.A1(net3474),
    .A2(net3476),
    .Z(_06205_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11675_ (.A1(net357),
    .A2(net3469),
    .A3(net390),
    .A4(_06205_),
    .Z(_06206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11676_ (.A1(net3646),
    .A2(_06206_),
    .ZN(_06207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11677_ (.A1(net3469),
    .A2(_06207_),
    .Z(_06208_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3475 (.I(\id_stage_i.controller_i.instr_i[5] ),
    .Z(net3475));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _11679_ (.I(\id_stage_i.controller_i.instr_i[4] ),
    .ZN(_06210_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3555 (.I(net3554),
    .Z(net3555));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11681_ (.A1(\id_stage_i.controller_i.instr_i[5] ),
    .A2(\id_stage_i.controller_i.instr_i[6] ),
    .ZN(_06212_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11682_ (.A1(net3478),
    .A2(_06212_),
    .A3(_06210_),
    .Z(_06213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11683_ (.A1(\id_stage_i.controller_i.instr_i[6] ),
    .A2(\id_stage_i.controller_i.instr_i[5] ),
    .Z(_06214_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11684_ (.A1(_06210_),
    .A2(net274),
    .Z(_06215_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3559 (.I(net3558),
    .Z(net3559));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11686_ (.A1(_06213_),
    .A2(_06215_),
    .B(net3481),
    .ZN(_06217_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_63_clk_i_regs (.I(clknet_6_60__leaf_clk_i_regs),
    .Z(clknet_leaf_63_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11688_ (.A1(net3476),
    .A2(net322),
    .Z(_06219_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11689_ (.I(net3475),
    .ZN(_06220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11690_ (.A1(net3474),
    .A2(_06220_),
    .B(net3481),
    .ZN(_06221_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11691_ (.I(net3478),
    .ZN(_06222_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11692_ (.A1(_06219_),
    .A2(_06221_),
    .B(_06222_),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11693_ (.A1(net3481),
    .A2(net3469),
    .Z(_06224_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3558 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(net3558));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3471 (.I(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(net3471));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11696_ (.A1(\id_stage_i.controller_i.instr_i[13] ),
    .A2(\id_stage_i.controller_i.instr_i[14] ),
    .Z(_06227_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11697_ (.A1(_06224_),
    .A2(_06213_),
    .A3(_06227_),
    .Z(_06228_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11698_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(\load_store_unit_i.ls_fsm_cs[1] ),
    .ZN(_06229_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11699_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_06229_),
    .ZN(_06230_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11700_ (.I(\load_store_unit_i.ls_fsm_cs[0] ),
    .ZN(_06231_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11701_ (.I(\load_store_unit_i.ls_fsm_cs[2] ),
    .ZN(_06232_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _11702_ (.A1(_06231_),
    .A2(\load_store_unit_i.handle_misaligned_q ),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .C(_06232_),
    .ZN(_06233_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11703_ (.A1(_06230_),
    .A2(_06233_),
    .ZN(_06234_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_62_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_62_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11705_ (.A1(_06217_),
    .A2(_06223_),
    .B(_06228_),
    .C(_06234_),
    .ZN(_06236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11706_ (.A1(_06208_),
    .A2(_06236_),
    .B(net3394),
    .ZN(_06237_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3645 (.I(net3644),
    .Z(net3645));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3526 (.I(net3513),
    .Z(net3526));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11709_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[12] ),
    .ZN(_06240_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _11710_ (.A1(net3478),
    .A2(_06210_),
    .A3(net322),
    .ZN(_06241_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11711_ (.I(net3649),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11712_ (.A1(\id_stage_i.controller_i.instr_i[13] ),
    .A2(\id_stage_i.controller_i.instr_i[14] ),
    .ZN(_06243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11713_ (.A1(_06242_),
    .A2(_06243_),
    .Z(_06244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11714_ (.A1(_06210_),
    .A2(net274),
    .ZN(_06245_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11715_ (.I(\id_stage_i.id_fsm_q ),
    .ZN(_06246_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11716_ (.A1(_06222_),
    .A2(net3473),
    .A3(_06246_),
    .Z(_06247_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11717_ (.A1(_06222_),
    .A2(net3477),
    .A3(net322),
    .ZN(_06248_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11718_ (.A1(_06241_),
    .A2(_06244_),
    .B1(_06245_),
    .B2(_06247_),
    .C(_06248_),
    .ZN(_06249_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11719_ (.A1(net3481),
    .A2(_06210_),
    .Z(_06250_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11720_ (.A1(net3478),
    .A2(net323),
    .A3(_06250_),
    .ZN(_06251_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11721_ (.A1(_06215_),
    .A2(_06221_),
    .B(_06222_),
    .ZN(_06252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11722_ (.A1(net3473),
    .A2(_06246_),
    .ZN(_06253_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11723_ (.A1(_06214_),
    .A2(_06198_),
    .A3(_06202_),
    .A4(_06210_),
    .Z(_06254_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11724_ (.A1(_06253_),
    .A2(net344),
    .Z(_06255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _11725_ (.A1(_06224_),
    .A2(_06249_),
    .B1(_06251_),
    .B2(_06252_),
    .C(_06255_),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11726_ (.A1(_06208_),
    .A2(_06256_),
    .ZN(_06257_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3537 (.I(net3534),
    .Z(net3537));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11728_ (.A1(_06237_),
    .A2(_06240_),
    .B(net3352),
    .ZN(_06259_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3577 (.I(net3576),
    .Z(net3577));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_57_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_57_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_56_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_56_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3587 (.I(net3583),
    .Z(net3587));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_1_0__f_clk_i (.I(clknet_0_clk_i),
    .Z(clknet_1_0__leaf_clk_i));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk_i_regs (.I(clknet_6_29__leaf_clk_i_regs),
    .Z(clknet_leaf_3_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk_i_regs (.I(clknet_6_29__leaf_clk_i_regs),
    .Z(clknet_leaf_2_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3608 (.I(net333),
    .Z(net3608));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11737_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S0(net3640),
    .S1(net3600),
    .Z(_06268_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk_i_regs (.I(clknet_6_29__leaf_clk_i_regs),
    .Z(clknet_leaf_1_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_54_clk_i_regs (.I(clknet_6_55__leaf_clk_i_regs),
    .Z(clknet_leaf_54_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11740_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(net3640),
    .Z(_06271_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3525 (.I(net423),
    .Z(net3525));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3513 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .Z(net3513));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11743_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .A2(net3640),
    .Z(_06274_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11744_ (.I(net3589),
    .ZN(_06275_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3502 (.I(net3500),
    .Z(net3502));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11746_ (.I0(_06271_),
    .I1(_06274_),
    .S(net3468),
    .Z(_06277_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3470 (.I(\load_store_unit_i.rdata_offset_q[1] ),
    .Z(net3470));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3505 (.I(net3503),
    .Z(net3505));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3491 (.I(net3490),
    .Z(net3491));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3512 (.I(net3509),
    .Z(net3512));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11751_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S0(net3640),
    .S1(net3600),
    .Z(_06282_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11752_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S0(net3640),
    .S1(net3600),
    .Z(_06283_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11753_ (.I(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .ZN(_06284_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3524 (.I(net314),
    .Z(net3524));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_53_clk_i_regs (.I(clknet_6_55__leaf_clk_i_regs),
    .Z(clknet_leaf_53_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3536 (.I(net3534),
    .Z(net3536));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3664 (.I(net3663),
    .Z(net3664));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _11758_ (.I0(_06268_),
    .I1(_06277_),
    .I2(_06282_),
    .I3(_06283_),
    .S0(net3459),
    .S1(net3579),
    .Z(_06289_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _11759_ (.I(net3576),
    .ZN(_06290_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3619 (.I(net3606),
    .Z(net3619));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3663 (.I(net3661),
    .Z(net3663));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3508 (.I(net3507),
    .Z(net3508));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3507 (.I(net3505),
    .Z(net3507));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3511 (.I(net3509),
    .Z(net3511));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3492 (.I(net3490),
    .Z(net3492));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11766_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S0(net3645),
    .S1(net3602),
    .Z(_06297_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11767_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S0(net3645),
    .S1(net3602),
    .Z(_06298_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3489 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .Z(net3489));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3501 (.I(net3500),
    .Z(net3501));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3500 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(net3500));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11771_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S0(net3640),
    .S1(net3597),
    .Z(_06302_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11772_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S0(net3640),
    .S1(net3597),
    .Z(_06303_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3499 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(net3499));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3510 (.I(net3509),
    .Z(net3510));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3618 (.I(net3616),
    .Z(net3618));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11776_ (.I0(_06297_),
    .I1(_06298_),
    .I2(_06302_),
    .I3(_06303_),
    .S0(net3461),
    .S1(net3578),
    .Z(_06307_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11777_ (.A1(_06290_),
    .A2(_06307_),
    .Z(_06308_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11778_ (.A1(net3577),
    .A2(_06289_),
    .B(_06308_),
    .ZN(_06309_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11779_ (.A1(_06208_),
    .A2(_06256_),
    .A3(_06236_),
    .Z(_06310_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3535 (.I(net3534),
    .Z(net3535));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11781_ (.A1(net3381),
    .A2(_06310_),
    .ZN(_06312_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11782_ (.A1(_06208_),
    .A2(_06236_),
    .Z(_06313_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_51_clk_i_regs (.I(clknet_6_55__leaf_clk_i_regs),
    .Z(clknet_leaf_51_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11784_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(_06313_),
    .Z(_06315_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11785_ (.A1(_06259_),
    .A2(_06312_),
    .A3(_06315_),
    .Z(_11494_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11786_ (.I(_11494_[0]),
    .ZN(_11490_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11787_ (.A1(_06213_),
    .A2(_06215_),
    .B(_06224_),
    .ZN(_06316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11788_ (.A1(net3469),
    .A2(_06202_),
    .Z(_06317_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11789_ (.A1(net3475),
    .A2(_06210_),
    .Z(_06318_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11790_ (.I(net277),
    .ZN(_06319_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11791_ (.A1(_06222_),
    .A2(_06319_),
    .A3(net3477),
    .A4(net270),
    .Z(_06320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11792_ (.A1(_06317_),
    .A2(_06318_),
    .B1(_06320_),
    .B2(net3481),
    .ZN(_06321_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11793_ (.A1(_06316_),
    .A2(_06321_),
    .B(_06234_),
    .ZN(_06322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11794_ (.A1(net3481),
    .A2(net270),
    .ZN(_06323_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11795_ (.A1(net320),
    .A2(_06243_),
    .Z(_06324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11796_ (.A1(_06215_),
    .A2(_06253_),
    .B1(_06324_),
    .B2(_06213_),
    .ZN(_06325_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11797_ (.A1(net3481),
    .A2(net3646),
    .Z(_06326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11798_ (.A1(net3481),
    .A2(net3477),
    .ZN(_06327_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11799_ (.A1(_06220_),
    .A2(net3477),
    .A3(_06326_),
    .B(_06327_),
    .ZN(_06328_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11800_ (.A1(_06222_),
    .A2(_06319_),
    .A3(net270),
    .Z(_06329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11801_ (.A1(_06328_),
    .A2(_06329_),
    .ZN(_06330_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11802_ (.A1(_06323_),
    .A2(_06325_),
    .B(_06330_),
    .ZN(_06331_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11803_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .A2(_06322_),
    .A3(_06331_),
    .Z(_06332_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3586 (.I(net3583),
    .Z(net3586));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _11805_ (.I(net3558),
    .ZN(_06334_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3465 (.I(_06275_),
    .Z(net3465));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11808_ (.A1(_06322_),
    .A2(_06331_),
    .B(net3449),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11809_ (.A1(_06253_),
    .A2(net262),
    .ZN(_06338_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3557 (.I(net3556),
    .Z(net3557));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11811_ (.I(\load_store_unit_i.ls_fsm_cs[1] ),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11812_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_11641_[0]),
    .B(_06340_),
    .C(\load_store_unit_i.ls_fsm_cs[2] ),
    .ZN(_06341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _11813_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_06229_),
    .B1(_06320_),
    .B2(net3481),
    .C(_06341_),
    .ZN(_06342_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11814_ (.A1(_06338_),
    .A2(_06342_),
    .Z(_06343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11815_ (.A1(net320),
    .A2(_06243_),
    .ZN(_06344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11816_ (.I(net3473),
    .ZN(_06345_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _11817_ (.A1(_06345_),
    .A2(net275),
    .B(_06214_),
    .C(_06210_),
    .ZN(_06346_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _11818_ (.A1(_06222_),
    .A2(_06245_),
    .B1(_06344_),
    .B2(_06241_),
    .C(_06346_),
    .ZN(_06347_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _11819_ (.A1(_06319_),
    .A2(net3476),
    .A3(_06345_),
    .A4(net275),
    .Z(_06348_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11820_ (.A1(net3476),
    .A2(net3646),
    .B(_06319_),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _11821_ (.A1(net3475),
    .A2(net3469),
    .A3(net266),
    .ZN(_06350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11822_ (.A1(_06348_),
    .A2(_06349_),
    .B(_06350_),
    .ZN(_06351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11823_ (.A1(_06224_),
    .A2(_06347_),
    .B(_06351_),
    .C(_06234_),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11824_ (.A1(_06332_),
    .A2(_06337_),
    .B(_06343_),
    .C(_06352_),
    .ZN(_06353_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11825_ (.A1(_06230_),
    .A2(_06233_),
    .Z(_06354_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11826_ (.A1(_06354_),
    .A2(_06351_),
    .Z(_06355_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3477 (.I(\id_stage_i.controller_i.instr_i[4] ),
    .Z(net3477));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3469 (.I(net268),
    .Z(net3469));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3644 (.I(net3606),
    .Z(net3644));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_67_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_67_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11831_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S0(net3529),
    .S1(net3510),
    .Z(_06360_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11832_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .S0(net3529),
    .S1(net3510),
    .Z(_06361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11833_ (.I0(_06360_),
    .I1(_06361_),
    .S(net3453),
    .Z(_06362_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_65_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_65_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3523 (.I(net3521),
    .Z(net3523));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11836_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S0(net3565),
    .S1(net3529),
    .Z(_06365_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11837_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .S0(net3565),
    .S1(net3529),
    .Z(_06366_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _11838_ (.I(net3503),
    .ZN(_06367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11839_ (.I0(_06365_),
    .I1(_06366_),
    .S(net3427),
    .Z(_06368_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11840_ (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .ZN(_06369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11841_ (.I0(_06362_),
    .I1(_06368_),
    .S(net3425),
    .Z(_06370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11842_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .S(net3530),
    .Z(_06371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11843_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S(net3530),
    .Z(_06372_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11844_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .A2(net3530),
    .Z(_06373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11845_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(net3530),
    .Z(_06374_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3495 (.I(net3490),
    .Z(net3495));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11847_ (.I0(_06371_),
    .I1(_06372_),
    .I2(_06373_),
    .I3(_06374_),
    .S0(net3563),
    .S1(net3427),
    .Z(_06376_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11848_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S0(net3529),
    .S1(net3510),
    .Z(_06377_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11849_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .S0(net3529),
    .S1(net3510),
    .Z(_06378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11850_ (.I0(_06377_),
    .I1(_06378_),
    .S(net3453),
    .Z(_06379_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3522 (.I(net3521),
    .Z(net3522));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11852_ (.I0(_06376_),
    .I1(_06379_),
    .S(net3491),
    .Z(_06381_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11853_ (.I(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .ZN(_06382_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk_i_regs (.I(clknet_6_23__leaf_clk_i_regs),
    .Z(clknet_leaf_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _11855_ (.I0(_06370_),
    .I1(_06381_),
    .S(net3423),
    .Z(_06384_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_49_clk_i_regs (.I(clknet_6_60__leaf_clk_i_regs),
    .Z(clknet_leaf_49_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11857_ (.A1(_06355_),
    .A2(_06384_),
    .ZN(_06386_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11858_ (.A1(_06353_),
    .A2(_06386_),
    .Z(_06387_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _11859_ (.I(_06387_),
    .ZN(_06388_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_48_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_48_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3521 (.I(net3513),
    .Z(net3521));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_47_clk_i_regs (.I(clknet_6_60__leaf_clk_i_regs),
    .Z(clknet_leaf_47_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3520 (.I(net423),
    .Z(net3520));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11864_ (.I(net3481),
    .ZN(_06391_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11865_ (.A1(\id_stage_i.controller_i.instr_i[0] ),
    .A2(\id_stage_i.controller_i.instr_i[1] ),
    .ZN(_06392_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _11866_ (.A1(net3478),
    .A2(net3474),
    .A3(_06210_),
    .A4(_06392_),
    .Z(_06393_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _11867_ (.A1(_06391_),
    .A2(_06393_),
    .B(_06233_),
    .C(_06230_),
    .ZN(_06394_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11868_ (.A1(_06230_),
    .A2(_06233_),
    .A3(_06328_),
    .A4(_06329_),
    .Z(_06395_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11869_ (.A1(_06255_),
    .A2(_06394_),
    .B(_06395_),
    .ZN(_06396_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11870_ (.A1(_06255_),
    .A2(_06394_),
    .A3(_06395_),
    .Z(_06397_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11871_ (.A1(_06352_),
    .A2(_06396_),
    .A3(_06397_),
    .Z(_06398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11872_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A2(_06398_),
    .ZN(_06399_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _11873_ (.A1(_06255_),
    .A2(_06234_),
    .A3(_06394_),
    .A4(_06351_),
    .Z(_06400_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3514 (.I(net423),
    .Z(net3514));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11875_ (.I(net3526),
    .ZN(_06402_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk_i_regs (.I(clknet_6_48__leaf_clk_i_regs),
    .Z(clknet_leaf_8_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11877_ (.A1(_06322_),
    .A2(_06331_),
    .B(_06400_),
    .C(net3419),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3493 (.I(net3490),
    .Z(net3493));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11879_ (.A1(_06241_),
    .A2(_06344_),
    .B(_06346_),
    .ZN(_06406_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11880_ (.A1(_06224_),
    .A2(_06406_),
    .Z(_06407_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11881_ (.A1(net3474),
    .A2(_06210_),
    .A3(net3473),
    .A4(_06246_),
    .Z(_06408_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11882_ (.I(\id_stage_i.controller_i.instr_i[14] ),
    .ZN(_06409_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11883_ (.A1(_06210_),
    .A2(net3416),
    .B(net3474),
    .ZN(_06410_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11884_ (.A1(net357),
    .A2(_06198_),
    .A3(net390),
    .Z(_06411_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11885_ (.A1(_06408_),
    .A2(_06410_),
    .B(_06411_),
    .ZN(_06412_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11886_ (.A1(_06354_),
    .A2(_06412_),
    .Z(_06413_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11887_ (.A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_06407_),
    .A3(_06343_),
    .A4(_06413_),
    .Z(_06414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11888_ (.A1(net3488),
    .A2(net3495),
    .ZN(_06415_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3625 (.I(net3624),
    .Z(net3625));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3519 (.I(net3516),
    .Z(net3519));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11891_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S0(net3514),
    .S1(net3501),
    .Z(_06418_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11892_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .S0(net3514),
    .S1(net3501),
    .Z(_06419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11893_ (.I0(_06418_),
    .I1(_06419_),
    .S(net3452),
    .Z(_06420_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11894_ (.A1(_06415_),
    .A2(_06420_),
    .Z(_06421_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11895_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S0(net3518),
    .S1(net3512),
    .Z(_06422_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11896_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .S0(net3518),
    .S1(net3512),
    .Z(_06423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11897_ (.I0(_06422_),
    .I1(_06423_),
    .S(net3452),
    .Z(_06424_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11898_ (.A1(net3488),
    .A2(net3426),
    .A3(_06424_),
    .Z(_06425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11899_ (.A1(net3488),
    .A2(net3426),
    .ZN(_06426_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11900_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S0(net3514),
    .S1(net3501),
    .Z(_06427_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11901_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .S0(net3514),
    .S1(net3501),
    .Z(_06428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11902_ (.I0(_06427_),
    .I1(_06428_),
    .S(net3452),
    .Z(_06429_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11903_ (.A1(_06426_),
    .A2(_06429_),
    .Z(_06430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11904_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S(net3518),
    .Z(_06431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11905_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .S(net3518),
    .Z(_06432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11906_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(net3518),
    .Z(_06433_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11907_ (.A1(net3518),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .Z(_06434_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11908_ (.I0(_06431_),
    .I1(_06432_),
    .I2(_06433_),
    .I3(_06434_),
    .S0(net3452),
    .S1(net3442),
    .Z(_06435_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11909_ (.A1(net3488),
    .A2(net3495),
    .A3(_06435_),
    .Z(_06436_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11910_ (.A1(_06436_),
    .A2(_06425_),
    .A3(_06430_),
    .A4(_06421_),
    .Z(_06437_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11911_ (.A1(_06355_),
    .A2(_06437_),
    .Z(_06438_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11912_ (.A1(_06404_),
    .A2(_06438_),
    .A3(_06414_),
    .ZN(_06439_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11913_ (.A1(_06399_),
    .A2(_06439_),
    .Z(_11391_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _11914_ (.I(_11391_[0]),
    .ZN(_06440_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3464 (.I(net3463),
    .Z(net3464));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11916_ (.A1(_06354_),
    .A2(_06351_),
    .ZN(_06441_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3454 (.I(_06284_),
    .Z(net3454));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11918_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S0(net3567),
    .S1(net3548),
    .Z(_06443_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11919_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .S0(net3575),
    .S1(net3548),
    .Z(_06444_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11920_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S0(net3567),
    .S1(net3548),
    .Z(_06445_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11921_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S0(net3567),
    .S1(net3548),
    .Z(_06446_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11922_ (.I0(_06443_),
    .I1(_06444_),
    .I2(_06445_),
    .I3(_06446_),
    .S0(net3436),
    .S1(net3425),
    .Z(_06447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11923_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .S(net3548),
    .Z(_06448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11924_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S(net3548),
    .Z(_06449_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11925_ (.A1(net3548),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .Z(_06450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11926_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(net3548),
    .Z(_06451_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11927_ (.I0(_06448_),
    .I1(_06449_),
    .I2(_06450_),
    .I3(_06451_),
    .S0(net3575),
    .S1(net3436),
    .Z(_06452_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11928_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S0(net3548),
    .S1(net3510),
    .Z(_06453_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11929_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .S0(net3548),
    .S1(net3510),
    .Z(_06454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11930_ (.I0(_06453_),
    .I1(_06454_),
    .S(net3445),
    .Z(_06455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11931_ (.I0(_06452_),
    .I1(_06455_),
    .S(net3494),
    .Z(_06456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _11932_ (.I0(_06447_),
    .I1(_06456_),
    .S(net3423),
    .Z(_06457_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11933_ (.A1(_06441_),
    .A2(_06457_),
    .Z(_06458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11934_ (.A1(_06338_),
    .A2(_06342_),
    .ZN(_06459_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3430 (.I(net3427),
    .Z(net3430));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3431 (.I(net3430),
    .Z(net3431));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11937_ (.A1(_06322_),
    .A2(_06331_),
    .B(_06459_),
    .C(net3440),
    .ZN(_06462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11938_ (.A1(_06224_),
    .A2(_06406_),
    .ZN(_06463_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11939_ (.A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_06463_),
    .A3(_06459_),
    .B(_06413_),
    .ZN(_06464_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11940_ (.A1(_06224_),
    .A2(_06347_),
    .B(_06234_),
    .ZN(_06465_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11941_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .A2(_06465_),
    .A3(_06396_),
    .A4(_06397_),
    .Z(_06466_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11942_ (.A1(_06462_),
    .A2(_06464_),
    .A3(_06466_),
    .Z(_06467_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11943_ (.A1(_06458_),
    .A2(_06467_),
    .Z(_11410_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11944_ (.I(_11410_[0]),
    .ZN(_11414_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3429 (.I(net3427),
    .Z(net3429));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11946_ (.A1(_06322_),
    .A2(_06331_),
    .B(_06400_),
    .C(net3425),
    .ZN(_06469_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11947_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S0(net3546),
    .S1(net3510),
    .Z(_06470_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11948_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .S0(net3546),
    .S1(net3510),
    .Z(_06471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11949_ (.I0(_06470_),
    .I1(_06471_),
    .S(net3453),
    .Z(_06472_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11950_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S0(net3567),
    .S1(net528),
    .Z(_06473_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11951_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .S0(net3567),
    .S1(net528),
    .Z(_06474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11952_ (.I0(_06473_),
    .I1(_06474_),
    .S(net3427),
    .Z(_06475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11953_ (.I0(_06472_),
    .I1(_06475_),
    .S(net3425),
    .Z(_06476_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11954_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S0(net528),
    .S1(net3510),
    .Z(_06477_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11955_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .S0(net3546),
    .S1(net3510),
    .Z(_06478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11956_ (.I0(_06477_),
    .I1(_06478_),
    .S(net3453),
    .Z(_06479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11957_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .S(net3546),
    .Z(_06480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11958_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S(net3546),
    .Z(_06481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11959_ (.A1(net528),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .Z(_06482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11960_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net3546),
    .Z(_06483_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3423 (.I(net3421),
    .Z(net3423));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11962_ (.I0(_06480_),
    .I1(_06481_),
    .I2(_06482_),
    .I3(_06483_),
    .S0(net3568),
    .S1(net3427),
    .Z(_06485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11963_ (.I0(_06479_),
    .I1(_06485_),
    .S(net3425),
    .Z(_06486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _11964_ (.I0(_06476_),
    .I1(_06486_),
    .S(net3423),
    .Z(_06487_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11965_ (.A1(_06355_),
    .A2(_06487_),
    .Z(_06488_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _11966_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .A2(_06352_),
    .A3(_06396_),
    .A4(_06397_),
    .Z(_06489_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _11967_ (.A1(_06469_),
    .A2(_06488_),
    .A3(_06489_),
    .ZN(_11422_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11968_ (.I(_11422_[0]),
    .ZN(_11418_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11969_ (.A1(_06382_),
    .A2(_06369_),
    .Z(_06490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11970_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .S(net575),
    .Z(_06491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11971_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S(net575),
    .Z(_06492_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11972_ (.A1(net3540),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .Z(_06493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11973_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net3540),
    .Z(_06494_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11974_ (.I0(_06491_),
    .I1(_06492_),
    .I2(_06493_),
    .I3(_06494_),
    .S0(net3566),
    .S1(net3433),
    .Z(_06495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11975_ (.A1(_06490_),
    .A2(_06495_),
    .ZN(_06496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11976_ (.A1(net3489),
    .A2(net3425),
    .Z(_06497_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11977_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S0(net3563),
    .S1(net3540),
    .Z(_06498_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11978_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S0(net3562),
    .S1(net3540),
    .Z(_06499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11979_ (.I0(_06498_),
    .I1(_06499_),
    .S(net3430),
    .Z(_06500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11980_ (.A1(_06497_),
    .A2(_06500_),
    .ZN(_06501_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3418 (.I(_06402_),
    .Z(net3418));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11982_ (.A1(net3554),
    .A2(net3526),
    .ZN(_06503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11983_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S(net3510),
    .Z(_06504_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11984_ (.A1(net3415),
    .A2(_06504_),
    .ZN(_06505_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3422 (.I(net3421),
    .Z(net3422));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11986_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .S(net3510),
    .Z(_06507_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _11987_ (.A1(net3448),
    .A2(net3527),
    .A3(_06507_),
    .ZN(_06508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11988_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .S(net3510),
    .Z(_06509_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _11989_ (.A1(net3562),
    .A2(net3420),
    .A3(_06509_),
    .ZN(_06510_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11990_ (.A1(net314),
    .A2(net3558),
    .Z(_06511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11991_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .S(net3510),
    .Z(_06512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11992_ (.A1(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .A2(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(_06513_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11993_ (.A1(net3411),
    .A2(_06512_),
    .B(net3410),
    .ZN(_06514_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _11994_ (.A1(_06505_),
    .A2(_06508_),
    .A3(_06510_),
    .A4(_06514_),
    .Z(_06515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11995_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S(net3510),
    .Z(_06516_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11996_ (.A1(net3415),
    .A2(_06516_),
    .ZN(_06517_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3412 (.I(net3411),
    .Z(net3412));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11998_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .S(net3510),
    .Z(_06519_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _11999_ (.A1(net3448),
    .A2(net3540),
    .A3(_06519_),
    .ZN(_06520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12000_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .S(net3510),
    .Z(_06521_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12001_ (.A1(net3562),
    .A2(net3420),
    .A3(_06521_),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12002_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .S(net3510),
    .Z(_06523_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12003_ (.A1(net3411),
    .A2(_06523_),
    .B(net3421),
    .C(net3491),
    .ZN(_06524_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12004_ (.A1(_06517_),
    .A2(_06520_),
    .A3(_06522_),
    .A4(_06524_),
    .Z(_06525_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12005_ (.A1(_06515_),
    .A2(_06501_),
    .A3(_06496_),
    .A4(_06525_),
    .ZN(_06526_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12006_ (.A1(_06355_),
    .A2(_06526_),
    .Z(_06527_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12007_ (.A1(_06322_),
    .A2(_06331_),
    .B(_06400_),
    .C(net3421),
    .ZN(_06528_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12008_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A2(_06352_),
    .A3(_06396_),
    .A4(_06397_),
    .Z(_06529_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _12009_ (.A1(_06527_),
    .A2(_06528_),
    .A3(_06529_),
    .ZN(_11430_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _12010_ (.I(_11430_[0]),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3415 (.I(net3414),
    .Z(net3415));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3420 (.I(net3418),
    .Z(net3420));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3419 (.I(net3418),
    .Z(net3419));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12014_ (.A1(_06224_),
    .A2(_06406_),
    .B(_06394_),
    .ZN(_06533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12015_ (.A1(_06441_),
    .A2(_06533_),
    .Z(_06534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12016_ (.A1(net3486),
    .A2(_06534_),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3426 (.I(_06369_),
    .Z(net3426));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3411 (.I(_06511_),
    .Z(net3411));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12019_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .S(net3526),
    .Z(_06538_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12020_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S(net3526),
    .Z(_06539_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3463 (.I(_06284_),
    .Z(net3463));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12022_ (.A1(net3526),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .Z(_06541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12023_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(net3526),
    .Z(_06542_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3404 (.I(_08646_),
    .Z(net3404));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3407 (.I(_08481_),
    .Z(net3407));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12026_ (.I0(_06538_),
    .I1(_06539_),
    .I2(_06541_),
    .I3(_06542_),
    .S0(net3556),
    .S1(net3443),
    .Z(_06545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12027_ (.A1(_06490_),
    .A2(_06545_),
    .ZN(_06546_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12028_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S0(net3556),
    .S1(net3526),
    .Z(_06547_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12029_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S0(net3556),
    .S1(net3526),
    .Z(_06548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12030_ (.I0(_06547_),
    .I1(_06548_),
    .S(net3443),
    .Z(_06549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12031_ (.A1(_06497_),
    .A2(_06549_),
    .ZN(_06550_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3408 (.I(_06735_),
    .Z(net3408));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3462 (.I(_06284_),
    .Z(net3462));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3413 (.I(net483),
    .Z(net3413));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12035_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S(net3510),
    .Z(_06554_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12036_ (.A1(net3415),
    .A2(_06554_),
    .ZN(_06555_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3397 (.I(_06717_),
    .Z(net3397));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12039_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .S(net3510),
    .Z(_06558_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12040_ (.A1(net3451),
    .A2(net3527),
    .A3(_06558_),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3396 (.I(_06933_),
    .Z(net3396));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12042_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .S(net3510),
    .Z(_06561_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12043_ (.A1(net3553),
    .A2(net3418),
    .A3(_06561_),
    .ZN(_06562_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3395 (.I(_05680_),
    .Z(net3395));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12045_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .S(net3510),
    .Z(_06564_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12046_ (.A1(net3411),
    .A2(_06564_),
    .B(net3410),
    .ZN(_06565_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12047_ (.A1(_06555_),
    .A2(_06559_),
    .A3(_06562_),
    .A4(_06565_),
    .Z(_06566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12048_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S(net3510),
    .Z(_06567_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12049_ (.A1(net3414),
    .A2(_06567_),
    .ZN(_06568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12050_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .S(net3510),
    .Z(_06569_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12051_ (.A1(net3451),
    .A2(net3527),
    .A3(_06569_),
    .ZN(_06570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12052_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .S(net3510),
    .Z(_06571_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12053_ (.A1(net3556),
    .A2(net3418),
    .A3(_06571_),
    .ZN(_06572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12054_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .S(net3510),
    .Z(_06573_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3394 (.I(_06234_),
    .Z(net3394));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12056_ (.A1(net3411),
    .A2(_06573_),
    .B(net3421),
    .C(net3490),
    .ZN(_06575_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12057_ (.A1(_06568_),
    .A2(_06570_),
    .A3(_06572_),
    .A4(_06575_),
    .Z(_06576_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12058_ (.A1(_06566_),
    .A2(_06550_),
    .A3(_06546_),
    .A4(_06576_),
    .ZN(_06577_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3393 (.I(_06586_),
    .Z(net3393));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12060_ (.A1(_06355_),
    .A2(net341),
    .ZN(_06579_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12061_ (.A1(_06535_),
    .A2(_06579_),
    .Z(_11438_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12062_ (.I(_11438_[0]),
    .ZN(_11434_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12063_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .S(net3527),
    .Z(_06580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12064_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S(net3527),
    .Z(_06581_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12065_ (.A1(net3527),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .Z(_06582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12066_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net3527),
    .Z(_06583_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12068_ (.I0(_06580_),
    .I1(_06581_),
    .I2(_06582_),
    .I3(_06583_),
    .S0(net3559),
    .S1(net3427),
    .Z(_06585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12069_ (.A1(net3399),
    .A2(_06585_),
    .ZN(_06586_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12070_ (.A1(net3554),
    .A2(_06513_),
    .Z(_06587_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3460 (.I(net3454),
    .Z(net3460));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3392 (.I(_06594_),
    .Z(net3392));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12073_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S0(net3532),
    .S1(net3504),
    .Z(_06590_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12074_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .S0(net3532),
    .S1(net3504),
    .Z(_06591_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3391 (.I(_06605_),
    .Z(net3391));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12076_ (.A1(net3450),
    .A2(_06513_),
    .Z(_06593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12077_ (.A1(_06587_),
    .A2(_06590_),
    .B1(_06591_),
    .B2(net3398),
    .ZN(_06594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12078_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S(net3506),
    .Z(_06595_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12079_ (.A1(net3414),
    .A2(_06595_),
    .ZN(_06596_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3390 (.I(_06614_),
    .Z(net3390));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12081_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .S(net3506),
    .Z(_06598_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12082_ (.A1(net3449),
    .A2(net3532),
    .A3(_06598_),
    .ZN(_06599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12083_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .S(net3506),
    .Z(_06600_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12084_ (.A1(net3559),
    .A2(net3419),
    .A3(_06600_),
    .ZN(_06601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12085_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .S(net3506),
    .Z(_06602_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3389 (.I(_06804_),
    .Z(net3389));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12087_ (.A1(net3412),
    .A2(_06602_),
    .B(net3489),
    .C(net3425),
    .ZN(_06604_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12088_ (.A1(_06596_),
    .A2(_06599_),
    .A3(_06601_),
    .A4(_06604_),
    .Z(_06605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12089_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S(net3505),
    .Z(_06606_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12090_ (.A1(net3414),
    .A2(_06606_),
    .ZN(_06607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12091_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .S(net3507),
    .Z(_06608_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12092_ (.A1(net3449),
    .A2(net3532),
    .A3(_06608_),
    .ZN(_06609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12093_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .S(net3505),
    .Z(_06610_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12094_ (.A1(net3559),
    .A2(net3419),
    .A3(_06610_),
    .ZN(_06611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12095_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .S(net3507),
    .Z(_06612_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12096_ (.A1(net3412),
    .A2(_06612_),
    .B(net3421),
    .C(net3490),
    .ZN(_06613_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12097_ (.A1(_06607_),
    .A2(_06609_),
    .A3(_06611_),
    .A4(_06613_),
    .Z(_06614_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12098_ (.A1(net3393),
    .A2(net3392),
    .A3(net3391),
    .A4(net3390),
    .Z(_06615_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3388 (.I(_06817_),
    .Z(net3388));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12100_ (.A1(net3485),
    .A2(_06533_),
    .ZN(_06617_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3387 (.I(_06821_),
    .Z(net3387));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12102_ (.I0(_06615_),
    .I1(_06617_),
    .S(_06441_),
    .Z(_11446_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12103_ (.I(_11446_[0]),
    .ZN(_11442_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3386 (.I(_06831_),
    .Z(net3386));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12105_ (.I(net3484),
    .ZN(_06620_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12106_ (.A1(_06323_),
    .A2(_06325_),
    .B1(_06412_),
    .B2(_06234_),
    .C(_06342_),
    .ZN(_06621_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12107_ (.A1(_06620_),
    .A2(_06621_),
    .ZN(_06622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12108_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .S(net3526),
    .Z(_06623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12109_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S(net3526),
    .Z(_06624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12110_ (.A1(net3526),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .Z(_06625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12111_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net3526),
    .Z(_06626_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12112_ (.I0(_06623_),
    .I1(_06624_),
    .I2(_06625_),
    .I3(_06626_),
    .S0(net3555),
    .S1(net3441),
    .Z(_06627_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12113_ (.A1(net3399),
    .A2(_06627_),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12114_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S0(net3531),
    .S1(net3504),
    .Z(_06629_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12115_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .S0(net3531),
    .S1(net3504),
    .Z(_06630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12116_ (.A1(_06587_),
    .A2(_06629_),
    .B1(_06630_),
    .B2(net3398),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3406 (.I(_08644_),
    .Z(net3406));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12118_ (.A1(net3559),
    .A2(net3505),
    .Z(_06633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12119_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .S(net3531),
    .Z(_06634_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12120_ (.A1(_06633_),
    .A2(_06634_),
    .ZN(_06635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12121_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S(net3531),
    .Z(_06636_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12122_ (.A1(net3450),
    .A2(net3510),
    .A3(_06636_),
    .ZN(_06637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12123_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .S(net3531),
    .Z(_06638_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12124_ (.A1(net3554),
    .A2(net3441),
    .A3(_06638_),
    .ZN(_06639_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12125_ (.A1(net3554),
    .A2(net3511),
    .ZN(_06640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12126_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S(net3531),
    .Z(_06641_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12127_ (.A1(_06640_),
    .A2(_06641_),
    .B(net3488),
    .C(net3425),
    .ZN(_06642_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12128_ (.A1(_06635_),
    .A2(_06637_),
    .A3(_06639_),
    .A4(_06642_),
    .Z(_06643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12129_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S(net3510),
    .Z(_06644_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12130_ (.A1(net3414),
    .A2(_06644_),
    .ZN(_06645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12131_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .S(net3510),
    .Z(_06646_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12132_ (.A1(net3451),
    .A2(net3527),
    .A3(_06646_),
    .ZN(_06647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12133_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .S(net3510),
    .Z(_06648_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12134_ (.A1(net3554),
    .A2(net3418),
    .A3(_06648_),
    .ZN(_06649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12135_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .S(net3510),
    .Z(_06650_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12136_ (.A1(net3411),
    .A2(_06650_),
    .B(net3421),
    .C(net3490),
    .ZN(_06651_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12137_ (.A1(_06645_),
    .A2(_06647_),
    .A3(_06649_),
    .A4(_06651_),
    .Z(_06652_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12138_ (.A1(_06643_),
    .A2(_06631_),
    .A3(_06628_),
    .A4(_06652_),
    .ZN(_06653_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12139_ (.A1(_06355_),
    .A2(_06653_),
    .Z(_06654_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _12140_ (.A1(_06622_),
    .A2(_06654_),
    .ZN(_11454_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12141_ (.I(_11454_[0]),
    .ZN(_11450_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12142_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .S(net3516),
    .Z(_06655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12143_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S(net3516),
    .Z(_06656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12144_ (.A1(net3516),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .Z(_06657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12145_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net3516),
    .Z(_06658_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12146_ (.I0(_06655_),
    .I1(_06656_),
    .I2(_06657_),
    .I3(_06658_),
    .S0(net3556),
    .S1(_06367_),
    .Z(_06659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12147_ (.A1(_06490_),
    .A2(_06659_),
    .ZN(_06660_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3384 (.I(_06926_),
    .Z(net3384));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12149_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S0(net3514),
    .S1(net3501),
    .Z(_06662_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12150_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .S0(net3514),
    .S1(net3501),
    .Z(_06663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12151_ (.A1(_06587_),
    .A2(_06662_),
    .B1(_06663_),
    .B2(_06593_),
    .ZN(_06664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12152_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S(net3500),
    .Z(_06665_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12153_ (.A1(_06503_),
    .A2(_06665_),
    .ZN(_06666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12154_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .S(net3500),
    .Z(_06667_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12155_ (.A1(net3450),
    .A2(net3517),
    .A3(_06667_),
    .ZN(_06668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12156_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .S(net3500),
    .Z(_06669_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12157_ (.A1(net3556),
    .A2(_06402_),
    .A3(_06669_),
    .ZN(_06670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12158_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .S(net3500),
    .Z(_06671_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12159_ (.A1(net483),
    .A2(_06671_),
    .B(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .C(_06369_),
    .ZN(_06672_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12160_ (.A1(_06666_),
    .A2(_06668_),
    .A3(_06670_),
    .A4(_06672_),
    .Z(_06673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12161_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S(net3509),
    .Z(_06674_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12162_ (.A1(_06503_),
    .A2(_06674_),
    .ZN(_06675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12163_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .S(net3509),
    .Z(_06676_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12164_ (.A1(net3450),
    .A2(net558),
    .A3(_06676_),
    .ZN(_06677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12165_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .S(net3509),
    .Z(_06678_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12166_ (.A1(net3556),
    .A2(_06402_),
    .A3(_06678_),
    .ZN(_06679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12167_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .S(net3509),
    .Z(_06680_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12168_ (.A1(_06511_),
    .A2(_06680_),
    .B(_06382_),
    .C(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .ZN(_06681_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12169_ (.A1(_06675_),
    .A2(_06677_),
    .A3(_06679_),
    .A4(_06681_),
    .Z(_06682_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12170_ (.A1(_06673_),
    .A2(_06664_),
    .A3(_06660_),
    .A4(_06682_),
    .ZN(_06683_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3383 (.I(net300),
    .Z(net3383));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3382 (.I(_08653_),
    .Z(net3382));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12173_ (.A1(net3483),
    .A2(_06441_),
    .A3(_06533_),
    .Z(_06686_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12174_ (.A1(_06355_),
    .A2(net412),
    .B(_06686_),
    .ZN(_11462_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12175_ (.I(_11462_[0]),
    .ZN(_11458_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12176_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .S(net3520),
    .Z(_06687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12177_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S(net3520),
    .Z(_06688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12178_ (.A1(net558),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .Z(_06689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12179_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(net3520),
    .Z(_06690_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12180_ (.I0(_06687_),
    .I1(_06688_),
    .I2(_06689_),
    .I3(_06690_),
    .S0(net3556),
    .S1(_06367_),
    .Z(_06691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12181_ (.A1(_06490_),
    .A2(_06691_),
    .ZN(_06692_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12182_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S0(net3514),
    .S1(net3501),
    .Z(_06693_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12183_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .S0(net3514),
    .S1(net3501),
    .Z(_06694_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12184_ (.A1(_06587_),
    .A2(_06693_),
    .B1(_06694_),
    .B2(_06593_),
    .ZN(_06695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12185_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S(net3502),
    .Z(_06696_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12186_ (.A1(_06503_),
    .A2(_06696_),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12187_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .S(net3502),
    .Z(_06698_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12188_ (.A1(net3450),
    .A2(net3517),
    .A3(_06698_),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12189_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .S(net3500),
    .Z(_06700_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12190_ (.A1(net3556),
    .A2(_06402_),
    .A3(_06700_),
    .ZN(_06701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12191_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .S(net3502),
    .Z(_06702_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12192_ (.A1(net3413),
    .A2(_06702_),
    .B(net3488),
    .C(_06369_),
    .ZN(_06703_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12193_ (.A1(_06697_),
    .A2(_06699_),
    .A3(_06701_),
    .A4(_06703_),
    .Z(_06704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12194_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S(net3512),
    .Z(_06705_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12195_ (.A1(_06503_),
    .A2(_06705_),
    .ZN(_06706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12196_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .S(net3512),
    .Z(_06707_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12197_ (.A1(net3450),
    .A2(net559),
    .A3(_06707_),
    .ZN(_06708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12198_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .S(net3512),
    .Z(_06709_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12199_ (.A1(net3556),
    .A2(_06402_),
    .A3(_06709_),
    .ZN(_06710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12200_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .S(net3512),
    .Z(_06711_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12201_ (.A1(net483),
    .A2(_06711_),
    .B(_06382_),
    .C(net3490),
    .ZN(_06712_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12202_ (.A1(_06706_),
    .A2(_06708_),
    .A3(_06710_),
    .A4(_06712_),
    .Z(_06713_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12203_ (.A1(_06704_),
    .A2(_06695_),
    .A3(_06692_),
    .A4(_06713_),
    .ZN(_06714_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3381 (.I(_06309_),
    .Z(net3381));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12205_ (.A1(net3482),
    .A2(_06441_),
    .A3(_06533_),
    .Z(_06716_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12206_ (.A1(_06355_),
    .A2(net407),
    .B(_06716_),
    .ZN(_11470_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12207_ (.I(_11470_[0]),
    .ZN(_11466_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12208_ (.A1(_06242_),
    .A2(_06243_),
    .ZN(_06717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12209_ (.A1(_06206_),
    .A2(net3397),
    .Z(_06718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12210_ (.A1(net3482),
    .A2(net3483),
    .ZN(_06719_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _12211_ (.A1(net3497),
    .A2(net3419),
    .A3(net3409),
    .A4(_06719_),
    .ZN(_06720_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3380 (.I(_06355_),
    .Z(net3380));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12213_ (.A1(net3484),
    .A2(net3485),
    .A3(net3479),
    .Z(_06722_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3379 (.I(_06413_),
    .Z(net3379));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12215_ (.A1(net3487),
    .A2(\id_stage_i.controller_i.instr_i[25] ),
    .A3(\id_stage_i.controller_i.instr_i[30] ),
    .Z(_06724_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12216_ (.A1(net3498),
    .A2(net3552),
    .A3(net3482),
    .Z(_06725_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12217_ (.A1(_06722_),
    .A2(_06724_),
    .A3(_06725_),
    .ZN(_06726_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12218_ (.A1(net3499),
    .A2(net3483),
    .ZN(_06727_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12219_ (.A1(net3560),
    .A2(net3499),
    .A3(net3483),
    .Z(_06728_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12220_ (.A1(_06727_),
    .A2(_06728_),
    .Z(_06729_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12221_ (.A1(_06726_),
    .A2(_06729_),
    .Z(_06730_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _12222_ (.A1(net3487),
    .A2(\id_stage_i.controller_i.instr_i[25] ),
    .A3(net3484),
    .A4(\id_stage_i.controller_i.instr_i[30] ),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12223_ (.A1(net3487),
    .A2(\id_stage_i.controller_i.instr_i[25] ),
    .A3(net3484),
    .A4(\id_stage_i.controller_i.instr_i[30] ),
    .Z(_06732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12224_ (.A1(_06731_),
    .A2(_06732_),
    .B(net3485),
    .C(net3479),
    .ZN(_06733_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3378 (.I(net448),
    .Z(net3378));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12226_ (.A1(net3576),
    .A2(net3578),
    .A3(net3581),
    .A4(net3596),
    .Z(_06735_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12227_ (.A1(net3607),
    .A2(net3408),
    .ZN(_06736_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _12228_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .ZN(_06737_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3377 (.I(_06880_),
    .Z(net3377));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12230_ (.I(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .ZN(_06739_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _12231_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12232_ (.A1(net3416),
    .A2(_06739_),
    .A3(_06740_),
    .Z(_06741_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12233_ (.A1(_06733_),
    .A2(_06736_),
    .A3(_06737_),
    .A4(_06741_),
    .Z(_06742_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _12234_ (.A1(_06720_),
    .A2(_06730_),
    .B(_06742_),
    .C(_06206_),
    .ZN(_06743_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _12235_ (.I(net304),
    .ZN(_06744_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3376 (.I(_06916_),
    .Z(net3376));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12237_ (.A1(_06744_),
    .A2(_06242_),
    .ZN(_06746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12238_ (.A1(net3478),
    .A2(_06220_),
    .B(net3474),
    .ZN(_06747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12239_ (.I0(net3481),
    .I1(net3474),
    .S(net3477),
    .Z(_06748_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _12240_ (.A1(_06747_),
    .A2(net3477),
    .A3(_06391_),
    .B1(_06748_),
    .B2(net3478),
    .ZN(_06749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12241_ (.A1(net3474),
    .A2(_06220_),
    .B(_06392_),
    .ZN(_06750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _12242_ (.A1(_06206_),
    .A2(_06746_),
    .B1(net328),
    .B2(_06750_),
    .ZN(_06751_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12243_ (.A1(_06222_),
    .A2(net3469),
    .ZN(_06752_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12244_ (.A1(net3649),
    .A2(net3646),
    .Z(_06753_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12245_ (.A1(net3648),
    .A2(net3416),
    .B1(_06753_),
    .B2(net3481),
    .ZN(_06754_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3374 (.I(_07012_),
    .Z(net3374));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12247_ (.A1(net3475),
    .A2(net3646),
    .B1(_06753_),
    .B2(net3648),
    .ZN(_06756_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12248_ (.A1(\id_stage_i.controller_i.instr_i[6] ),
    .A2(\id_stage_i.controller_i.instr_i[4] ),
    .ZN(_06757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _12249_ (.A1(net3469),
    .A2(_06202_),
    .A3(_06757_),
    .ZN(_06758_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _12250_ (.A1(_06245_),
    .A2(_06752_),
    .A3(_06754_),
    .B1(_06756_),
    .B2(_06758_),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3405 (.I(_08645_),
    .Z(net3405));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12252_ (.A1(_06744_),
    .A2(net3649),
    .Z(_06761_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _12253_ (.I(\id_stage_i.controller_i.instr_i[30] ),
    .ZN(_06762_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _12254_ (.A1(\id_stage_i.controller_i.instr_i[29] ),
    .A2(\id_stage_i.controller_i.instr_i[28] ),
    .A3(\id_stage_i.controller_i.instr_i[31] ),
    .ZN(_06763_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12255_ (.A1(\id_stage_i.controller_i.instr_i[25] ),
    .A2(\id_stage_i.controller_i.instr_i[27] ),
    .A3(\id_stage_i.controller_i.instr_i[26] ),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12256_ (.A1(net3646),
    .A2(_06762_),
    .B(_06763_),
    .C(_06764_),
    .ZN(_06765_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12257_ (.A1(net3477),
    .A2(net269),
    .A3(net265),
    .A4(_06212_),
    .Z(_06766_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12258_ (.A1(_06761_),
    .A2(_06765_),
    .A3(_06766_),
    .Z(_06767_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12259_ (.A1(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .A2(_06228_),
    .A3(_06759_),
    .A4(_06767_),
    .Z(_06768_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12260_ (.A1(\id_stage_i.controller_i.instr_i[27] ),
    .A2(\id_stage_i.controller_i.instr_i[26] ),
    .ZN(_06769_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12261_ (.A1(net3486),
    .A2(net3480),
    .ZN(_06770_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12262_ (.A1(\id_stage_i.controller_i.instr_i[13] ),
    .A2(_06763_),
    .A3(_06769_),
    .A4(_06770_),
    .Z(_06771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12263_ (.A1(net320),
    .A2(_06771_),
    .ZN(_06772_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12264_ (.I(net3486),
    .ZN(_06773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12265_ (.A1(net3649),
    .A2(_06773_),
    .B(net3480),
    .ZN(_06774_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12266_ (.A1(net3649),
    .A2(net3646),
    .ZN(_06775_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12267_ (.A1(_06773_),
    .A2(_06775_),
    .Z(_06776_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12268_ (.A1(_06763_),
    .A2(_06769_),
    .Z(_06777_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12269_ (.A1(_06744_),
    .A2(_06774_),
    .B1(_06776_),
    .B2(_06762_),
    .C(_06777_),
    .ZN(_06778_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12270_ (.A1(_06319_),
    .A2(\id_stage_i.controller_i.instr_i[4] ),
    .Z(_06779_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12271_ (.A1(_06411_),
    .A2(_06779_),
    .Z(_06780_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12272_ (.A1(_06772_),
    .A2(_06778_),
    .A3(net324),
    .Z(_06781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _12273_ (.A1(_06743_),
    .A2(_06751_),
    .B(_06768_),
    .C(_06781_),
    .ZN(_06782_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12274_ (.A1(_06718_),
    .A2(_06782_),
    .Z(_06783_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3375 (.I(net3374),
    .Z(net3375));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12276_ (.A1(_11466_[0]),
    .A2(_06783_),
    .Z(_11157_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12277_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S0(net3525),
    .S1(net3511),
    .Z(_06785_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12278_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .S0(net3525),
    .S1(net3511),
    .Z(_06786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12279_ (.I0(_06785_),
    .I1(_06786_),
    .S(net3450),
    .Z(_06787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12280_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .S(net3525),
    .Z(_06788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12281_ (.A1(net3555),
    .A2(_06788_),
    .ZN(_06789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12282_ (.A1(net3525),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .Z(_06790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12283_ (.A1(net3451),
    .A2(_06790_),
    .B(net3511),
    .ZN(_06791_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12284_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .S(net3525),
    .Z(_06792_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12285_ (.A1(net3555),
    .A2(net3441),
    .A3(_06792_),
    .ZN(_06793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12286_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S(net3525),
    .Z(_06794_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12287_ (.A1(_06640_),
    .A2(_06794_),
    .B(net3425),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12288_ (.A1(_06789_),
    .A2(_06791_),
    .B(_06793_),
    .C(_06795_),
    .ZN(_06796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12289_ (.A1(net3495),
    .A2(_06787_),
    .B(net3488),
    .C(_06796_),
    .ZN(_06797_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12290_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S0(net3554),
    .S1(net3514),
    .Z(_06798_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12291_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .S0(net3554),
    .S1(net314),
    .Z(_06799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12292_ (.I0(_06798_),
    .I1(_06799_),
    .S(net3441),
    .Z(_06800_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12293_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S0(net3515),
    .S1(net3511),
    .Z(_06801_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12294_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .S0(net3515),
    .S1(net3511),
    .Z(_06802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12295_ (.I0(_06801_),
    .I1(_06802_),
    .S(net3450),
    .Z(_06803_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _12296_ (.A1(_06415_),
    .A2(_06800_),
    .B1(_06803_),
    .B2(_06426_),
    .ZN(_06804_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _12297_ (.A1(_06804_),
    .A2(_06797_),
    .ZN(_06805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _12298_ (.A1(net3480),
    .A2(_06534_),
    .B1(_06805_),
    .B2(_06355_),
    .ZN(_11478_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12299_ (.I(_11478_[0]),
    .ZN(_11474_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12300_ (.A1(_06322_),
    .A2(_06331_),
    .Z(_06806_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12301_ (.A1(net3449),
    .A2(_06255_),
    .A3(_06394_),
    .Z(_06807_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12302_ (.A1(_06255_),
    .A2(_06394_),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .ZN(_06808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12303_ (.I0(_06807_),
    .I1(_06808_),
    .S(_06465_),
    .Z(_06809_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12304_ (.A1(net3479),
    .A2(_06343_),
    .A3(_06465_),
    .ZN(_06810_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _12305_ (.A1(_06806_),
    .A2(_06809_),
    .B(_06810_),
    .C(_06441_),
    .ZN(_06811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12306_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .S(net3533),
    .Z(_06812_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12307_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S(net3533),
    .Z(_06813_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12308_ (.A1(net3533),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .Z(_06814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12309_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(net3533),
    .Z(_06815_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12310_ (.I0(_06812_),
    .I1(_06813_),
    .I2(_06814_),
    .I3(_06815_),
    .S0(net3561),
    .S1(net3427),
    .Z(_06816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12311_ (.A1(_06490_),
    .A2(_06816_),
    .ZN(_06817_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12312_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S0(net3561),
    .S1(net3533),
    .Z(_06818_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12313_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .S0(net3561),
    .S1(net3533),
    .Z(_06819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12314_ (.I0(_06818_),
    .I1(_06819_),
    .S(net3427),
    .Z(_06820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12315_ (.A1(net3410),
    .A2(_06820_),
    .ZN(_06821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12316_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .S(net3531),
    .Z(_06822_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12317_ (.A1(_06633_),
    .A2(_06822_),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12318_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S(net3531),
    .Z(_06824_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12319_ (.A1(net3448),
    .A2(net3507),
    .A3(_06824_),
    .ZN(_06825_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3370 (.I(_07066_),
    .Z(net3370));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12321_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .S(net3531),
    .Z(_06827_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12322_ (.A1(net3559),
    .A2(net3440),
    .A3(_06827_),
    .ZN(_06828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12323_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S(net3531),
    .Z(_06829_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12324_ (.A1(_06640_),
    .A2(_06829_),
    .B(net3489),
    .C(net3425),
    .ZN(_06830_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12325_ (.A1(_06823_),
    .A2(_06825_),
    .A3(_06828_),
    .A4(_06830_),
    .Z(_06831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12326_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S(net3505),
    .Z(_06832_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12327_ (.A1(net3414),
    .A2(_06832_),
    .ZN(_06833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12328_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .S(net3505),
    .Z(_06834_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12329_ (.A1(net3448),
    .A2(net3532),
    .A3(_06834_),
    .ZN(_06835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12330_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .S(net3505),
    .Z(_06836_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12331_ (.A1(net3561),
    .A2(net3418),
    .A3(_06836_),
    .ZN(_06837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12332_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .S(net3505),
    .Z(_06838_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12333_ (.A1(net3411),
    .A2(_06838_),
    .B(net3421),
    .C(net3490),
    .ZN(_06839_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12334_ (.A1(_06833_),
    .A2(_06835_),
    .A3(_06837_),
    .A4(_06839_),
    .Z(_06840_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12335_ (.A1(net3388),
    .A2(net3387),
    .A3(net3386),
    .A4(net3385),
    .Z(_06841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12336_ (.A1(_06355_),
    .A2(_06841_),
    .Z(_06842_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12337_ (.I(_06842_),
    .ZN(_06843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12338_ (.A1(_06811_),
    .A2(_06843_),
    .ZN(_11486_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12339_ (.I(_11486_[0]),
    .ZN(_11482_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3369 (.I(_07087_),
    .Z(net3369));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12341_ (.A1(\id_stage_i.controller_i.instr_i[13] ),
    .A2(_06736_),
    .ZN(_06845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _12342_ (.A1(\id_stage_i.controller_i.instr_i[12] ),
    .A2(_06206_),
    .A3(_06845_),
    .ZN(_11147_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12343_ (.I(_11147_[0]),
    .ZN(_11150_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3368 (.I(_07105_),
    .Z(net3368));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3367 (.I(_07132_),
    .Z(net3367));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3366 (.I(net858),
    .Z(net3366));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _12347_ (.A1(net3607),
    .A2(net3408),
    .B(_06206_),
    .C(net303),
    .ZN(_06849_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3365 (.I(_07172_),
    .Z(net3365));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3364 (.I(_07220_),
    .Z(net3364));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12350_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[11] ),
    .ZN(_06851_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3363 (.I(net443),
    .Z(net3363));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12352_ (.A1(_06237_),
    .A2(_06851_),
    .B(_06257_),
    .ZN(_06853_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3362 (.I(_07278_),
    .Z(net3362));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3361 (.I(_07368_),
    .Z(net3361));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12355_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S0(net3633),
    .S1(net3591),
    .Z(_06856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12356_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(net3633),
    .Z(_06857_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3360 (.I(_07525_),
    .Z(net3360));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12358_ (.A1(net3633),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .Z(_06859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12359_ (.I0(_06857_),
    .I1(_06859_),
    .S(net3465),
    .Z(_06860_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3358 (.I(_07711_),
    .Z(net3358));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12361_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S0(net453),
    .S1(net3591),
    .Z(_06862_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12362_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .S0(net453),
    .S1(net3591),
    .Z(_06863_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3357 (.I(_08038_),
    .Z(net3357));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12364_ (.I0(_06856_),
    .I1(_06860_),
    .I2(_06862_),
    .I3(_06863_),
    .S0(net3458),
    .S1(net3578),
    .Z(_06865_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3353 (.I(_06237_),
    .Z(net3353));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3354 (.I(_08656_),
    .Z(net3354));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3352 (.I(_06257_),
    .Z(net3352));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3351 (.I(net470),
    .Z(net3351));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12369_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S0(net3615),
    .S1(net3591),
    .Z(_06870_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3350 (.I(_07470_),
    .Z(net3350));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12371_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S0(net3615),
    .S1(net3591),
    .Z(_06872_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3349 (.I(net445),
    .Z(net3349));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3348 (.I(_07659_),
    .Z(net3348));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12374_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S0(net3633),
    .S1(net3591),
    .Z(_06875_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3347 (.I(_07756_),
    .Z(net3347));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12376_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .S0(net3633),
    .S1(net3591),
    .Z(_06877_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12377_ (.I0(_06870_),
    .I1(_06872_),
    .I2(_06875_),
    .I3(_06877_),
    .S0(net3458),
    .S1(net3578),
    .Z(_06878_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12378_ (.A1(_06290_),
    .A2(_06878_),
    .Z(_06879_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12379_ (.A1(net3576),
    .A2(_06865_),
    .B(_06879_),
    .ZN(_06880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12380_ (.A1(_06310_),
    .A2(net3377),
    .ZN(_06881_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3346 (.I(net411),
    .Z(net3346));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12382_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(_06313_),
    .Z(_06883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12383_ (.A1(_06853_),
    .A2(_06881_),
    .A3(_06883_),
    .Z(_11481_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _12384_ (.I(_11481_[0]),
    .ZN(_11485_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12385_ (.A1(net3469),
    .A2(_06207_),
    .ZN(_06884_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12386_ (.A1(net3478),
    .A2(_06345_),
    .A3(net275),
    .Z(_06885_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12387_ (.A1(_06222_),
    .A2(net3477),
    .A3(net322),
    .Z(_06886_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12388_ (.A1(_06213_),
    .A2(_06717_),
    .B1(_06215_),
    .B2(_06885_),
    .C(_06886_),
    .ZN(_06887_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12389_ (.A1(net3478),
    .A2(net321),
    .A3(_06250_),
    .Z(_06888_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12390_ (.A1(_06319_),
    .A2(net3475),
    .B(_06391_),
    .ZN(_06889_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12391_ (.A1(_06245_),
    .A2(_06889_),
    .B(net3478),
    .ZN(_06890_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12392_ (.A1(_06323_),
    .A2(_06887_),
    .B1(_06888_),
    .B2(_06890_),
    .C(_06338_),
    .ZN(_06891_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12393_ (.A1(_06884_),
    .A2(_06891_),
    .B(_06354_),
    .ZN(_06892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12394_ (.A1(net3607),
    .A2(_06718_),
    .ZN(_06893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12395_ (.A1(_06208_),
    .A2(_06256_),
    .B(net3394),
    .C(_06893_),
    .ZN(_06894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _12396_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .A2(_06892_),
    .B(_06894_),
    .C(_06313_),
    .ZN(_06895_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3345 (.I(net469),
    .Z(net3345));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3344 (.I(net439),
    .Z(net3344));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3343 (.I(_07957_),
    .Z(net3343));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3359 (.I(_07624_),
    .Z(net3359));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12401_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S0(net3626),
    .S1(net3593),
    .Z(_06900_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12402_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .S0(net3626),
    .S1(net3593),
    .Z(_06901_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3342 (.I(_08001_),
    .Z(net3342));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3459 (.I(net3454),
    .Z(net3459));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12405_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S0(net3626),
    .S1(net3593),
    .Z(_06904_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12406_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .S0(net3626),
    .S1(net3593),
    .Z(_06905_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3458 (.I(net3454),
    .Z(net3458));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3402 (.I(_08650_),
    .Z(net3402));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12409_ (.I0(_06900_),
    .I1(_06901_),
    .I2(_06904_),
    .I3(_06905_),
    .S0(net3457),
    .S1(net3578),
    .Z(_06908_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12410_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S0(net3624),
    .S1(net3603),
    .Z(_06909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12411_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(net3624),
    .Z(_06910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12412_ (.A1(net3624),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .Z(_06911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12413_ (.I0(_06910_),
    .I1(_06911_),
    .S(net3466),
    .Z(_06912_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12414_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S0(net3625),
    .S1(net3593),
    .Z(_06913_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12415_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .S0(net3625),
    .S1(net3593),
    .Z(_06914_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12416_ (.I0(_06909_),
    .I1(_06912_),
    .I2(_06913_),
    .I3(_06914_),
    .S0(net3456),
    .S1(net3578),
    .Z(_06915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12417_ (.I0(_06908_),
    .I1(_06915_),
    .S(_06290_),
    .Z(_06916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12418_ (.A1(_06208_),
    .A2(_06236_),
    .ZN(_06917_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12419_ (.A1(_06892_),
    .A2(net3376),
    .B(_06917_),
    .ZN(_06918_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _12420_ (.A1(_06895_),
    .A2(_06918_),
    .ZN(_11395_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12421_ (.I(_11395_[0]),
    .ZN(_11399_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12422_ (.I(\cs_registers_i.pc_id_i[1] ),
    .ZN(_06919_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12423_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S0(net3613),
    .S1(net3583),
    .Z(_06920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12424_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(net416),
    .Z(_06921_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12425_ (.A1(net333),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .Z(_06922_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12426_ (.I0(_06921_),
    .I1(_06922_),
    .S(_06275_),
    .Z(_06923_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12427_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S0(net333),
    .S1(net3583),
    .Z(_06924_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12428_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .S0(net333),
    .S1(net3583),
    .Z(_06925_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12429_ (.I0(_06920_),
    .I1(_06923_),
    .I2(_06924_),
    .I3(_06925_),
    .S0(net3462),
    .S1(net3578),
    .Z(_06926_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3425 (.I(_06369_),
    .Z(net3425));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12431_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S0(net333),
    .S1(net3583),
    .Z(_06928_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12432_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .S0(net416),
    .S1(net3583),
    .Z(_06929_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3410 (.I(_06513_),
    .Z(net3410));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12434_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S0(net333),
    .S1(net3583),
    .Z(_06931_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12435_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .S0(net333),
    .S1(net3583),
    .Z(_06932_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12436_ (.I0(_06928_),
    .I1(_06929_),
    .I2(_06931_),
    .I3(_06932_),
    .S0(net3463),
    .S1(net3578),
    .Z(_06933_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12437_ (.A1(_06290_),
    .A2(net3396),
    .Z(_06934_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12438_ (.A1(net3576),
    .A2(net3384),
    .B(_06934_),
    .ZN(_06935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12439_ (.I0(_06919_),
    .I1(_06935_),
    .S(_06892_),
    .Z(_06936_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3341 (.I(_08094_),
    .Z(net3341));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12441_ (.A1(_06208_),
    .A2(_06256_),
    .B(net3394),
    .ZN(_06938_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3409 (.I(_06633_),
    .Z(net3409));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3356 (.I(_08215_),
    .Z(net3356));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3355 (.I(_08505_),
    .Z(net3355));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12445_ (.A1(net3605),
    .A2(_06718_),
    .Z(_06942_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12446_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A2(net3394),
    .B1(_06938_),
    .B2(_06942_),
    .ZN(_06943_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12447_ (.A1(_06917_),
    .A2(_06936_),
    .B(_06943_),
    .ZN(_11402_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12448_ (.I(_11402_[0]),
    .ZN(_11406_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3400 (.I(_03079_),
    .Z(net3400));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3398 (.I(_06593_),
    .Z(net3398));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12451_ (.A1(net3649),
    .A2(\id_stage_i.controller_i.instr_i[14] ),
    .A3(_06762_),
    .Z(_06946_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3372 (.I(_07060_),
    .Z(net3372));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3339 (.I(_08177_),
    .Z(net3339));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12454_ (.A1(_06242_),
    .A2(_06409_),
    .A3(\id_stage_i.controller_i.instr_i[30] ),
    .Z(_06949_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12455_ (.A1(_06946_),
    .A2(_06949_),
    .B(_06744_),
    .ZN(_06950_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12456_ (.A1(_06744_),
    .A2(net3649),
    .A3(net3480),
    .B(_06950_),
    .ZN(_06951_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12457_ (.A1(_06763_),
    .A2(_06764_),
    .A3(_06780_),
    .A4(_06951_),
    .Z(_06952_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12458_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(_06246_),
    .Z(_06953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12459_ (.A1(_06254_),
    .A2(_06953_),
    .Z(_06954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12460_ (.I0(_06766_),
    .I1(_06954_),
    .S(_06744_),
    .Z(_06955_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12461_ (.A1(_06242_),
    .A2(_06955_),
    .Z(_06956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12462_ (.A1(_06953_),
    .A2(_06254_),
    .ZN(_06957_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _12463_ (.A1(\id_stage_i.controller_i.instr_i[27] ),
    .A2(\id_stage_i.controller_i.instr_i[29] ),
    .A3(\id_stage_i.controller_i.instr_i[28] ),
    .A4(\id_stage_i.controller_i.instr_i[31] ),
    .ZN(_06958_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _12464_ (.A1(net3649),
    .A2(_06762_),
    .A3(_06766_),
    .A4(_06958_),
    .ZN(_06959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12465_ (.A1(_06957_),
    .A2(_06959_),
    .B(net3648),
    .C(net3416),
    .ZN(_06960_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _12466_ (.A1(_06952_),
    .A2(_06956_),
    .A3(_06960_),
    .ZN(_11003_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12467_ (.I(_11003_[0]),
    .ZN(_11006_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12468_ (.A1(net3648),
    .A2(_06958_),
    .ZN(_06961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12469_ (.A1(net3649),
    .A2(net3646),
    .ZN(_06962_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12470_ (.A1(_06961_),
    .A2(_06962_),
    .B(_06753_),
    .C(_06766_),
    .ZN(_06963_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12471_ (.A1(net3481),
    .A2(_06227_),
    .Z(_06964_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12472_ (.A1(net3474),
    .A2(_06220_),
    .B1(_06213_),
    .B2(_06964_),
    .C(_06392_),
    .ZN(_06965_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12473_ (.A1(_06965_),
    .A2(_06749_),
    .Z(_06966_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12474_ (.A1(net3648),
    .A2(net3486),
    .B(net3480),
    .ZN(_06967_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12475_ (.A1(net3486),
    .A2(_06775_),
    .B(_06967_),
    .C(_06777_),
    .ZN(_06968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12476_ (.A1(net326),
    .A2(_06968_),
    .ZN(_06969_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3401 (.I(_08651_),
    .Z(net3401));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12478_ (.A1(net3648),
    .A2(_06242_),
    .A3(net3646),
    .Z(_06971_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12479_ (.A1(_06761_),
    .A2(_06957_),
    .A3(_06971_),
    .Z(_06972_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12480_ (.A1(_06963_),
    .A2(_06969_),
    .A3(_06966_),
    .A4(_06972_),
    .ZN(_11002_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _12481_ (.I(_11002_[0]),
    .ZN(_11009_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12482_ (.A1(net3648),
    .A2(net3416),
    .Z(_06973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12483_ (.A1(_06973_),
    .A2(net3383),
    .ZN(_06974_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _12484_ (.A1(_06242_),
    .A2(net3416),
    .A3(_06771_),
    .A4(net325),
    .ZN(_06975_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12485_ (.A1(net3649),
    .A2(net3646),
    .Z(_06976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12486_ (.A1(_06319_),
    .A2(net3476),
    .ZN(_06977_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12487_ (.A1(_06771_),
    .A2(_06976_),
    .B(_06350_),
    .C(_06977_),
    .ZN(_06978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12488_ (.A1(net3648),
    .A2(net3416),
    .ZN(_06979_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12489_ (.A1(net3648),
    .A2(_06958_),
    .A3(_06962_),
    .B(_06979_),
    .ZN(_06980_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _12490_ (.A1(_06778_),
    .A2(_06978_),
    .B1(_06980_),
    .B2(_06766_),
    .ZN(_06981_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12491_ (.A1(net353),
    .A2(_06975_),
    .A3(_06981_),
    .Z(_06982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12492_ (.A1(net3469),
    .A2(net266),
    .ZN(_06983_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12493_ (.A1(_06210_),
    .A2(net3473),
    .A3(_06246_),
    .A4(net274),
    .Z(_06984_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12494_ (.A1(net3648),
    .A2(net3473),
    .A3(_06246_),
    .Z(_06985_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12495_ (.A1(net3476),
    .A2(net3648),
    .A3(net3649),
    .A4(net322),
    .Z(_06986_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12496_ (.A1(_06775_),
    .A2(_06984_),
    .B1(_06985_),
    .B2(_06215_),
    .C(_06986_),
    .ZN(_06987_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12497_ (.A1(_06983_),
    .A2(_06987_),
    .ZN(_06988_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12498_ (.A1(_06350_),
    .A2(_06977_),
    .A3(_06765_),
    .Z(_06989_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12499_ (.A1(net3476),
    .A2(net322),
    .A3(_06958_),
    .Z(_06990_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12500_ (.A1(_06219_),
    .A2(_06984_),
    .B1(_06990_),
    .B2(net3416),
    .ZN(_06991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12501_ (.A1(_06317_),
    .A2(_06761_),
    .ZN(_06992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12502_ (.A1(_06989_),
    .A2(_06991_),
    .B(_06992_),
    .ZN(_06993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12503_ (.A1(_06317_),
    .A2(_06215_),
    .ZN(_06994_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12504_ (.A1(_11007_[0]),
    .A2(_06253_),
    .A3(_06994_),
    .A4(_06973_),
    .Z(_06995_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12505_ (.A1(_06995_),
    .A2(_06993_),
    .A3(_06988_),
    .Z(_06996_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12506_ (.A1(_06974_),
    .A2(_06982_),
    .A3(_06996_),
    .Z(_06997_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12507_ (.A1(_06983_),
    .A2(_06987_),
    .Z(_06998_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _12508_ (.A1(_06411_),
    .A2(_06779_),
    .A3(_06771_),
    .A4(_06976_),
    .ZN(_06999_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12509_ (.A1(_06998_),
    .A2(_06999_),
    .Z(_07000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12510_ (.A1(_06979_),
    .A2(net3383),
    .Z(_07001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _12511_ (.A1(_07000_),
    .A2(_06982_),
    .B(_11005_[0]),
    .C(_07001_),
    .ZN(_07002_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12512_ (.A1(_06957_),
    .A2(net353),
    .A3(_06975_),
    .A4(_06981_),
    .Z(_07003_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12513_ (.I(_11012_[0]),
    .ZN(_07004_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12514_ (.A1(_06983_),
    .A2(_06987_),
    .B(_06999_),
    .ZN(_07005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3371 (.I(_07066_),
    .Z(net3371));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12516_ (.A1(_07004_),
    .A2(_07005_),
    .A3(_06993_),
    .Z(_07007_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12517_ (.A1(_07007_),
    .A2(_07003_),
    .ZN(_07008_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12518_ (.A1(_06997_),
    .A2(_07002_),
    .B(_07008_),
    .ZN(_07009_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3340 (.I(_08129_),
    .Z(net3340));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12520_ (.A1(\id_stage_i.controller_i.instr_i[25] ),
    .A2(_06762_),
    .Z(_07011_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _12521_ (.A1(_06777_),
    .A2(net327),
    .A3(_07011_),
    .ZN(_07012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12522_ (.A1(_07009_),
    .A2(_07012_),
    .ZN(_07013_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3334 (.I(net3333),
    .Z(net3334));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12524_ (.I(net3195),
    .ZN(_09746_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12525_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .ZN(_07015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _12526_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .ZN(_07016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12527_ (.A1(_07015_),
    .A2(_07016_),
    .ZN(_07017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3333 (.I(_08488_),
    .Z(net3333));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12529_ (.A1(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .A2(_07017_),
    .ZN(_07019_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12530_ (.A1(_06777_),
    .A2(net327),
    .A3(_07011_),
    .Z(_07020_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3403 (.I(_08649_),
    .Z(net3403));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12532_ (.I0(_11399_[0]),
    .I1(_07019_),
    .S(net3373),
    .Z(_09745_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12533_ (.I(_09745_[0]),
    .ZN(_11015_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3416 (.I(_06409_),
    .Z(net3416));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3414 (.I(_06503_),
    .Z(net3414));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3417 (.I(net3416),
    .Z(net3417));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _12537_ (.I(net3376),
    .ZN(_07025_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3336 (.I(net3335),
    .Z(net3336));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _12539_ (.I(net3658),
    .ZN(_07027_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3421 (.I(_06382_),
    .Z(net3421));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12541_ (.A1(_07015_),
    .A2(_07016_),
    .Z(_07029_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3329 (.I(_08500_),
    .Z(net3329));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12543_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A3(_07017_),
    .Z(_07031_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _12544_ (.A1(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .A2(_07027_),
    .B1(\ex_block_i.alu_i.imd_val_q_i[0] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net334),
    .ZN(_07032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12545_ (.A1(net3655),
    .A2(_07025_),
    .B(_07032_),
    .ZN(_07033_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12546_ (.A1(net3374),
    .A2(_07033_),
    .ZN(_07034_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12547_ (.I(_07034_),
    .ZN(_07035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12548_ (.I0(net3196),
    .I1(net267),
    .S(_06388_),
    .Z(_07036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12549_ (.A1(_07036_),
    .A2(_07035_),
    .ZN(_11014_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12550_ (.I(_11014_[0]),
    .ZN(_09744_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12551_ (.A1(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .A2(_07017_),
    .Z(_07037_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3330 (.I(net3329),
    .Z(net3330));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12553_ (.I0(_11402_[0]),
    .I1(_07037_),
    .S(net3373),
    .Z(_11019_[0]));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12554_ (.A1(_09747_[0]),
    .A2(_11021_[0]),
    .ZN(\alu_adder_result_ex[1] ));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12555_ (.I(\alu_adder_result_ex[1] ),
    .ZN(_11653_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer321 (.I(net3530),
    .Z(net576));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3325 (.I(net3324),
    .Z(net3325));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12558_ (.A1(net3582),
    .A2(_06718_),
    .Z(_07041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12559_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .I1(_07041_),
    .S(_06938_),
    .Z(_07042_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3327 (.I(_08501_),
    .Z(net3327));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12561_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07044_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12562_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07045_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3328 (.I(_08501_),
    .Z(net3328));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12564_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07047_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12565_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07048_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3322 (.I(_08511_),
    .Z(net3322));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3424 (.I(_06382_),
    .Z(net3424));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12568_ (.I0(_07044_),
    .I1(_07045_),
    .I2(_07047_),
    .I3(_07048_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12569_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12570_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(net3622),
    .Z(_07053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12571_ (.A1(net3622),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .Z(_07054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12572_ (.I0(_07053_),
    .I1(_07054_),
    .S(net3467),
    .Z(_07055_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3324 (.I(_08508_),
    .Z(net3324));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12574_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07057_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12575_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07058_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12576_ (.I0(_07052_),
    .I1(_07055_),
    .I2(_07057_),
    .I3(_07058_),
    .S0(net3460),
    .S1(net3578),
    .Z(_07059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12577_ (.I0(_07051_),
    .I1(_07059_),
    .S(_06290_),
    .Z(_07060_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12578_ (.I(net3372),
    .ZN(_07061_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12579_ (.A1(_06884_),
    .A2(_06891_),
    .B(_06354_),
    .C(\cs_registers_i.pc_id_i[2] ),
    .ZN(_07062_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12580_ (.A1(_06938_),
    .A2(_07061_),
    .B(_07062_),
    .ZN(_07063_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3319 (.I(net3317),
    .Z(net3319));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12582_ (.I0(_07042_),
    .I1(_07063_),
    .S(_06313_),
    .Z(_11409_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12583_ (.I(_11409_[0]),
    .ZN(_11413_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12584_ (.A1(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .A2(_07017_),
    .Z(_07065_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12585_ (.A1(_06777_),
    .A2(net327),
    .A3(_07011_),
    .Z(_07066_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3318 (.I(net3317),
    .Z(net3318));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3457 (.I(net3454),
    .Z(net3457));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3455 (.I(net3454),
    .Z(net3455));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3337 (.I(net3336),
    .Z(net3337));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12590_ (.I0(_11409_[0]),
    .I1(_07065_),
    .S(net3370),
    .Z(_11023_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12591_ (.A1(net3580),
    .A2(_06718_),
    .Z(_07071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12592_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .I1(_07071_),
    .S(_06938_),
    .Z(_07072_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12593_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07073_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12594_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07074_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3326 (.I(_08508_),
    .Z(net3326));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12596_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07076_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12597_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07077_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12598_ (.I0(_07073_),
    .I1(_07074_),
    .I2(_07076_),
    .I3(_07077_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07078_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12599_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12600_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net3622),
    .Z(_07080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12601_ (.A1(net3622),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .Z(_07081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12602_ (.I0(_07080_),
    .I1(_07081_),
    .S(net3467),
    .Z(_07082_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12603_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07083_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12604_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_07084_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3315 (.I(net3314),
    .Z(net3315));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12606_ (.I0(_07079_),
    .I1(_07082_),
    .I2(_07083_),
    .I3(_07084_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12607_ (.I0(_07078_),
    .I1(_07086_),
    .S(_06290_),
    .Z(_07087_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12608_ (.I(net3369),
    .ZN(_07088_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12609_ (.A1(_06884_),
    .A2(_06891_),
    .B(_06354_),
    .C(\cs_registers_i.pc_id_i[3] ),
    .ZN(_07089_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12610_ (.A1(_06938_),
    .A2(_07088_),
    .B(_07089_),
    .ZN(_07090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12611_ (.I0(_07072_),
    .I1(_07090_),
    .S(_06313_),
    .Z(_11417_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12612_ (.I(_11417_[0]),
    .ZN(_11421_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12613_ (.A1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A2(_07017_),
    .Z(_07091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12614_ (.I0(_11417_[0]),
    .I1(_07091_),
    .S(net3370),
    .Z(_11027_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12615_ (.A1(\cs_registers_i.pc_id_i[4] ),
    .A2(_06256_),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12616_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S0(net3622),
    .S1(net3596),
    .Z(_07093_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12617_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S0(net3622),
    .S1(net3596),
    .Z(_07094_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12618_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S0(net3620),
    .S1(net3592),
    .Z(_07095_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12619_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .S0(net3620),
    .S1(net3592),
    .Z(_07096_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12620_ (.I0(_07093_),
    .I1(_07094_),
    .I2(_07095_),
    .I3(_07096_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07097_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12621_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S0(net3622),
    .S1(net3596),
    .Z(_07098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12622_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net3622),
    .Z(_07099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12623_ (.A1(net3622),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .Z(_07100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12624_ (.I0(_07099_),
    .I1(_07100_),
    .S(net3465),
    .Z(_07101_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12625_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S0(net3620),
    .S1(net3592),
    .Z(_07102_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12626_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S0(net3620),
    .S1(net3592),
    .Z(_07103_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12627_ (.I0(_07098_),
    .I1(_07101_),
    .I2(_07102_),
    .I3(_07103_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12628_ (.I0(_07097_),
    .I1(_07104_),
    .S(_06290_),
    .Z(_07105_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12629_ (.I(net3368),
    .ZN(_07106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12630_ (.I0(_07092_),
    .I1(_07106_),
    .S(_06892_),
    .Z(_07107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12631_ (.A1(net3576),
    .A2(_06718_),
    .ZN(_07108_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3531 (.I(net314),
    .Z(net3531));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12633_ (.A1(\cs_registers_i.pc_id_i[4] ),
    .A2(_06256_),
    .Z(_07110_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12634_ (.A1(_06917_),
    .A2(_07110_),
    .B(_06354_),
    .ZN(_07111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12635_ (.I(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .ZN(_07112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _12636_ (.A1(_06313_),
    .A2(_07107_),
    .B1(_07108_),
    .B2(_06237_),
    .C1(_07111_),
    .C2(_07112_),
    .ZN(_11425_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12637_ (.I(net3252),
    .ZN(_11429_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12638_ (.A1(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .A2(_07017_),
    .Z(_07113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12639_ (.I0(_11425_[0]),
    .I1(_07113_),
    .S(net3370),
    .Z(_11031_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12640_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[5] ),
    .ZN(_07114_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12641_ (.A1(_06237_),
    .A2(_07114_),
    .B(_06257_),
    .ZN(_07115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3313 (.I(net447),
    .Z(net3313));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12643_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S0(net3619),
    .S1(net3581),
    .Z(_07117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12644_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .S(net3619),
    .Z(_07118_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12645_ (.A1(net3619),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .Z(_07119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12646_ (.I0(_07118_),
    .I1(_07119_),
    .S(net3454),
    .Z(_07120_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3320 (.I(_08515_),
    .Z(net3320));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12648_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S0(net3619),
    .S1(net3581),
    .Z(_07122_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12649_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .S0(net3619),
    .S1(net3581),
    .Z(_07123_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12650_ (.I0(_07117_),
    .I1(_07120_),
    .I2(_07122_),
    .I3(_07123_),
    .S0(net3466),
    .S1(net3578),
    .Z(_07124_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3317 (.I(_08520_),
    .Z(net3317));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12652_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S0(net3616),
    .S1(net3591),
    .Z(_07126_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12653_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S0(net3616),
    .S1(net3591),
    .Z(_07127_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12654_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S0(net3616),
    .S1(net3591),
    .Z(_07128_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12655_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .S0(net3616),
    .S1(net3591),
    .Z(_07129_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12656_ (.I0(_07126_),
    .I1(_07127_),
    .I2(_07128_),
    .I3(_07129_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07130_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12657_ (.A1(_06290_),
    .A2(_07130_),
    .Z(_07131_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12658_ (.A1(net3576),
    .A2(_07124_),
    .B(_07131_),
    .ZN(_07132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12659_ (.A1(_06310_),
    .A2(net3367),
    .ZN(_07133_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12660_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(_06313_),
    .Z(_07134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12661_ (.A1(_07115_),
    .A2(_07133_),
    .A3(_07134_),
    .Z(_11433_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12662_ (.I(_11433_[0]),
    .ZN(_11437_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12663_ (.A1(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .A2(_07017_),
    .Z(_07135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12664_ (.I0(_11433_[0]),
    .I1(_07135_),
    .S(net3370),
    .Z(_11035_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12665_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[6] ),
    .ZN(_07136_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12666_ (.A1(_06237_),
    .A2(_07136_),
    .B(_06257_),
    .ZN(_07137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12667_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S0(net3617),
    .S1(net3592),
    .Z(_07138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12668_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net3633),
    .Z(_07139_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3312 (.I(_08547_),
    .Z(net3312));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12670_ (.A1(net3633),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .Z(_07141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12671_ (.I0(_07139_),
    .I1(_07141_),
    .S(net3465),
    .Z(_07142_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12672_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S0(net3615),
    .S1(net3590),
    .Z(_07143_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12673_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .S0(net3615),
    .S1(net3591),
    .Z(_07144_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12674_ (.I0(_07138_),
    .I1(_07142_),
    .I2(_07143_),
    .I3(_07144_),
    .S0(net3458),
    .S1(net3578),
    .Z(_07145_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3428 (.I(net3427),
    .Z(net3428));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12676_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S0(net3615),
    .S1(net3590),
    .Z(_07147_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12677_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .S0(net3615),
    .S1(net3590),
    .Z(_07148_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12678_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S0(net3615),
    .S1(net3590),
    .Z(_07149_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12679_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .S0(net3615),
    .S1(net3590),
    .Z(_07150_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12680_ (.I0(_07147_),
    .I1(_07148_),
    .I2(_07149_),
    .I3(_07150_),
    .S0(net3464),
    .S1(net3578),
    .Z(_07151_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12681_ (.A1(_06290_),
    .A2(_07151_),
    .Z(_07152_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12682_ (.A1(_07145_),
    .A2(net3576),
    .B(_07152_),
    .ZN(_07153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12683_ (.A1(_06310_),
    .A2(net3366),
    .ZN(_07154_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12684_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(_06313_),
    .Z(_07155_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12685_ (.A1(_07137_),
    .A2(_07154_),
    .A3(_07155_),
    .Z(_11441_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12686_ (.I(_11441_[0]),
    .ZN(_11445_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12687_ (.A1(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A2(_07017_),
    .Z(_07156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12688_ (.I0(_11441_[0]),
    .I1(_07156_),
    .S(net3371),
    .Z(_11039_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12689_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[7] ),
    .ZN(_07157_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12690_ (.A1(_06237_),
    .A2(_07157_),
    .B(_06257_),
    .ZN(_07158_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12691_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S0(net3609),
    .S1(net3591),
    .Z(_07159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12692_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net3609),
    .Z(_07160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12693_ (.A1(net3609),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .Z(_07161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12694_ (.I0(_07160_),
    .I1(_07161_),
    .S(net3466),
    .Z(_07162_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12695_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S0(net3617),
    .S1(net3591),
    .Z(_07163_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12696_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .S0(net3617),
    .S1(net3591),
    .Z(_07164_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12697_ (.I0(_07159_),
    .I1(_07162_),
    .I2(_07163_),
    .I3(_07164_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07165_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12698_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S0(net3608),
    .S1(net3584),
    .Z(_07166_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12699_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S0(net3608),
    .S1(net3584),
    .Z(_07167_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12700_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S0(net3608),
    .S1(net3584),
    .Z(_07168_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12701_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .S0(net3608),
    .S1(net3584),
    .Z(_07169_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12702_ (.I0(_07166_),
    .I1(_07167_),
    .I2(_07168_),
    .I3(_07169_),
    .S0(net3464),
    .S1(net3578),
    .Z(_07170_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12703_ (.A1(_06290_),
    .A2(_07170_),
    .Z(_07171_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12704_ (.A1(net3576),
    .A2(_07165_),
    .B(_07171_),
    .ZN(_07172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12705_ (.A1(_06310_),
    .A2(net3365),
    .ZN(_07173_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12706_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(_06313_),
    .Z(_07174_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12707_ (.A1(_07158_),
    .A2(_07173_),
    .A3(_07174_),
    .Z(_11449_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12708_ (.I(_11449_[0]),
    .ZN(_11453_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12709_ (.I(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .ZN(_07175_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3323 (.I(net3322),
    .Z(net3323));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _12711_ (.A1(_07175_),
    .A2(net3374),
    .A3(_07029_),
    .B1(_11453_[0]),
    .B2(net3373),
    .ZN(_11043_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12712_ (.I(_09747_[0]),
    .ZN(_07177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _12713_ (.A1(_11021_[0]),
    .A2(_07177_),
    .B(_11020_[0]),
    .C(_11024_[0]),
    .ZN(_07178_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12714_ (.A1(_11025_[0]),
    .A2(_11024_[0]),
    .B(_11029_[0]),
    .ZN(_07179_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12715_ (.A1(_11028_[0]),
    .A2(_11032_[0]),
    .ZN(_07180_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12716_ (.I(_11036_[0]),
    .ZN(_07181_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12717_ (.A1(_07178_),
    .A2(_07179_),
    .B(_07180_),
    .C(_07181_),
    .ZN(_07182_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12718_ (.A1(_11032_[0]),
    .A2(_11033_[0]),
    .B(_11037_[0]),
    .ZN(_07183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12719_ (.A1(_07181_),
    .A2(_07183_),
    .ZN(_07184_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12720_ (.A1(_11041_[0]),
    .A2(_07182_),
    .A3(_07184_),
    .Z(_07185_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12721_ (.A1(_11040_[0]),
    .A2(_07185_),
    .ZN(_07186_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12722_ (.A1(net312),
    .A2(_07186_),
    .ZN(net178));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12723_ (.A1(_11017_[0]),
    .A2(net382),
    .A3(net389),
    .A4(net400),
    .Z(_07187_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12724_ (.A1(_11033_[0]),
    .A2(net455),
    .A3(_07187_),
    .Z(_07188_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12725_ (.A1(_06997_),
    .A2(net465),
    .B(net473),
    .C(_07188_),
    .ZN(_07189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12726_ (.I(_11033_[0]),
    .ZN(_07190_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12727_ (.I(_11025_[0]),
    .ZN(_07191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12728_ (.A1(_11021_[0]),
    .A2(_11016_[0]),
    .B(_11020_[0]),
    .ZN(_07192_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _12729_ (.I(_11024_[0]),
    .ZN(_07193_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12730_ (.A1(_07191_),
    .A2(_07192_),
    .B(_07193_),
    .ZN(_07194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12731_ (.A1(net400),
    .A2(_07194_),
    .B(_11028_[0]),
    .ZN(_07195_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12732_ (.I(_11032_[0]),
    .ZN(_07196_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12733_ (.A1(_07190_),
    .A2(_07195_),
    .B(_07196_),
    .ZN(_07197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12734_ (.A1(net455),
    .A2(net350),
    .ZN(_07198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12735_ (.A1(_07181_),
    .A2(_07198_),
    .ZN(_07199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12736_ (.A1(net3373),
    .A2(_07188_),
    .B(_07199_),
    .ZN(_07200_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12737_ (.I(net288),
    .ZN(_07201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12738_ (.A1(_07189_),
    .A2(_07200_),
    .B(_07201_),
    .ZN(_07202_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12739_ (.A1(_07201_),
    .A2(_07189_),
    .A3(_07200_),
    .Z(_07203_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _12740_ (.A1(_07202_),
    .A2(_07203_),
    .ZN(net177));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12741_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[8] ),
    .ZN(_07204_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12742_ (.A1(_06237_),
    .A2(_07204_),
    .B(_06257_),
    .ZN(_07205_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12743_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S0(net3614),
    .S1(net3588),
    .Z(_07206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12744_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net3614),
    .Z(_07207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12745_ (.A1(net3614),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .Z(_07208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12746_ (.I0(_07207_),
    .I1(_07208_),
    .S(net3466),
    .Z(_07209_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3314 (.I(_08535_),
    .Z(net3314));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12748_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S0(net3610),
    .S1(net3585),
    .Z(_07211_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12749_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .S0(net3609),
    .S1(net3585),
    .Z(_07212_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12750_ (.I0(_07206_),
    .I1(_07209_),
    .I2(_07211_),
    .I3(_07212_),
    .S0(net3462),
    .S1(net3578),
    .Z(_07213_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12751_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S0(net333),
    .S1(net3583),
    .Z(_07214_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12752_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07215_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12753_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S0(net3612),
    .S1(net3587),
    .Z(_07216_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12754_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .S0(net3612),
    .S1(net3587),
    .Z(_07217_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12755_ (.I0(_07214_),
    .I1(_07215_),
    .I2(_07216_),
    .I3(_07217_),
    .S0(net3464),
    .S1(net3578),
    .Z(_07218_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12756_ (.A1(_06290_),
    .A2(_07218_),
    .Z(_07219_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12757_ (.A1(_07213_),
    .A2(net3576),
    .B(_07219_),
    .ZN(_07220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12758_ (.A1(_06310_),
    .A2(net3364),
    .ZN(_07221_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12759_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(_06313_),
    .Z(_07222_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12760_ (.A1(_07205_),
    .A2(_07221_),
    .A3(_07222_),
    .Z(_11457_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12761_ (.I(_11457_[0]),
    .ZN(_11461_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12762_ (.A1(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .A2(_07017_),
    .Z(_07223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12763_ (.I0(_11457_[0]),
    .I1(_07223_),
    .S(net3371),
    .Z(_11047_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12764_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[9] ),
    .ZN(_07224_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12765_ (.A1(_06237_),
    .A2(_07224_),
    .B(_06257_),
    .ZN(_07225_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12766_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S0(net3614),
    .S1(net3585),
    .Z(_07226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12767_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(net3609),
    .Z(_07227_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12768_ (.A1(net3609),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .Z(_07228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12769_ (.I0(_07227_),
    .I1(_07228_),
    .S(net3466),
    .Z(_07229_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12770_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S0(net3610),
    .S1(net3585),
    .Z(_07230_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12771_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .S0(net3610),
    .S1(net3585),
    .Z(_07231_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12772_ (.I0(_07226_),
    .I1(_07229_),
    .I2(_07230_),
    .I3(_07231_),
    .S0(net3462),
    .S1(net3578),
    .Z(_07232_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12773_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07233_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12774_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07234_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12775_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07235_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12776_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07236_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12777_ (.I0(_07233_),
    .I1(_07234_),
    .I2(_07235_),
    .I3(_07236_),
    .S0(net3464),
    .S1(net3578),
    .Z(_07237_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12778_ (.A1(_06290_),
    .A2(_07237_),
    .Z(_07238_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12779_ (.A1(_07232_),
    .A2(net3576),
    .B(_07238_),
    .ZN(_07239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12780_ (.A1(_06310_),
    .A2(net3363),
    .ZN(_07240_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12781_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(_06313_),
    .Z(_07241_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12782_ (.A1(_07225_),
    .A2(_07240_),
    .A3(_07241_),
    .Z(_11465_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12783_ (.I(_11465_[0]),
    .ZN(_11469_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12784_ (.A1(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .A2(_07017_),
    .Z(_07242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12785_ (.I0(_11465_[0]),
    .I1(_07242_),
    .S(net3371),
    .Z(_11051_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12786_ (.I(_11021_[0]),
    .ZN(_07243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12787_ (.I(_11020_[0]),
    .ZN(_07244_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _12788_ (.A1(net458),
    .A2(_07243_),
    .B(_07244_),
    .C(_07193_),
    .ZN(_07245_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _12789_ (.I(_07179_),
    .ZN(_07246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12790_ (.A1(_07181_),
    .A2(_07180_),
    .ZN(_07247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12791_ (.A1(_07246_),
    .A2(_07245_),
    .B(_07247_),
    .ZN(_07248_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12792_ (.A1(_11041_[0]),
    .A2(net310),
    .A3(_07184_),
    .ZN(_07249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12793_ (.A1(_11045_[0]),
    .A2(_11040_[0]),
    .ZN(_07250_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12794_ (.I(_11044_[0]),
    .ZN(_07251_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12795_ (.A1(_07248_),
    .A2(_07249_),
    .B(_07250_),
    .C(_07251_),
    .ZN(_07252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12796_ (.A1(_11049_[0]),
    .A2(_07252_),
    .B(_11048_[0]),
    .ZN(_07253_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12797_ (.A1(net315),
    .A2(_07253_),
    .Z(_07254_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _12798_ (.I(_07254_),
    .ZN(net180));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12799_ (.A1(_11041_[0]),
    .A2(_11045_[0]),
    .ZN(_07255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12800_ (.A1(net401),
    .A2(_07197_),
    .B(_11036_[0]),
    .ZN(_07256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12801_ (.A1(net311),
    .A2(_11040_[0]),
    .B(_11044_[0]),
    .ZN(_07257_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12802_ (.A1(net284),
    .A2(_07256_),
    .B(_07257_),
    .ZN(_07258_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12803_ (.A1(net292),
    .A2(net455),
    .A3(_07187_),
    .ZN(_07259_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12804_ (.A1(net305),
    .A2(net3374),
    .B(net284),
    .C(_07259_),
    .ZN(_07260_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12805_ (.A1(net3104),
    .A2(_07260_),
    .B(net293),
    .ZN(_07261_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12806_ (.A1(net293),
    .A2(net3104),
    .A3(_07260_),
    .Z(_07262_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12807_ (.A1(_07261_),
    .A2(_07262_),
    .Z(net179));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12808_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[10] ),
    .ZN(_07263_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12809_ (.A1(_06237_),
    .A2(_07263_),
    .B(_06257_),
    .ZN(_07264_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12810_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S0(net3608),
    .S1(net3584),
    .Z(_07265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12811_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .S(net3609),
    .Z(_07266_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12812_ (.A1(net3609),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .Z(_07267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12813_ (.I0(_07266_),
    .I1(_07267_),
    .S(net3466),
    .Z(_07268_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12814_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S0(net3609),
    .S1(net3585),
    .Z(_07269_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12815_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .S0(net3609),
    .S1(net3585),
    .Z(_07270_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12816_ (.I0(_07265_),
    .I1(_07268_),
    .I2(_07269_),
    .I3(_07270_),
    .S0(net3462),
    .S1(net3578),
    .Z(_07271_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12817_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07272_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12818_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07273_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12819_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07274_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12820_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .S0(net3611),
    .S1(net3586),
    .Z(_07275_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12821_ (.I0(_07272_),
    .I1(_07273_),
    .I2(_07274_),
    .I3(_07275_),
    .S0(net3464),
    .S1(net3578),
    .Z(_07276_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12822_ (.A1(_06290_),
    .A2(_07276_),
    .Z(_07277_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12823_ (.A1(net3576),
    .A2(_07271_),
    .B(_07277_),
    .ZN(_07278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12824_ (.A1(_06310_),
    .A2(net3362),
    .ZN(_07279_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12825_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(_06313_),
    .Z(_07280_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12826_ (.A1(_07264_),
    .A2(_07279_),
    .A3(_07280_),
    .Z(_11473_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12827_ (.I(_11473_[0]),
    .ZN(_11477_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12828_ (.A1(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .A2(_07017_),
    .Z(_07281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12829_ (.I0(_11473_[0]),
    .I1(_07281_),
    .S(net3371),
    .Z(_11055_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12830_ (.I(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .ZN(_07282_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _12831_ (.A1(_07282_),
    .A2(net3374),
    .A3(_07029_),
    .B1(net3373),
    .B2(_11485_[0]),
    .ZN(_11059_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _12832_ (.I(_11049_[0]),
    .ZN(_07283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12833_ (.A1(_11057_[0]),
    .A2(_11052_[0]),
    .B(_11056_[0]),
    .C(_11048_[0]),
    .ZN(_07284_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12834_ (.A1(_07283_),
    .A2(_07251_),
    .B(_07284_),
    .ZN(_07285_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12835_ (.A1(_07283_),
    .A2(_07250_),
    .ZN(_07286_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12836_ (.A1(_07285_),
    .A2(_07286_),
    .ZN(_07287_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _12837_ (.A1(net318),
    .A2(_07248_),
    .A3(_07249_),
    .B(_07287_),
    .ZN(_07288_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12838_ (.A1(_11053_[0]),
    .A2(_11052_[0]),
    .Z(_07289_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12839_ (.A1(net281),
    .A2(_07289_),
    .Z(_07290_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12840_ (.A1(_07290_),
    .A2(_11056_[0]),
    .Z(_07291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12841_ (.A1(_07288_),
    .A2(_07291_),
    .ZN(_07292_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12842_ (.A1(_11061_[0]),
    .A2(_07292_),
    .ZN(net152));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12843_ (.A1(_06974_),
    .A2(_06982_),
    .A3(net332),
    .ZN(_07293_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _12844_ (.A1(net353),
    .A2(_06975_),
    .A3(_06981_),
    .ZN(_07294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12845_ (.A1(_06979_),
    .A2(net3383),
    .ZN(_07295_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12846_ (.I(_11005_[0]),
    .ZN(_07296_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12847_ (.A1(_07005_),
    .A2(_07294_),
    .B(_07295_),
    .C(_07296_),
    .ZN(_07297_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12848_ (.A1(net292),
    .A2(net455),
    .A3(net288),
    .A4(_11045_[0]),
    .Z(_07298_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12849_ (.A1(_07187_),
    .A2(_07298_),
    .Z(_07299_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12850_ (.I(_07299_),
    .ZN(_07300_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _12851_ (.A1(_07293_),
    .A2(_07297_),
    .B1(_07003_),
    .B2(_07007_),
    .C(_07300_),
    .ZN(_07301_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12852_ (.A1(net3373),
    .A2(_07299_),
    .Z(_07302_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12853_ (.A1(_11052_[0]),
    .A2(_07258_),
    .A3(_11048_[0]),
    .Z(_07303_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12854_ (.A1(_07303_),
    .A2(_07301_),
    .A3(_07302_),
    .Z(_07304_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12855_ (.A1(net294),
    .A2(_11048_[0]),
    .A3(_11052_[0]),
    .Z(_07305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12856_ (.A1(_07289_),
    .A2(_07305_),
    .Z(_07306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12857_ (.I(net281),
    .ZN(_07307_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12858_ (.A1(net286),
    .A2(_07306_),
    .B(_07307_),
    .ZN(_07308_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12859_ (.A1(_07307_),
    .A2(net286),
    .A3(_07306_),
    .Z(_07309_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12860_ (.A1(_07308_),
    .A2(_07309_),
    .Z(net151));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3316 (.I(_08527_),
    .Z(net3316));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12862_ (.A1(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .A2(_07017_),
    .Z(_07311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12863_ (.I0(_11494_[0]),
    .I1(_07311_),
    .S(net3371),
    .Z(_11063_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3427 (.I(_06367_),
    .Z(net3427));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3309 (.I(net481),
    .Z(net3309));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3310 (.I(_08558_),
    .Z(net3310));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3321 (.I(_08511_),
    .Z(net3321));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3311 (.I(net3310),
    .Z(net3311));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3303 (.I(_08583_),
    .Z(net3303));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place3307 (.I(_08573_),
    .Z(net3307));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3306 (.I(net3304),
    .Z(net3306));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12872_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S0(net3574),
    .S1(net3549),
    .Z(_07320_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3298 (.I(_08600_),
    .Z(net3298));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3293 (.I(_08613_),
    .Z(net3293));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3292 (.I(_08615_),
    .Z(net3292));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12876_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S0(net3574),
    .S1(net3549),
    .Z(_07324_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12877_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S0(net3574),
    .S1(net3551),
    .Z(_07325_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12878_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S0(net3574),
    .S1(net3551),
    .Z(_07326_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3297 (.I(net3296),
    .Z(net3297));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3294 (.I(net3293),
    .Z(net3294));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3291 (.I(_08662_),
    .Z(net3291));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3296 (.I(_08605_),
    .Z(net3296));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12883_ (.I0(_07320_),
    .I1(_07324_),
    .I2(_07325_),
    .I3(_07326_),
    .S0(net3437),
    .S1(net3490),
    .Z(_07331_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12884_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S0(net3574),
    .S1(net3551),
    .Z(_07332_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3304 (.I(_08578_),
    .Z(net3304));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3302 (.I(net3301),
    .Z(net3302));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12887_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(net3550),
    .Z(_07335_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3290 (.I(_02398_),
    .Z(net3290));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3289 (.I(_02570_),
    .Z(net3289));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12890_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .A2(_06334_),
    .A3(net314),
    .Z(_07338_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12891_ (.A1(_07335_),
    .A2(net3574),
    .B(_07338_),
    .ZN(_07339_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12892_ (.I(_07339_),
    .ZN(_07340_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12893_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S0(net3574),
    .S1(net3551),
    .Z(_07341_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12894_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S0(net3574),
    .S1(net3551),
    .Z(_07342_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12895_ (.I0(_07332_),
    .I1(_07340_),
    .I2(_07341_),
    .I3(_07342_),
    .S0(net3434),
    .S1(net3493),
    .Z(_07343_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3287 (.I(_11430_[0]),
    .Z(net3287));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3301 (.I(_08586_),
    .Z(net3301));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12898_ (.I0(_07331_),
    .I1(_07343_),
    .S(net3421),
    .Z(_07346_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12899_ (.A1(net3479),
    .A2(_06396_),
    .Z(_07347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12900_ (.A1(_06465_),
    .A2(_07347_),
    .ZN(_07348_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _12901_ (.A1(_06806_),
    .A2(_06459_),
    .A3(_06465_),
    .B(_06396_),
    .ZN(_07349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12902_ (.A1(net320),
    .A2(_07349_),
    .ZN(_07350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12903_ (.A1(_07348_),
    .A2(_07350_),
    .ZN(_07351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12904_ (.I0(net420),
    .I1(_07351_),
    .S(_06441_),
    .Z(_11493_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12905_ (.I(_11493_[0]),
    .ZN(_11489_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12906_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[13] ),
    .ZN(_07352_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12907_ (.A1(_06237_),
    .A2(_07352_),
    .B(net3352),
    .ZN(_07353_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3456 (.I(net3454),
    .Z(net3456));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12909_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S0(net3640),
    .S1(net3602),
    .Z(_07355_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12910_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S0(net3640),
    .S1(net3602),
    .Z(_07356_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer305 (.I(net3115),
    .Z(net560));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12912_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S0(net3640),
    .S1(net3597),
    .Z(_07358_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12913_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .S0(net3640),
    .S1(net3597),
    .Z(_07359_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12914_ (.I0(_07355_),
    .I1(_07356_),
    .I2(_07358_),
    .I3(_07359_),
    .S0(net3461),
    .S1(net3578),
    .Z(_07360_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12915_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S0(net3640),
    .S1(net3601),
    .Z(_07361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12916_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net3640),
    .Z(_07362_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12917_ (.A1(net3640),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .Z(_07363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12918_ (.I0(_07362_),
    .I1(_07363_),
    .S(net3468),
    .Z(_07364_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12919_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S0(net3640),
    .S1(net3596),
    .Z(_07365_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12920_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S0(net3640),
    .S1(net3596),
    .Z(_07366_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12921_ (.I0(_07361_),
    .I1(_07364_),
    .I2(_07365_),
    .I3(_07366_),
    .S0(net3459),
    .S1(net3579),
    .Z(_07367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12922_ (.I0(_07360_),
    .I1(_07367_),
    .S(_06290_),
    .Z(_07368_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12923_ (.I(net3361),
    .ZN(_07369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12924_ (.A1(_06310_),
    .A2(_07369_),
    .ZN(_07370_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12925_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(_06313_),
    .Z(_07371_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12926_ (.A1(_07353_),
    .A2(_07370_),
    .A3(_07371_),
    .Z(_11502_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _12927_ (.I(_11502_[0]),
    .ZN(_11498_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _12928_ (.I(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .ZN(_07372_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _12929_ (.A1(_07372_),
    .A2(net3374),
    .A3(_07029_),
    .B1(_11498_[0]),
    .B2(net3373),
    .ZN(_11067_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3300 (.I(net3298),
    .Z(net3300));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3286 (.I(_11003_[0]),
    .Z(net3286));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12932_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S0(net3574),
    .S1(net3549),
    .Z(_07375_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12933_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S0(net3574),
    .S1(net3549),
    .Z(_07376_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 place3530 (.I(net3513),
    .Z(net3530));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12935_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S0(net3574),
    .S1(net3551),
    .Z(_07378_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12936_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .S0(net3574),
    .S1(net3551),
    .Z(_07379_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12937_ (.I0(_07375_),
    .I1(_07376_),
    .I2(_07378_),
    .I3(_07379_),
    .S0(net3437),
    .S1(net3490),
    .Z(_07380_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12938_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S0(net3569),
    .S1(net3543),
    .Z(_07381_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3295 (.I(_08605_),
    .Z(net3295));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12940_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net3541),
    .Z(_07383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12941_ (.A1(net3541),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .Z(_07384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12942_ (.I0(_07383_),
    .I1(_07384_),
    .S(net3446),
    .Z(_07385_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12943_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S0(net3569),
    .S1(net3541),
    .Z(_07386_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12944_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S0(net3569),
    .S1(net3541),
    .Z(_07387_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12945_ (.I0(_07381_),
    .I1(_07385_),
    .I2(_07386_),
    .I3(_07387_),
    .S0(net3434),
    .S1(net3492),
    .Z(_07388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12946_ (.I0(_07380_),
    .I1(_07388_),
    .S(net3422),
    .Z(_07389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12947_ (.A1(net3648),
    .A2(_07349_),
    .ZN(_07390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12948_ (.A1(_07348_),
    .A2(_07390_),
    .ZN(_07391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12949_ (.I0(net424),
    .I1(_07391_),
    .S(_06441_),
    .Z(_11501_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12950_ (.I(_11501_[0]),
    .ZN(_11497_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3433 (.I(_06367_),
    .Z(net3433));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3494 (.I(net3490),
    .Z(net3494));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12953_ (.A1(_11061_[0]),
    .A2(net3187),
    .A3(_07291_),
    .Z(_07394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _12954_ (.A1(net394),
    .A2(_11060_[0]),
    .B1(_07394_),
    .B2(_07288_),
    .C(_11064_[0]),
    .ZN(_07395_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12955_ (.A1(_11069_[0]),
    .A2(net399),
    .ZN(net154));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12956_ (.A1(_11056_[0]),
    .A2(_11061_[0]),
    .B(_11060_[0]),
    .ZN(_07396_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12957_ (.A1(net315),
    .A2(_11048_[0]),
    .Z(_07397_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12958_ (.A1(_11061_[0]),
    .A2(net281),
    .Z(_07398_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12959_ (.A1(_11052_[0]),
    .A2(_07397_),
    .B(_07398_),
    .ZN(_07399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12960_ (.A1(net359),
    .A2(_07399_),
    .ZN(_07400_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12961_ (.A1(net393),
    .A2(_07258_),
    .A3(_07400_),
    .Z(_07401_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12962_ (.A1(_07301_),
    .A2(_07302_),
    .A3(_07401_),
    .Z(_07402_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12963_ (.A1(net294),
    .A2(net315),
    .A3(_07398_),
    .Z(_07403_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12964_ (.A1(_07301_),
    .A2(_07302_),
    .B(_07403_),
    .C(net393),
    .ZN(_07404_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12965_ (.A1(_07400_),
    .A2(_07403_),
    .Z(_07405_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12966_ (.A1(net3104),
    .A2(_07403_),
    .B(_07400_),
    .ZN(_07406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12967_ (.I0(_07405_),
    .I1(_07406_),
    .S(net393),
    .Z(_07407_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12968_ (.A1(_07402_),
    .A2(_07404_),
    .A3(_07407_),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12969_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[14] ),
    .ZN(_07408_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12970_ (.A1(_06237_),
    .A2(_07408_),
    .B(net3352),
    .ZN(_07409_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12971_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S0(net3618),
    .S1(net3581),
    .Z(_07410_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12972_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .S0(net3618),
    .S1(net3581),
    .Z(_07411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12973_ (.I0(_07410_),
    .I1(_07411_),
    .S(net3466),
    .Z(_07412_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12974_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S0(net3618),
    .S1(net3588),
    .Z(_07413_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12975_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S0(net3618),
    .S1(net3588),
    .Z(_07414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12976_ (.I0(_07413_),
    .I1(_07414_),
    .S(net3455),
    .Z(_07415_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _12977_ (.I(net3578),
    .ZN(_07416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12978_ (.I0(_07412_),
    .I1(_07415_),
    .S(_07416_),
    .Z(_07417_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12979_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S0(net3621),
    .S1(net3593),
    .Z(_07418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12980_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(net3616),
    .Z(_07419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12981_ (.A1(net3618),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .Z(_07420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12982_ (.I0(_07419_),
    .I1(_07420_),
    .S(net3466),
    .Z(_07421_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12983_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S0(net3616),
    .S1(net3593),
    .Z(_07422_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12984_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S0(net3621),
    .S1(net3593),
    .Z(_07423_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12985_ (.I0(_07418_),
    .I1(_07421_),
    .I2(_07422_),
    .I3(_07423_),
    .S0(net3455),
    .S1(net3578),
    .Z(_07424_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12986_ (.A1(_06290_),
    .A2(_07424_),
    .Z(_07425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12987_ (.A1(_07417_),
    .A2(net3576),
    .B(_07425_),
    .ZN(_07426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12988_ (.A1(_06310_),
    .A2(net3351),
    .ZN(_07427_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12989_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(_06313_),
    .Z(_07428_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12990_ (.A1(_07409_),
    .A2(_07427_),
    .A3(_07428_),
    .Z(_11510_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12991_ (.I(_11510_[0]),
    .ZN(_11506_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12992_ (.A1(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .A2(_07017_),
    .Z(_07429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12993_ (.I0(_11510_[0]),
    .I1(_07429_),
    .S(net3371),
    .Z(_11071_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3461 (.I(net3454),
    .Z(net3461));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3285 (.I(net451),
    .Z(net3285));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12996_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S0(net3557),
    .S1(net3523),
    .Z(_07432_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12997_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S0(net3557),
    .S1(net3523),
    .Z(_07433_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3468 (.I(net3467),
    .Z(net3468));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3283 (.I(_08512_),
    .Z(net3283));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3280 (.I(_08524_),
    .Z(net3280));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13001_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S0(net3557),
    .S1(net3523),
    .Z(_07437_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13002_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .S0(net3557),
    .S1(net3523),
    .Z(_07438_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3277 (.I(_08528_),
    .Z(net3277));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13004_ (.I0(_07432_),
    .I1(_07433_),
    .I2(_07437_),
    .I3(_07438_),
    .S0(net3444),
    .S1(net3496),
    .Z(_07440_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13005_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S0(net3557),
    .S1(net3523),
    .Z(_07441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13006_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(net3523),
    .Z(_07442_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13007_ (.A1(net3523),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .Z(_07443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13008_ (.I0(_07442_),
    .I1(_07443_),
    .S(net3453),
    .Z(_07444_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13009_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S0(net3557),
    .S1(net3523),
    .Z(_07445_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13010_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S0(net3557),
    .S1(net3523),
    .Z(_07446_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3279 (.I(net3278),
    .Z(net3279));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13012_ (.I0(_07441_),
    .I1(_07444_),
    .I2(_07445_),
    .I3(_07446_),
    .S0(net3444),
    .S1(net3496),
    .Z(_07448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13013_ (.I0(_07440_),
    .I1(_07448_),
    .S(net3424),
    .Z(_07449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13014_ (.A1(net3647),
    .A2(_07349_),
    .ZN(_07450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13015_ (.A1(_07348_),
    .A2(_07450_),
    .ZN(_07451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13016_ (.I0(_07449_),
    .I1(_07451_),
    .S(_06441_),
    .Z(_11509_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13017_ (.I(_11509_[0]),
    .ZN(_11505_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13018_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(net3394),
    .Z(_07452_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13019_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S0(net444),
    .S1(net3594),
    .Z(_07453_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place3276 (.I(net3275),
    .Z(net3276));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13021_ (.A1(net3456),
    .A2(net3594),
    .ZN(_07455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13022_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net444),
    .Z(_07456_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13023_ (.A1(net3456),
    .A2(_07453_),
    .B1(_07455_),
    .B2(_07456_),
    .C(_07416_),
    .ZN(_07457_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13024_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S0(net444),
    .S1(net3594),
    .Z(_07458_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13025_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S0(net444),
    .S1(net3594),
    .Z(_07459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13026_ (.I0(_07458_),
    .I1(_07459_),
    .S(net3456),
    .Z(_07460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13027_ (.A1(net3578),
    .A2(_07460_),
    .ZN(_07461_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13028_ (.A1(_07457_),
    .A2(_07461_),
    .Z(_07462_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13029_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S0(net3632),
    .S1(net3594),
    .Z(_07463_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13030_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S0(net3632),
    .S1(net3594),
    .Z(_07464_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13031_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S0(net3632),
    .S1(net3594),
    .Z(_07465_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13032_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .S0(net3632),
    .S1(net3594),
    .Z(_07466_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13033_ (.I0(_07463_),
    .I1(_07464_),
    .I2(_07465_),
    .I3(_07466_),
    .S0(net3456),
    .S1(net3578),
    .Z(_07467_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13034_ (.A1(_06290_),
    .A2(_07467_),
    .ZN(_07468_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13035_ (.A1(net444),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .B(_06735_),
    .ZN(_07469_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13036_ (.A1(_06290_),
    .A2(_07462_),
    .B(_07468_),
    .C(_07469_),
    .ZN(_07470_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13037_ (.A1(_06310_),
    .A2(net3350),
    .Z(_07471_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13038_ (.A1(\cs_registers_i.pc_id_i[15] ),
    .A2(_06313_),
    .A3(_06938_),
    .Z(_07472_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13039_ (.A1(_07452_),
    .A2(_07471_),
    .A3(_07472_),
    .Z(_11518_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _13040_ (.I(_11518_[0]),
    .ZN(_11514_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13041_ (.A1(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .A2(_07017_),
    .Z(_07473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13042_ (.I0(_11518_[0]),
    .I1(_07473_),
    .S(net3373),
    .Z(_11075_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13043_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S0(net3564),
    .S1(net3523),
    .Z(_07474_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13044_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S0(net3564),
    .S1(net3523),
    .Z(_07475_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13045_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S0(net3564),
    .S1(net3523),
    .Z(_07476_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13046_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .S0(net3564),
    .S1(net3523),
    .Z(_07477_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13047_ (.I0(_07474_),
    .I1(_07475_),
    .I2(_07476_),
    .I3(_07477_),
    .S0(net3444),
    .S1(net3496),
    .Z(_07478_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13048_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S0(net3564),
    .S1(net3523),
    .Z(_07479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13049_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net3523),
    .Z(_07480_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13050_ (.A1(net3523),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .Z(_07481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13051_ (.I0(_07480_),
    .I1(_07481_),
    .S(net3453),
    .Z(_07482_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13052_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S0(net3564),
    .S1(net3523),
    .Z(_07483_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13053_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S0(net3564),
    .S1(net3523),
    .Z(_07484_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13054_ (.I0(_07479_),
    .I1(_07482_),
    .I2(_07483_),
    .I3(_07484_),
    .S0(net3444),
    .S1(net3496),
    .Z(_07485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13055_ (.I0(_07478_),
    .I1(_07485_),
    .S(net3424),
    .Z(_07486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13056_ (.A1(net3607),
    .A2(_07349_),
    .ZN(_07487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13057_ (.A1(_07348_),
    .A2(_07487_),
    .ZN(_07488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13058_ (.I0(_07486_),
    .I1(_07488_),
    .S(_06441_),
    .Z(_11517_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13059_ (.I(_11517_[0]),
    .ZN(_11513_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13060_ (.A1(_07181_),
    .A2(_07183_),
    .B(_07255_),
    .ZN(_07489_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13061_ (.A1(_07489_),
    .A2(_11049_[0]),
    .Z(_07490_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13062_ (.A1(_07286_),
    .A2(_07285_),
    .Z(_07491_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13063_ (.A1(_07182_),
    .A2(_07490_),
    .B(_07491_),
    .ZN(_07492_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _13064_ (.A1(net348),
    .A2(net3187),
    .A3(_07291_),
    .ZN(_07493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13065_ (.A1(net3187),
    .A2(_11060_[0]),
    .ZN(_07494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13066_ (.I(_11064_[0]),
    .ZN(_07495_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _13067_ (.A1(_07492_),
    .A2(_07493_),
    .B(_07494_),
    .C(_07495_),
    .ZN(_07496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13068_ (.A1(_11069_[0]),
    .A2(_07496_),
    .Z(_07497_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13069_ (.A1(_11068_[0]),
    .A2(_07497_),
    .Z(_07498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13070_ (.A1(net3186),
    .A2(_07498_),
    .B(_11072_[0]),
    .ZN(_07499_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _13071_ (.A1(net271),
    .A2(_07499_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13072_ (.A1(_07304_),
    .A2(_07306_),
    .Z(_07500_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _13073_ (.A1(net3187),
    .A2(_11069_[0]),
    .A3(net3186),
    .A4(_07398_),
    .Z(_07501_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13074_ (.I(_11065_[0]),
    .ZN(_07502_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13075_ (.A1(_07502_),
    .A2(_07396_),
    .B(_07495_),
    .ZN(_07503_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13076_ (.A1(_11069_[0]),
    .A2(_07503_),
    .Z(_07504_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13077_ (.A1(_11068_[0]),
    .A2(_07504_),
    .Z(_07505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13078_ (.A1(net388),
    .A2(_07306_),
    .B(_07505_),
    .C(net3186),
    .ZN(_07506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13079_ (.A1(net3187),
    .A2(_11069_[0]),
    .B(net3186),
    .ZN(_07507_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13080_ (.A1(_11069_[0]),
    .A2(_07503_),
    .B(_11068_[0]),
    .ZN(_07508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13081_ (.I0(net3186),
    .I1(_07507_),
    .S(net352),
    .Z(_07509_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13082_ (.A1(net3186),
    .A2(_07398_),
    .A3(_07505_),
    .ZN(_07510_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13083_ (.A1(_07509_),
    .A2(_07510_),
    .Z(_07511_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13084_ (.A1(_07500_),
    .A2(_07501_),
    .B(_07506_),
    .C(_07511_),
    .ZN(net155));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13085_ (.I(\cs_registers_i.pc_id_i[16] ),
    .ZN(_07512_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13086_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S0(net3629),
    .S1(net3597),
    .Z(_07513_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13087_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .S0(net3629),
    .S1(net3597),
    .Z(_07514_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13088_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S0(net3629),
    .S1(net3597),
    .Z(_07515_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13089_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S0(net3629),
    .S1(net3597),
    .Z(_07516_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13090_ (.I0(_07513_),
    .I1(_07514_),
    .I2(_07515_),
    .I3(_07516_),
    .S0(net3457),
    .S1(net3578),
    .Z(_07517_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13091_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S0(net3629),
    .S1(net3595),
    .Z(_07518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13092_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(net3624),
    .Z(_07519_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13093_ (.A1(net3624),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .Z(_07520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13094_ (.I0(_07519_),
    .I1(_07520_),
    .S(net3467),
    .Z(_07521_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13095_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S0(net3629),
    .S1(net3595),
    .Z(_07522_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13096_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S0(net3629),
    .S1(net3595),
    .Z(_07523_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13097_ (.I0(_07518_),
    .I1(_07521_),
    .I2(_07522_),
    .I3(_07523_),
    .S0(net3457),
    .S1(net3578),
    .Z(_07524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13098_ (.I0(_07517_),
    .I1(_07524_),
    .S(_06290_),
    .Z(_07525_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _13099_ (.I(net3360),
    .ZN(_07526_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _13100_ (.A1(_07512_),
    .A2(_06892_),
    .B1(_07526_),
    .B2(net3352),
    .ZN(_07527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13101_ (.A1(_06313_),
    .A2(_07527_),
    .ZN(_07528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13102_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(net3394),
    .ZN(_07529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13103_ (.A1(_07528_),
    .A2(_07529_),
    .ZN(_11526_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _13104_ (.I(_11526_[0]),
    .ZN(_11522_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13105_ (.A1(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .A2(_07017_),
    .Z(_07530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13106_ (.I0(_11526_[0]),
    .I1(_07530_),
    .S(net3373),
    .Z(_11079_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3272 (.I(_08540_),
    .Z(net3272));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13108_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S0(net3565),
    .S1(net3529),
    .Z(_07532_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13109_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .S0(net3565),
    .S1(net3529),
    .Z(_07533_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13110_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S0(net3563),
    .S1(net3529),
    .Z(_07534_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13111_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S0(net3565),
    .S1(net3529),
    .Z(_07535_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13112_ (.I0(_07532_),
    .I1(_07533_),
    .I2(_07534_),
    .I3(_07535_),
    .S0(net3432),
    .S1(net3491),
    .Z(_07536_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13113_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S0(net3565),
    .S1(net3529),
    .Z(_07537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13114_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(net3529),
    .Z(_07538_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13115_ (.A1(net3529),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .Z(_07539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13116_ (.I0(_07538_),
    .I1(_07539_),
    .S(net3453),
    .Z(_07540_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13117_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S0(net3565),
    .S1(net3529),
    .Z(_07541_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13118_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S0(net3565),
    .S1(net3529),
    .Z(_07542_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13119_ (.I0(_07537_),
    .I1(_07540_),
    .I2(_07541_),
    .I3(_07542_),
    .S0(net3432),
    .S1(net3491),
    .Z(_07543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13120_ (.I0(_07536_),
    .I1(_07543_),
    .S(net3423),
    .Z(_07544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13121_ (.A1(net3605),
    .A2(_07349_),
    .ZN(_07545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13122_ (.A1(_07348_),
    .A2(_07545_),
    .ZN(_07546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13123_ (.I0(_07544_),
    .I1(_07546_),
    .S(_06441_),
    .Z(_11525_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13124_ (.I(_11525_[0]),
    .ZN(_11521_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13125_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(net3394),
    .ZN(_07547_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13126_ (.A1(net333),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .Z(_07548_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13127_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .S0(net3624),
    .S1(net3593),
    .Z(_07549_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13128_ (.A1(net3581),
    .A2(_07549_),
    .Z(_07550_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13129_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S0(net3624),
    .S1(net3593),
    .Z(_07551_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13130_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S0(net3624),
    .S1(net3593),
    .Z(_07552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13131_ (.I0(_07551_),
    .I1(_07552_),
    .S(net3454),
    .Z(_07553_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13132_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S0(net3631),
    .S1(net3593),
    .Z(_07554_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13133_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .S0(net3631),
    .S1(net3593),
    .Z(_07555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13134_ (.I0(_07554_),
    .I1(_07555_),
    .S(net3454),
    .Z(_07556_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13135_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S0(net3630),
    .S1(net3589),
    .Z(_07557_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13136_ (.A1(net3454),
    .A2(_07557_),
    .Z(_07558_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13137_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net333),
    .Z(_07559_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13138_ (.A1(net3581),
    .A2(_06275_),
    .A3(_07559_),
    .Z(_07560_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13139_ (.A1(_07558_),
    .A2(_07560_),
    .Z(_07561_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _13140_ (.I0(_07550_),
    .I1(_07553_),
    .I2(_07556_),
    .I3(_07561_),
    .S0(_07416_),
    .S1(_06290_),
    .Z(_07562_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13141_ (.A1(_07416_),
    .A2(_07551_),
    .Z(_07563_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13142_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S0(net3624),
    .S1(net3593),
    .Z(_07564_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _13143_ (.A1(_06290_),
    .A2(net3454),
    .A3(_07563_),
    .A4(_07564_),
    .Z(_07565_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _13144_ (.A1(_06735_),
    .A2(_07548_),
    .B(_07565_),
    .C(_07562_),
    .ZN(_07566_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13145_ (.A1(net3352),
    .A2(_06917_),
    .A3(net3349),
    .Z(_07567_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13146_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(_06313_),
    .A3(_06938_),
    .ZN(_07568_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _13147_ (.A1(_07547_),
    .A2(_07567_),
    .A3(_07568_),
    .ZN(_11534_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13148_ (.I(_11534_[0]),
    .ZN(_11530_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13149_ (.A1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .A2(_07017_),
    .Z(_07569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13150_ (.I0(_11534_[0]),
    .I1(_07569_),
    .S(net3373),
    .Z(_11083_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13151_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S0(net3563),
    .S1(net3528),
    .Z(_07570_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13152_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S0(net3563),
    .S1(net3528),
    .Z(_07571_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13153_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S0(net3563),
    .S1(net3528),
    .Z(_07572_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13154_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .S0(net3563),
    .S1(net3528),
    .Z(_07573_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13155_ (.I0(_07570_),
    .I1(_07571_),
    .I2(_07572_),
    .I3(_07573_),
    .S0(net3431),
    .S1(net3491),
    .Z(_07574_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13156_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S0(net3563),
    .S1(net3528),
    .Z(_07575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13157_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net3540),
    .Z(_07576_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13158_ (.A1(net3540),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .Z(_07577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13159_ (.I0(_07576_),
    .I1(_07577_),
    .S(net3448),
    .Z(_07578_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13160_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S0(net3563),
    .S1(net3528),
    .Z(_07579_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13161_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .S0(net3563),
    .S1(net3528),
    .Z(_07580_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13162_ (.I0(_07575_),
    .I1(_07578_),
    .I2(_07579_),
    .I3(_07580_),
    .S0(net3431),
    .S1(net3491),
    .Z(_07581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13163_ (.I0(_07574_),
    .I1(_07581_),
    .S(net3423),
    .Z(_07582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13164_ (.A1(net3582),
    .A2(_07349_),
    .ZN(_07583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13165_ (.A1(_07348_),
    .A2(_07583_),
    .ZN(_07584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13166_ (.I0(_07582_),
    .I1(_07584_),
    .S(_06441_),
    .Z(_11533_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13167_ (.I(_11533_[0]),
    .ZN(_11529_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13168_ (.I(_11077_[0]),
    .ZN(_07585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13169_ (.A1(_11073_[0]),
    .A2(_11068_[0]),
    .B(_11072_[0]),
    .ZN(_07586_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13170_ (.I(_11076_[0]),
    .ZN(_07587_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13171_ (.A1(_07586_),
    .A2(_07585_),
    .B(_07587_),
    .ZN(_07588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13172_ (.A1(_11081_[0]),
    .A2(_07588_),
    .B(_11080_[0]),
    .ZN(_07589_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13173_ (.A1(net3186),
    .A2(net271),
    .A3(_11081_[0]),
    .Z(_07590_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13174_ (.A1(_11069_[0]),
    .A2(_07496_),
    .A3(_07590_),
    .ZN(_07591_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13175_ (.A1(_07589_),
    .A2(_07591_),
    .Z(_07592_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13176_ (.A1(_11085_[0]),
    .A2(_07592_),
    .ZN(net158));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _13177_ (.A1(net3187),
    .A2(_11069_[0]),
    .A3(net3186),
    .A4(net271),
    .Z(_07593_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13178_ (.A1(_11081_[0]),
    .A2(_07489_),
    .A3(_07403_),
    .A4(_07593_),
    .Z(_07594_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13179_ (.A1(_07187_),
    .A2(_07594_),
    .Z(_07595_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13180_ (.I(_07595_),
    .ZN(_07596_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13181_ (.A1(net305),
    .A2(_07596_),
    .Z(_07597_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13182_ (.A1(net3186),
    .A2(net271),
    .ZN(_07598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13183_ (.A1(_11069_[0]),
    .A2(_11064_[0]),
    .B(_11068_[0]),
    .ZN(_07599_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13184_ (.A1(net271),
    .A2(_11072_[0]),
    .B(_11076_[0]),
    .ZN(_07600_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13185_ (.A1(_07598_),
    .A2(_07599_),
    .B(_07600_),
    .ZN(_07601_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13186_ (.A1(_07405_),
    .A2(_07593_),
    .Z(_07602_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13187_ (.I(_07257_),
    .ZN(_07603_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13188_ (.A1(_07603_),
    .A2(_07403_),
    .Z(_07604_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13189_ (.A1(_07400_),
    .A2(_07604_),
    .Z(_07605_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13190_ (.A1(_07593_),
    .A2(_07605_),
    .Z(_07606_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13191_ (.A1(net379),
    .A2(_07606_),
    .B(_11081_[0]),
    .ZN(_07607_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13192_ (.A1(_11081_[0]),
    .A2(net379),
    .A3(_07602_),
    .B(_07607_),
    .ZN(_07608_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13193_ (.A1(_07199_),
    .A2(_07594_),
    .B1(_07595_),
    .B2(net3371),
    .C(_07608_),
    .ZN(_07609_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13194_ (.A1(_11081_[0]),
    .A2(_07258_),
    .A3(_07400_),
    .A4(net379),
    .Z(_07610_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13195_ (.A1(_07301_),
    .A2(_07302_),
    .A3(_07610_),
    .Z(_07611_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13196_ (.A1(_07609_),
    .A2(_07597_),
    .A3(_07611_),
    .Z(net157));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13197_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S0(net3634),
    .S1(net3597),
    .Z(_07612_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13198_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S0(net3634),
    .S1(net3597),
    .Z(_07613_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13199_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S0(net3634),
    .S1(net3597),
    .Z(_07614_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13200_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S0(net3634),
    .S1(net3597),
    .Z(_07615_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13201_ (.I0(_07612_),
    .I1(_07613_),
    .I2(_07614_),
    .I3(_07615_),
    .S0(net3461),
    .S1(net3579),
    .Z(_07616_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13202_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S0(net3634),
    .S1(net3601),
    .Z(_07617_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13203_ (.A1(net480),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .Z(_07618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13204_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(net3634),
    .Z(_07619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13205_ (.I0(_07618_),
    .I1(_07619_),
    .S(net3601),
    .Z(_07620_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13206_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S0(net3634),
    .S1(net3601),
    .Z(_07621_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13207_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S0(net3634),
    .S1(net3601),
    .Z(_07622_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13208_ (.I0(_07617_),
    .I1(_07620_),
    .I2(_07621_),
    .I3(_07622_),
    .S0(net3459),
    .S1(net3579),
    .Z(_07623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13209_ (.I0(_07616_),
    .I1(_07623_),
    .S(_06290_),
    .Z(_07624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13210_ (.A1(_06208_),
    .A2(_06256_),
    .Z(_07625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13211_ (.A1(\cs_registers_i.pc_id_i[18] ),
    .A2(_06938_),
    .B1(net3359),
    .B2(_07625_),
    .ZN(_07626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13212_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(net3394),
    .ZN(_07627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13213_ (.A1(_06917_),
    .A2(_07626_),
    .B(_07627_),
    .ZN(_11542_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13214_ (.I(_11542_[0]),
    .ZN(_11538_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13215_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(_07017_),
    .Z(_07628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13216_ (.I0(_11542_[0]),
    .I1(_07628_),
    .S(net3373),
    .Z(_11087_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13217_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S0(net3573),
    .S1(net3543),
    .Z(_07629_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13218_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S0(net3573),
    .S1(net3543),
    .Z(_07630_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13219_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S0(net3573),
    .S1(net3543),
    .Z(_07631_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13220_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S0(net3573),
    .S1(net3543),
    .Z(_07632_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13221_ (.I0(_07629_),
    .I1(_07630_),
    .I2(_07631_),
    .I3(_07632_),
    .S0(net3438),
    .S1(net3492),
    .Z(_07633_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13222_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S0(net3573),
    .S1(net3543),
    .Z(_07634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13223_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(net3543),
    .Z(_07635_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13224_ (.A1(net3543),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .Z(_07636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13225_ (.I0(_07635_),
    .I1(_07636_),
    .S(net3447),
    .Z(_07637_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13226_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S0(net3573),
    .S1(net3543),
    .Z(_07638_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13227_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S0(net3573),
    .S1(net3543),
    .Z(_07639_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13228_ (.I0(_07634_),
    .I1(_07637_),
    .I2(_07638_),
    .I3(_07639_),
    .S0(net3435),
    .S1(net3492),
    .Z(_07640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13229_ (.I0(_07633_),
    .I1(_07640_),
    .S(net3422),
    .Z(_07641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13230_ (.A1(net3580),
    .A2(_07349_),
    .ZN(_07642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13231_ (.A1(_07348_),
    .A2(_07642_),
    .ZN(_07643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13232_ (.I0(net414),
    .I1(_07643_),
    .S(_06441_),
    .Z(_11541_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13233_ (.I(_11541_[0]),
    .ZN(_11537_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13234_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[19] ),
    .ZN(_07644_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13235_ (.A1(net3353),
    .A2(_07644_),
    .B(net3352),
    .ZN(_07645_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13236_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S0(net3644),
    .S1(net3597),
    .Z(_07646_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13237_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S0(net3644),
    .S1(net3597),
    .Z(_07647_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13238_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S0(net3644),
    .S1(net3597),
    .Z(_07648_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13239_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .S0(net3644),
    .S1(net3597),
    .Z(_07649_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _13240_ (.I0(_07646_),
    .I1(_07647_),
    .I2(_07648_),
    .I3(_07649_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07650_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13241_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S0(net3644),
    .S1(net3597),
    .Z(_07651_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13242_ (.A1(net333),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .Z(_07652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13243_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .S(net449),
    .Z(_07653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13244_ (.I0(_07652_),
    .I1(_07653_),
    .S(net3597),
    .Z(_07654_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13245_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S0(net3643),
    .S1(net3597),
    .Z(_07655_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13246_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S0(net3643),
    .S1(net3597),
    .Z(_07656_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13247_ (.I0(_07651_),
    .I1(_07654_),
    .I2(_07655_),
    .I3(_07656_),
    .S0(net3454),
    .S1(net3578),
    .Z(_07657_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13248_ (.A1(net3576),
    .A2(_07657_),
    .Z(_07658_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13249_ (.A1(_06290_),
    .A2(_07650_),
    .B(_07658_),
    .ZN(_07659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13250_ (.A1(_06310_),
    .A2(net3348),
    .ZN(_07660_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13251_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(_06313_),
    .Z(_07661_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13252_ (.A1(_07645_),
    .A2(_07660_),
    .A3(_07661_),
    .Z(_11550_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _13253_ (.I(_11550_[0]),
    .ZN(_11546_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13254_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(_07017_),
    .Z(_07662_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3271 (.I(net3270),
    .Z(net3271));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13256_ (.I0(_11550_[0]),
    .I1(_07662_),
    .S(net3371),
    .Z(_11091_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13257_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S0(net3575),
    .S1(net3549),
    .Z(_07664_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13258_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S0(net3575),
    .S1(net3549),
    .Z(_07665_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13259_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S0(net3575),
    .S1(net3549),
    .Z(_07666_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13260_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .S0(net3575),
    .S1(net3548),
    .Z(_07667_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13261_ (.I0(_07664_),
    .I1(_07665_),
    .I2(_07666_),
    .I3(_07667_),
    .S0(net3439),
    .S1(net3494),
    .Z(_07668_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13262_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S0(net3575),
    .S1(net3549),
    .Z(_07669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13263_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .S(net3549),
    .Z(_07670_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13264_ (.A1(net3549),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .Z(_07671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13265_ (.I0(_07670_),
    .I1(_07671_),
    .S(net3445),
    .Z(_07672_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13266_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S0(net3575),
    .S1(net3549),
    .Z(_07673_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13267_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S0(net3575),
    .S1(net3549),
    .Z(_07674_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13268_ (.I0(_07669_),
    .I1(_07672_),
    .I2(_07673_),
    .I3(_07674_),
    .S0(net3436),
    .S1(net3494),
    .Z(_07675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13269_ (.I0(_07668_),
    .I1(_07675_),
    .S(net3423),
    .Z(_07676_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13270_ (.A1(net3576),
    .A2(_07349_),
    .ZN(_07677_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13271_ (.A1(_07348_),
    .A2(_07677_),
    .ZN(_07678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13272_ (.I0(net441),
    .I1(_07678_),
    .S(_06441_),
    .Z(_11549_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13273_ (.I(_11549_[0]),
    .ZN(_11545_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13274_ (.A1(_11069_[0]),
    .A2(_11085_[0]),
    .A3(_11089_[0]),
    .A4(_07590_),
    .Z(_07679_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place3275 (.I(_08533_),
    .Z(net3275));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13276_ (.I(_11085_[0]),
    .ZN(_07681_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13277_ (.I(_11084_[0]),
    .ZN(_07682_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13278_ (.A1(_07589_),
    .A2(_07681_),
    .B(_07682_),
    .ZN(_07683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13279_ (.A1(_11089_[0]),
    .A2(_07683_),
    .Z(_07684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13280_ (.A1(_07496_),
    .A2(_07679_),
    .B(_07684_),
    .C(_11088_[0]),
    .ZN(_07685_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13281_ (.A1(_11093_[0]),
    .A2(_07685_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13282_ (.A1(_11081_[0]),
    .A2(_11085_[0]),
    .Z(_07686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13283_ (.A1(_07593_),
    .A2(_07686_),
    .Z(_07687_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13284_ (.A1(_11089_[0]),
    .A2(_07398_),
    .A3(_07687_),
    .Z(_07688_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13285_ (.A1(_11085_[0]),
    .A2(_11080_[0]),
    .Z(_07689_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13286_ (.A1(_07508_),
    .A2(_07598_),
    .B(_07600_),
    .ZN(_07690_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13287_ (.A1(_07686_),
    .A2(_07690_),
    .Z(_07691_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13288_ (.A1(_11084_[0]),
    .A2(_07689_),
    .A3(_07691_),
    .Z(_07692_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _13289_ (.A1(_07304_),
    .A2(_07306_),
    .B(_07692_),
    .C(_11089_[0]),
    .ZN(_07693_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13290_ (.A1(_11089_[0]),
    .A2(_07692_),
    .A3(_07687_),
    .ZN(_07694_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13291_ (.A1(_11089_[0]),
    .A2(_07692_),
    .B(_07694_),
    .ZN(_07695_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13292_ (.A1(_11089_[0]),
    .A2(_07398_),
    .A3(_07692_),
    .B(_07695_),
    .ZN(_07696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13293_ (.A1(_07500_),
    .A2(_07688_),
    .B(_07696_),
    .C(_07693_),
    .ZN(net159));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13294_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[20] ),
    .ZN(_07697_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13295_ (.A1(net3353),
    .A2(_07697_),
    .B(net3352),
    .ZN(_07698_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13296_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S0(net3634),
    .S1(net3597),
    .Z(_07699_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13297_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S0(net480),
    .S1(net3597),
    .Z(_07700_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13298_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S0(net480),
    .S1(net3596),
    .Z(_07701_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13299_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S0(net480),
    .S1(net3596),
    .Z(_07702_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13300_ (.I0(_07699_),
    .I1(_07700_),
    .I2(_07701_),
    .I3(_07702_),
    .S0(net3459),
    .S1(net3579),
    .Z(_07703_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13301_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S0(net480),
    .S1(net3596),
    .Z(_07704_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13302_ (.A1(net480),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .Z(_07705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13303_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net3634),
    .Z(_07706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13304_ (.I0(_07705_),
    .I1(_07706_),
    .S(net3596),
    .Z(_07707_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13305_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S0(net3641),
    .S1(net3596),
    .Z(_07708_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13306_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S0(net3641),
    .S1(net3596),
    .Z(_07709_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13307_ (.I0(_07704_),
    .I1(_07707_),
    .I2(_07708_),
    .I3(_07709_),
    .S0(net3459),
    .S1(net3579),
    .Z(_07710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13308_ (.I0(_07703_),
    .I1(_07710_),
    .S(_06290_),
    .Z(_07711_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _13309_ (.I(net3358),
    .ZN(_07712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13310_ (.A1(_06310_),
    .A2(_07712_),
    .ZN(_07713_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13311_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(_06313_),
    .Z(_07714_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13312_ (.A1(_07698_),
    .A2(_07713_),
    .A3(_07714_),
    .Z(_11558_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13313_ (.I(_11558_[0]),
    .ZN(_11554_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13314_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(_07017_),
    .Z(_07715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13315_ (.I0(_11558_[0]),
    .I1(_07715_),
    .S(net3371),
    .Z(_11095_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3504 (.I(net3503),
    .Z(net3504));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13317_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S0(net3569),
    .S1(net3544),
    .Z(_07717_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13318_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S0(net3569),
    .S1(net3544),
    .Z(_07718_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3268 (.I(_08562_),
    .Z(net3268));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3267 (.I(_08566_),
    .Z(net3267));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13321_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S0(net3569),
    .S1(net3544),
    .Z(_07721_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3509 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(net3509));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13323_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S0(net3569),
    .S1(net3544),
    .Z(_07723_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13324_ (.I0(_07717_),
    .I1(_07718_),
    .I2(_07721_),
    .I3(_07723_),
    .S0(net3435),
    .S1(net3492),
    .Z(_07724_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13325_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S0(net3569),
    .S1(net3544),
    .Z(_07725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13326_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net3543),
    .Z(_07726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13327_ (.A1(net3543),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .Z(_07727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13328_ (.I0(_07726_),
    .I1(_07727_),
    .S(net3447),
    .Z(_07728_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13329_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S0(net3569),
    .S1(net3543),
    .Z(_07729_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13330_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S0(net3569),
    .S1(net3543),
    .Z(_07730_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13331_ (.I0(_07725_),
    .I1(_07728_),
    .I2(_07729_),
    .I3(_07730_),
    .S0(net3435),
    .S1(net3492),
    .Z(_07731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13332_ (.I0(_07724_),
    .I1(_07731_),
    .S(net3422),
    .Z(_07732_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3266 (.I(net3265),
    .Z(net3266));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13334_ (.A1(_06459_),
    .A2(_06395_),
    .Z(_07734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3503 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(net3503));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13336_ (.A1(_06354_),
    .A2(_06463_),
    .Z(_07736_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13337_ (.A1(_07736_),
    .A2(_07347_),
    .Z(_07737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13338_ (.A1(net3560),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_07738_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13339_ (.I(_07738_),
    .ZN(_07739_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3273 (.I(net3272),
    .Z(net3273));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _13341_ (.A1(net3380),
    .A2(net410),
    .B1(_07739_),
    .B2(net3379),
    .ZN(_11553_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13342_ (.I(_11553_[0]),
    .ZN(_11557_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13343_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[21] ),
    .ZN(_07741_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13344_ (.A1(net3353),
    .A2(_07741_),
    .B(net3352),
    .ZN(_07742_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13345_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .S0(net3642),
    .S1(net3581),
    .Z(_07743_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13346_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .S0(net3642),
    .S1(net3581),
    .Z(_07744_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13347_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S0(net3642),
    .S1(net3581),
    .Z(_07745_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13348_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S0(net3642),
    .S1(net3581),
    .Z(_07746_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _13349_ (.I0(_07743_),
    .I1(_07744_),
    .I2(_07745_),
    .I3(_07746_),
    .S0(net3578),
    .S1(net3596),
    .Z(_07747_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13350_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S0(net3642),
    .S1(net3599),
    .Z(_07748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13351_ (.A1(net3622),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .Z(_07749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13352_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net3622),
    .Z(_07750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13353_ (.I0(_07749_),
    .I1(_07750_),
    .S(net3599),
    .Z(_07751_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13354_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S0(net3622),
    .S1(net3599),
    .Z(_07752_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13355_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S0(net3642),
    .S1(net3599),
    .Z(_07753_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13356_ (.I0(_07748_),
    .I1(_07751_),
    .I2(_07752_),
    .I3(_07753_),
    .S0(net3460),
    .S1(net3578),
    .Z(_07754_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13357_ (.A1(net3577),
    .A2(_07754_),
    .Z(_07755_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13358_ (.A1(_06290_),
    .A2(_07747_),
    .B(_07755_),
    .ZN(_07756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13359_ (.A1(_06310_),
    .A2(net3347),
    .ZN(_07757_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13360_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(_06313_),
    .Z(_07758_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13361_ (.A1(_07742_),
    .A2(_07757_),
    .A3(_07758_),
    .Z(_11566_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13362_ (.I(_11566_[0]),
    .ZN(_11562_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13363_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(_07017_),
    .Z(_07759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13364_ (.I0(_11566_[0]),
    .I1(_07759_),
    .S(net3371),
    .Z(_11099_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13365_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S0(net3570),
    .S1(net3542),
    .Z(_07760_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13366_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .S0(net3570),
    .S1(net3542),
    .Z(_07761_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3263 (.I(_08571_),
    .Z(net3263));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3467 (.I(_06275_),
    .Z(net3467));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13369_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S0(net3570),
    .S1(net3542),
    .Z(_07764_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13370_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .S0(net3570),
    .S1(net3542),
    .Z(_07765_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3466 (.I(_06275_),
    .Z(net3466));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3579 (.I(net3578),
    .Z(net3579));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13373_ (.I0(_07760_),
    .I1(_07761_),
    .I2(_07764_),
    .I3(_07765_),
    .S0(net3433),
    .S1(net3493),
    .Z(_07768_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13374_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S0(net3575),
    .S1(net3549),
    .Z(_07769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13375_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net3549),
    .Z(_07770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13376_ (.A1(net3548),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .Z(_07771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13377_ (.I0(_07770_),
    .I1(_07771_),
    .S(net3445),
    .Z(_07772_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13378_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S0(net3575),
    .S1(net3548),
    .Z(_07773_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13379_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S0(net3575),
    .S1(net3548),
    .Z(_07774_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13380_ (.I0(_07769_),
    .I1(_07772_),
    .I2(_07773_),
    .I3(_07774_),
    .S0(net3433),
    .S1(net3493),
    .Z(_07775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13381_ (.I0(_07768_),
    .I1(_07775_),
    .S(net3421),
    .Z(_07776_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3534 (.I(net3513),
    .Z(net3534));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13383_ (.A1(net3531),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_07778_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13384_ (.I(_07778_),
    .ZN(_07779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13385_ (.A1(net3380),
    .A2(net442),
    .B1(_07779_),
    .B2(net3379),
    .ZN(_11561_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13386_ (.I(_11561_[0]),
    .ZN(_11565_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13387_ (.I(_11097_[0]),
    .ZN(_07780_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _13388_ (.A1(_11069_[0]),
    .A2(_11085_[0]),
    .A3(_11089_[0]),
    .A4(_07590_),
    .ZN(_07781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13389_ (.A1(_11089_[0]),
    .A2(net316),
    .B(_11088_[0]),
    .ZN(_07782_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13390_ (.A1(_07781_),
    .A2(_07395_),
    .B(_07782_),
    .ZN(_07783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13391_ (.A1(_07783_),
    .A2(_11093_[0]),
    .B(_11092_[0]),
    .ZN(_07784_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13392_ (.I(_11096_[0]),
    .ZN(_07785_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13393_ (.A1(_07780_),
    .A2(_07784_),
    .B(_07785_),
    .ZN(_07786_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13394_ (.A1(_07786_),
    .A2(_11101_[0]),
    .ZN(_07787_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _13395_ (.I(_07787_),
    .ZN(net162));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _13396_ (.A1(net290),
    .A2(net471),
    .B(net472),
    .C(_07299_),
    .ZN(_07788_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13397_ (.A1(net3373),
    .A2(_07299_),
    .ZN(_07789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13398_ (.A1(_11089_[0]),
    .A2(_11093_[0]),
    .ZN(_07790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _13399_ (.A1(_07601_),
    .A2(_07686_),
    .B(_07689_),
    .C(_11084_[0]),
    .ZN(_07791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13400_ (.A1(_11093_[0]),
    .A2(_11088_[0]),
    .B(_11092_[0]),
    .ZN(_07792_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13401_ (.A1(_07791_),
    .A2(_07790_),
    .B(_07792_),
    .ZN(_07793_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _13402_ (.A1(net349),
    .A2(_07400_),
    .A3(_07793_),
    .ZN(_07794_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13403_ (.A1(_07788_),
    .A2(_07789_),
    .A3(_07794_),
    .Z(_07795_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13404_ (.A1(_11089_[0]),
    .A2(_11093_[0]),
    .A3(_07687_),
    .Z(_07796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13405_ (.A1(_07405_),
    .A2(_07796_),
    .B(net378),
    .ZN(_07797_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13406_ (.A1(_07795_),
    .A2(net386),
    .B(net343),
    .ZN(_07798_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13407_ (.A1(net343),
    .A2(_07795_),
    .A3(net386),
    .Z(_07799_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13408_ (.A1(_07798_),
    .A2(_07799_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13409_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[22] ),
    .ZN(_07800_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13410_ (.A1(net3353),
    .A2(_07800_),
    .B(net3352),
    .ZN(_07801_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13411_ (.A1(net3627),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .Z(_07802_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13412_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S0(net3627),
    .S1(net3597),
    .Z(_07803_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13413_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S0(net3627),
    .S1(net3597),
    .Z(_07804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13414_ (.I0(_07803_),
    .I1(_07804_),
    .S(net3454),
    .Z(_07805_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13415_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S0(net3628),
    .S1(net3597),
    .Z(_07806_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13416_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .S0(net3627),
    .S1(net3604),
    .Z(_07807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13417_ (.I0(_07806_),
    .I1(_07807_),
    .S(net3454),
    .Z(_07808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13418_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .S(net3628),
    .Z(_07809_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13419_ (.A1(net3454),
    .A2(_07809_),
    .Z(_07810_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13420_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S0(net3628),
    .S1(net3581),
    .Z(_07811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13421_ (.I0(_07810_),
    .I1(_07811_),
    .S(net3604),
    .Z(_07812_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13422_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S0(net3627),
    .S1(net3603),
    .Z(_07813_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13423_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S0(net3627),
    .S1(net3604),
    .Z(_07814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13424_ (.I0(_07813_),
    .I1(_07814_),
    .S(net3454),
    .Z(_07815_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _13425_ (.I0(_07805_),
    .I1(_07808_),
    .I2(_07812_),
    .I3(_07815_),
    .S0(net3578),
    .S1(_06290_),
    .Z(_07816_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13426_ (.A1(_06735_),
    .A2(_07802_),
    .B(_07816_),
    .ZN(_07817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13427_ (.A1(_06310_),
    .A2(net3346),
    .ZN(_07818_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13428_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(_06313_),
    .Z(_07819_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13429_ (.A1(_07801_),
    .A2(_07818_),
    .A3(_07819_),
    .Z(_11574_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13430_ (.I(_11574_[0]),
    .ZN(_11570_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13431_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(_07017_),
    .Z(_07820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13432_ (.I0(_11574_[0]),
    .I1(_07820_),
    .S(net3371),
    .Z(_11103_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3617 (.I(net3616),
    .Z(net3617));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3265 (.I(_08570_),
    .Z(net3265));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13435_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S0(net3563),
    .S1(net576),
    .Z(_07823_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3274 (.I(_08533_),
    .Z(net3274));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3258 (.I(net3257),
    .Z(net3258));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13438_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S0(net3563),
    .S1(net576),
    .Z(_07826_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13439_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S0(net3563),
    .S1(net576),
    .Z(_07827_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13440_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .S0(net3563),
    .S1(net576),
    .Z(_07828_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13441_ (.I0(_07823_),
    .I1(_07826_),
    .I2(_07827_),
    .I3(_07828_),
    .S0(net3427),
    .S1(net3491),
    .Z(_07829_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3578 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .Z(net3578));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13443_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S0(net3563),
    .S1(net3530),
    .Z(_07831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13444_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .S(net3530),
    .Z(_07832_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13445_ (.A1(net3530),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .Z(_07833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13446_ (.I0(_07832_),
    .I1(_07833_),
    .S(net3453),
    .Z(_07834_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13447_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S0(net3563),
    .S1(net3530),
    .Z(_07835_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13448_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S0(net3563),
    .S1(net3530),
    .Z(_07836_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13449_ (.I0(_07831_),
    .I1(_07834_),
    .I2(_07835_),
    .I3(_07836_),
    .S0(net3427),
    .S1(net3491),
    .Z(_07837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13450_ (.I0(_07829_),
    .I1(_07837_),
    .S(net3423),
    .Z(_07838_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13452_ (.A1(net3508),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_07840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13453_ (.I(_07840_),
    .ZN(_07841_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _13454_ (.A1(net3380),
    .A2(_07838_),
    .B1(_07841_),
    .B2(net3379),
    .ZN(_11569_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13455_ (.I(_11569_[0]),
    .ZN(_11573_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13456_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[23] ),
    .ZN(_07842_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13457_ (.A1(net3353),
    .A2(_07842_),
    .B(net3352),
    .ZN(_07843_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13458_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .S0(net3614),
    .S1(net3581),
    .Z(_07844_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13459_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S0(net3614),
    .S1(net3581),
    .Z(_07845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13460_ (.I0(_07844_),
    .I1(_07845_),
    .S(net3588),
    .Z(_07846_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13461_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S0(net3614),
    .S1(net3588),
    .Z(_07847_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13462_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S0(net3614),
    .S1(net3588),
    .Z(_07848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13463_ (.I0(_07847_),
    .I1(_07848_),
    .S(net3455),
    .Z(_07849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13464_ (.I0(_07846_),
    .I1(_07849_),
    .S(_07416_),
    .Z(_07850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13465_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .S(net3616),
    .Z(_07851_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13466_ (.A1(net3616),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .Z(_07852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13467_ (.I0(_07851_),
    .I1(_07852_),
    .S(net3454),
    .Z(_07853_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13468_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .S0(net3616),
    .S1(net3581),
    .Z(_07854_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13469_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S0(net3616),
    .S1(net3581),
    .Z(_07855_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13470_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S0(net3616),
    .S1(net3581),
    .Z(_07856_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13471_ (.I0(_07853_),
    .I1(_07854_),
    .I2(_07855_),
    .I3(_07856_),
    .S0(net3578),
    .S1(net3591),
    .Z(_07857_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13472_ (.A1(_06290_),
    .A2(_07857_),
    .Z(_07858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13473_ (.A1(_07850_),
    .A2(net3576),
    .B(_07858_),
    .ZN(_07859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13474_ (.A1(_06310_),
    .A2(net3345),
    .ZN(_07860_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13475_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(_06313_),
    .Z(_07861_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13476_ (.A1(_07843_),
    .A2(_07860_),
    .A3(_07861_),
    .Z(_11582_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _13477_ (.I(_11582_[0]),
    .ZN(_11578_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13478_ (.I(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .ZN(_07862_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _13479_ (.A1(_07862_),
    .A2(net3375),
    .A3(_07029_),
    .B1(_11578_[0]),
    .B2(net3373),
    .ZN(_11107_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13480_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S0(net3556),
    .S1(net3522),
    .Z(_07863_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13481_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S0(net3556),
    .S1(net3519),
    .Z(_07864_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13482_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S0(net3556),
    .S1(net3522),
    .Z(_07865_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13483_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .S0(net3556),
    .S1(net3522),
    .Z(_07866_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13484_ (.I0(_07863_),
    .I1(_07864_),
    .I2(_07865_),
    .I3(_07866_),
    .S0(net3443),
    .S1(net3496),
    .Z(_07867_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13485_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S0(net3556),
    .S1(net3521),
    .Z(_07868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13486_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(net3521),
    .Z(_07869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13487_ (.A1(net3521),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .Z(_07870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13488_ (.I0(_07869_),
    .I1(_07870_),
    .S(net3453),
    .Z(_07871_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13489_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S0(net3556),
    .S1(net3522),
    .Z(_07872_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13490_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S0(net3556),
    .S1(net3522),
    .Z(_07873_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13491_ (.I0(_07868_),
    .I1(_07871_),
    .I2(_07872_),
    .I3(_07873_),
    .S0(net3443),
    .S1(net3496),
    .Z(_07874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13492_ (.I0(_07867_),
    .I1(_07874_),
    .S(net3424),
    .Z(_07875_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13494_ (.A1(net3497),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_07877_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13495_ (.I(_07877_),
    .ZN(_07878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _13496_ (.A1(net3380),
    .A2(_07875_),
    .B1(_07878_),
    .B2(net3379),
    .ZN(_11577_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13497_ (.I(_11577_[0]),
    .ZN(_11581_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13498_ (.A1(_11097_[0]),
    .A2(_11101_[0]),
    .Z(_07879_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13499_ (.A1(_11105_[0]),
    .A2(_07879_),
    .Z(_07880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13500_ (.A1(_11093_[0]),
    .A2(_07880_),
    .Z(_07881_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13501_ (.I(_11104_[0]),
    .ZN(_07882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13502_ (.A1(_11097_[0]),
    .A2(_11092_[0]),
    .ZN(_07883_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13503_ (.I(_11101_[0]),
    .ZN(_07884_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13504_ (.A1(_07785_),
    .A2(_07883_),
    .B(_07884_),
    .ZN(_07885_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13505_ (.A1(_11100_[0]),
    .A2(_07885_),
    .B(_11105_[0]),
    .ZN(_07886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13506_ (.A1(_07882_),
    .A2(_07886_),
    .ZN(_07887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13507_ (.A1(_07881_),
    .A2(_07783_),
    .B(_07887_),
    .ZN(_07888_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _13508_ (.A1(_07888_),
    .A2(_11109_[0]),
    .ZN(net164));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13509_ (.A1(net462),
    .A2(_11096_[0]),
    .B(_11100_[0]),
    .ZN(_07889_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _13510_ (.A1(_07690_),
    .A2(_07686_),
    .B(_07689_),
    .C(_11084_[0]),
    .ZN(_07890_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13511_ (.A1(_07890_),
    .A2(_07790_),
    .B(_07792_),
    .ZN(_07891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13512_ (.A1(_07879_),
    .A2(net632),
    .ZN(_07892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13513_ (.A1(_07889_),
    .A2(_07892_),
    .ZN(_07893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _13514_ (.A1(net287),
    .A2(_07306_),
    .B(_07893_),
    .C(_11105_[0]),
    .ZN(_07894_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13515_ (.A1(_07796_),
    .A2(_07879_),
    .Z(_07895_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13516_ (.A1(_11105_[0]),
    .A2(_07398_),
    .Z(_07896_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _13517_ (.A1(net287),
    .A2(_07306_),
    .A3(_07895_),
    .A4(_07896_),
    .Z(_07897_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _13518_ (.I(_11105_[0]),
    .ZN(_07898_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13519_ (.A1(_11105_[0]),
    .A2(_07895_),
    .Z(_07899_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _13520_ (.A1(_11101_[0]),
    .A2(_11096_[0]),
    .B1(_07891_),
    .B2(_07879_),
    .C(_11100_[0]),
    .ZN(_07900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13521_ (.I0(_07898_),
    .I1(_07899_),
    .S(_07900_),
    .Z(_07901_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13522_ (.A1(_11105_[0]),
    .A2(_07398_),
    .A3(_07893_),
    .B(_07901_),
    .ZN(_07902_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _13523_ (.A1(_07894_),
    .A2(_07897_),
    .A3(_07902_),
    .ZN(net163));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13524_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[24] ),
    .ZN(_07903_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13525_ (.A1(net3353),
    .A2(_07903_),
    .B(net3352),
    .ZN(_07904_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13526_ (.A1(net3625),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .Z(_07905_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13527_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S0(net3632),
    .S1(net3594),
    .Z(_07906_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13528_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .S0(net444),
    .S1(net3594),
    .Z(_07907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13529_ (.I0(_07906_),
    .I1(_07907_),
    .S(net3456),
    .Z(_07908_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13530_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S0(net3632),
    .S1(net3594),
    .Z(_07909_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13531_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .S0(net3632),
    .S1(net3594),
    .Z(_07910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13532_ (.I0(_07909_),
    .I1(_07910_),
    .S(net3456),
    .Z(_07911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13533_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .S(net3632),
    .Z(_07912_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13534_ (.A1(net3456),
    .A2(_07912_),
    .Z(_07913_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13535_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S0(net3632),
    .S1(net3581),
    .Z(_07914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13536_ (.I0(_07913_),
    .I1(_07914_),
    .S(net3594),
    .Z(_07915_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13537_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S0(net444),
    .S1(net3594),
    .Z(_07916_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13538_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .S0(net444),
    .S1(net3594),
    .Z(_07917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13539_ (.I0(_07916_),
    .I1(_07917_),
    .S(net3456),
    .Z(_07918_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _13540_ (.I0(_07908_),
    .I1(_07911_),
    .I2(_07915_),
    .I3(_07918_),
    .S0(net3578),
    .S1(_06290_),
    .Z(_07919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13541_ (.A1(_06735_),
    .A2(_07905_),
    .B(_07919_),
    .ZN(_07920_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13542_ (.A1(_06310_),
    .A2(net3344),
    .ZN(_07921_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13543_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(_06313_),
    .Z(_07922_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13544_ (.A1(_07904_),
    .A2(_07921_),
    .A3(_07922_),
    .Z(_11590_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13545_ (.I(_11590_[0]),
    .ZN(_11586_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13546_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(_07017_),
    .Z(_07923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13547_ (.I0(_11590_[0]),
    .I1(_07923_),
    .S(net3371),
    .Z(_11111_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13548_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S0(net3558),
    .S1(net314),
    .Z(_07924_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13549_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .S0(net3558),
    .S1(net314),
    .Z(_07925_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13550_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S0(net3558),
    .S1(net314),
    .Z(_07926_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13551_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .S0(net3558),
    .S1(net314),
    .Z(_07927_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13552_ (.I0(_07924_),
    .I1(_07925_),
    .I2(_07926_),
    .I3(_07927_),
    .S0(_06367_),
    .S1(net3496),
    .Z(_07928_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13553_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S0(net3558),
    .S1(net3524),
    .Z(_07929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13554_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .S(net314),
    .Z(_07930_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13555_ (.A1(net314),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .Z(_07931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13556_ (.I0(_07930_),
    .I1(_07931_),
    .S(_06334_),
    .Z(_07932_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13557_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S0(net3558),
    .S1(net3524),
    .Z(_07933_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13558_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .S0(net3558),
    .S1(net314),
    .Z(_07934_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13559_ (.I0(_07929_),
    .I1(_07932_),
    .I2(_07933_),
    .I3(_07934_),
    .S0(_06367_),
    .S1(net3496),
    .Z(_07935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13560_ (.I0(_07928_),
    .I1(_07935_),
    .S(net3424),
    .Z(_07936_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3264 (.I(net3263),
    .Z(net3264));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13562_ (.A1(net3489),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_07938_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13563_ (.I(_07938_),
    .ZN(_07939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _13564_ (.A1(net3380),
    .A2(_07936_),
    .B1(_07939_),
    .B2(net3379),
    .ZN(_11585_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13565_ (.I(_11585_[0]),
    .ZN(_11589_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13566_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[25] ),
    .ZN(_07940_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13567_ (.A1(net3353),
    .A2(_07940_),
    .B(net3352),
    .ZN(_07941_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13568_ (.A1(net480),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .Z(_07942_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13569_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S0(net3635),
    .S1(net3596),
    .Z(_07943_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13570_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .S0(net3635),
    .S1(net3596),
    .Z(_07944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13571_ (.I0(_07943_),
    .I1(_07944_),
    .S(net3459),
    .Z(_07945_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13572_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S0(net3635),
    .S1(net3596),
    .Z(_07946_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13573_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .S0(net3635),
    .S1(net3596),
    .Z(_07947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13574_ (.I0(_07946_),
    .I1(_07947_),
    .S(net3459),
    .Z(_07948_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13575_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .S(net480),
    .Z(_07949_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13576_ (.A1(net3459),
    .A2(_07949_),
    .Z(_07950_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13577_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S0(net480),
    .S1(net3581),
    .Z(_07951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13578_ (.I0(_07950_),
    .I1(_07951_),
    .S(net3596),
    .Z(_07952_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13579_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S0(net480),
    .S1(net3596),
    .Z(_07953_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13580_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .S0(net480),
    .S1(net3596),
    .Z(_07954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13581_ (.I0(_07953_),
    .I1(_07954_),
    .S(net3459),
    .Z(_07955_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13582_ (.I0(_07945_),
    .I1(_07948_),
    .I2(_07952_),
    .I3(_07955_),
    .S0(net3579),
    .S1(_06290_),
    .Z(_07956_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13583_ (.A1(net3408),
    .A2(_07942_),
    .B(_07956_),
    .ZN(_07957_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13584_ (.A1(_06310_),
    .A2(net3343),
    .ZN(_07958_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13585_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(_06313_),
    .Z(_07959_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13586_ (.A1(_07941_),
    .A2(_07958_),
    .A3(_07959_),
    .Z(_11598_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _13587_ (.I(_11598_[0]),
    .ZN(_11594_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13588_ (.I(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .ZN(_07960_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _13589_ (.A1(_07960_),
    .A2(net3375),
    .A3(_07029_),
    .B1(_11594_[0]),
    .B2(net3373),
    .ZN(_11115_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13590_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S0(net3571),
    .S1(net3542),
    .Z(_07961_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13591_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .S0(net3571),
    .S1(net3542),
    .Z(_07962_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13592_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S0(net3571),
    .S1(net3542),
    .Z(_07963_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13593_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .S0(net3569),
    .S1(net3541),
    .Z(_07964_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13594_ (.I0(_07961_),
    .I1(_07962_),
    .I2(_07963_),
    .I3(_07964_),
    .S0(net3429),
    .S1(net3492),
    .Z(_07965_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13595_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S0(net3569),
    .S1(net3541),
    .Z(_07966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13596_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .S(net3541),
    .Z(_07967_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13597_ (.A1(net3541),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .Z(_07968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13598_ (.I0(_07967_),
    .I1(_07968_),
    .S(net3446),
    .Z(_07969_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13599_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S0(net3569),
    .S1(net3542),
    .Z(_07970_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13600_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .S0(net3569),
    .S1(net3542),
    .Z(_07971_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13601_ (.I0(_07966_),
    .I1(_07969_),
    .I2(_07970_),
    .I3(_07971_),
    .S0(net3429),
    .S1(net3492),
    .Z(_07972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13602_ (.I0(_07965_),
    .I1(_07972_),
    .S(net3421),
    .Z(_07973_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3270 (.I(_08553_),
    .Z(net3270));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13604_ (.A1(net3486),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_07975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13605_ (.I(_07975_),
    .ZN(_07976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _13606_ (.A1(net3380),
    .A2(_07973_),
    .B1(_07976_),
    .B2(net3379),
    .ZN(_11593_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13607_ (.I(_11593_[0]),
    .ZN(_11597_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _13608_ (.I(_11117_[0]),
    .ZN(_07977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13609_ (.A1(_11109_[0]),
    .A2(_11113_[0]),
    .ZN(_07978_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13610_ (.A1(_11113_[0]),
    .A2(_11108_[0]),
    .B(_11112_[0]),
    .ZN(_07979_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13611_ (.A1(_07888_),
    .A2(_07978_),
    .B(_07979_),
    .ZN(_07980_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _13612_ (.A1(_07977_),
    .A2(_07980_),
    .ZN(net166));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13613_ (.I(_11113_[0]),
    .ZN(_07981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13614_ (.A1(_11109_[0]),
    .A2(_07880_),
    .ZN(_07982_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13615_ (.A1(_07898_),
    .A2(_07889_),
    .B(_07882_),
    .ZN(_07983_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13616_ (.A1(_11109_[0]),
    .A2(_07983_),
    .B(_11108_[0]),
    .ZN(_07984_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13617_ (.A1(_07795_),
    .A2(_07797_),
    .A3(_07982_),
    .B(_07984_),
    .ZN(_07985_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _13618_ (.A1(_07985_),
    .A2(_07981_),
    .ZN(net165));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13619_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[26] ),
    .ZN(_07986_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13620_ (.A1(net3353),
    .A2(_07986_),
    .B(net3352),
    .ZN(_07987_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13621_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S0(net3635),
    .S1(net3596),
    .Z(_07988_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13622_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S0(net480),
    .S1(net3596),
    .Z(_07989_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13623_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S0(net3635),
    .S1(net3596),
    .Z(_07990_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13624_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S0(net480),
    .S1(net3596),
    .Z(_07991_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13625_ (.I0(_07988_),
    .I1(_07989_),
    .I2(_07990_),
    .I3(_07991_),
    .S0(net3459),
    .S1(net3579),
    .Z(_07992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13626_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .S(net480),
    .Z(_07993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13627_ (.A1(net480),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .Z(_07994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13628_ (.I0(_07993_),
    .I1(_07994_),
    .S(net3459),
    .Z(_07995_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13629_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .S0(net3642),
    .S1(net3581),
    .Z(_07996_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13630_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S0(net480),
    .S1(net3581),
    .Z(_07997_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13631_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S0(net454),
    .S1(net3581),
    .Z(_07998_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13632_ (.I0(_07995_),
    .I1(_07996_),
    .I2(_07997_),
    .I3(_07998_),
    .S0(net3579),
    .S1(net3596),
    .Z(_07999_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13633_ (.A1(net3577),
    .A2(_07999_),
    .Z(_08000_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13634_ (.A1(_06290_),
    .A2(_07992_),
    .B(_08000_),
    .ZN(_08001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13635_ (.A1(_06310_),
    .A2(net3342),
    .ZN(_08002_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13636_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(_06313_),
    .Z(_08003_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13637_ (.A1(_07987_),
    .A2(_08002_),
    .A3(_08003_),
    .Z(_11606_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _13638_ (.I(_11606_[0]),
    .ZN(_11602_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13639_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(_07017_),
    .Z(_08004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13640_ (.I0(_11606_[0]),
    .I1(_08004_),
    .S(net3371),
    .Z(_11119_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13641_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S0(net3566),
    .S1(net3535),
    .Z(_08005_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13642_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S0(net3566),
    .S1(net3535),
    .Z(_08006_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13643_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S0(net3566),
    .S1(net3535),
    .Z(_08007_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13644_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S0(net3566),
    .S1(net3535),
    .Z(_08008_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13645_ (.I0(_08005_),
    .I1(_08006_),
    .I2(_08007_),
    .I3(_08008_),
    .S0(net3427),
    .S1(net3492),
    .Z(_08009_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13646_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S0(net3566),
    .S1(net3535),
    .Z(_08010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13647_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .S(net3533),
    .Z(_08011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13648_ (.A1(net3533),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .Z(_08012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13649_ (.I0(_08011_),
    .I1(_08012_),
    .S(net3445),
    .Z(_08013_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13650_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S0(net3566),
    .S1(net3533),
    .Z(_08014_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13651_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S0(net3566),
    .S1(net3533),
    .Z(_08015_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13652_ (.I0(_08010_),
    .I1(_08013_),
    .I2(_08014_),
    .I3(_08015_),
    .S0(net3427),
    .S1(net3492),
    .Z(_08016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13653_ (.I0(_08009_),
    .I1(_08016_),
    .S(net3421),
    .Z(_08017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3533 (.I(net423),
    .Z(net3533));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13655_ (.A1(net3485),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_08019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13656_ (.I(_08019_),
    .ZN(_08020_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13657_ (.A1(net3380),
    .A2(_08017_),
    .B1(_08020_),
    .B2(net3379),
    .ZN(_11601_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13658_ (.I(_11601_[0]),
    .ZN(_11605_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13659_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[27] ),
    .ZN(_08021_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13660_ (.A1(net3353),
    .A2(_08021_),
    .B(net3352),
    .ZN(_08022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13661_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .S(net3637),
    .Z(_08023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13662_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S(net3637),
    .Z(_08024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13663_ (.A1(net3637),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .Z(_08025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13664_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net3637),
    .Z(_08026_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13665_ (.I0(_08023_),
    .I1(_08024_),
    .I2(_08025_),
    .I3(_08026_),
    .S0(net3596),
    .S1(net3459),
    .Z(_08027_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13666_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .S0(net3637),
    .S1(net3581),
    .Z(_08028_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13667_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S0(net3636),
    .S1(net3581),
    .Z(_08029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13668_ (.I0(_08028_),
    .I1(_08029_),
    .S(net3596),
    .Z(_08030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13669_ (.I0(_08027_),
    .I1(_08030_),
    .S(net3579),
    .Z(_08031_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13670_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08032_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13671_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08033_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13672_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08034_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13673_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08035_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13674_ (.I0(_08032_),
    .I1(_08033_),
    .I2(_08034_),
    .I3(_08035_),
    .S0(net3459),
    .S1(net3579),
    .Z(_08036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13675_ (.A1(net3577),
    .A2(_08036_),
    .Z(_08037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13676_ (.A1(_06290_),
    .A2(_08031_),
    .B(_08037_),
    .ZN(_08038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13677_ (.A1(_06310_),
    .A2(net3357),
    .ZN(_08039_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13678_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(_06313_),
    .Z(_08040_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13679_ (.A1(_08022_),
    .A2(_08039_),
    .A3(_08040_),
    .Z(_11614_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _13680_ (.I(_11614_[0]),
    .ZN(_11610_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _13681_ (.I(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .ZN(_08041_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _13682_ (.A1(_08041_),
    .A2(net3375),
    .A3(_07029_),
    .B1(_11610_[0]),
    .B2(net3373),
    .ZN(_11123_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3261 (.I(_08576_),
    .Z(net3261));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13684_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S0(net3566),
    .S1(net3536),
    .Z(_08043_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13685_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S0(net3566),
    .S1(net3536),
    .Z(_08044_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13686_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S0(net3566),
    .S1(net3536),
    .Z(_08045_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13687_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .S0(net3566),
    .S1(net3536),
    .Z(_08046_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13688_ (.I0(_08043_),
    .I1(_08044_),
    .I2(_08045_),
    .I3(_08046_),
    .S0(net3427),
    .S1(net3492),
    .Z(_08047_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13689_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S0(net3566),
    .S1(net3534),
    .Z(_08048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13690_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net3534),
    .Z(_08049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13691_ (.A1(net3534),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .Z(_08050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13692_ (.I0(_08049_),
    .I1(_08050_),
    .S(net3445),
    .Z(_08051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13693_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S0(net3566),
    .S1(net3535),
    .Z(_08052_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13694_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .S0(net3566),
    .S1(net3535),
    .Z(_08053_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13695_ (.I0(_08048_),
    .I1(_08051_),
    .I2(_08052_),
    .I3(_08053_),
    .S0(net3427),
    .S1(net3492),
    .Z(_08054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13696_ (.I0(_08047_),
    .I1(_08054_),
    .S(net3421),
    .Z(_08055_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13698_ (.A1(net3484),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_08057_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13699_ (.I(_08057_),
    .ZN(_08058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _13700_ (.A1(net3380),
    .A2(net419),
    .B1(_08058_),
    .B2(net3379),
    .ZN(_11609_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13701_ (.I(_11609_[0]),
    .ZN(_11613_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13702_ (.A1(_07977_),
    .A2(_07978_),
    .ZN(_08059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13703_ (.A1(_07880_),
    .A2(_08059_),
    .Z(_08060_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13704_ (.A1(_11093_[0]),
    .A2(_08060_),
    .ZN(_08061_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13705_ (.A1(_07977_),
    .A2(_07979_),
    .ZN(_08062_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13706_ (.A1(_11116_[0]),
    .A2(_11120_[0]),
    .A3(_08062_),
    .Z(_08063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13707_ (.A1(_07887_),
    .A2(_08059_),
    .B(_08063_),
    .ZN(_08064_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13708_ (.A1(_07685_),
    .A2(_08061_),
    .B(_08064_),
    .ZN(_08065_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13709_ (.A1(_11121_[0]),
    .A2(_11120_[0]),
    .Z(_08066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13710_ (.A1(_08066_),
    .A2(net345),
    .ZN(_08067_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _13711_ (.A1(_11125_[0]),
    .A2(_08067_),
    .ZN(net168));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13712_ (.I(_08059_),
    .ZN(_08068_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13713_ (.A1(_11109_[0]),
    .A2(_11104_[0]),
    .B(_11108_[0]),
    .ZN(_08069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13714_ (.I(_11112_[0]),
    .ZN(_08070_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13715_ (.A1(_07981_),
    .A2(_08069_),
    .B(_08070_),
    .ZN(_08071_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13716_ (.A1(_11117_[0]),
    .A2(_08071_),
    .B(_11116_[0]),
    .ZN(_08072_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13717_ (.A1(_07900_),
    .A2(_07898_),
    .A3(_08068_),
    .B(_08072_),
    .ZN(_08073_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13718_ (.A1(_11105_[0]),
    .A2(_07398_),
    .A3(_07895_),
    .A4(_08059_),
    .Z(_08074_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13719_ (.A1(_07304_),
    .A2(_07306_),
    .A3(_08074_),
    .Z(_08075_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13720_ (.A1(net395),
    .A2(_08075_),
    .B(_11121_[0]),
    .ZN(_08076_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13721_ (.A1(_08075_),
    .A2(net395),
    .A3(_11121_[0]),
    .Z(_08077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13722_ (.A1(_08077_),
    .A2(_08076_),
    .ZN(_08078_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _13723_ (.I(net347),
    .ZN(net167));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13724_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[28] ),
    .ZN(_08079_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13725_ (.A1(net3353),
    .A2(_08079_),
    .B(net3352),
    .ZN(_08080_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13726_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S0(net3639),
    .S1(net3596),
    .Z(_08081_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13727_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08082_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13728_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08083_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13729_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08084_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13730_ (.I0(_08081_),
    .I1(_08082_),
    .I2(_08083_),
    .I3(_08084_),
    .S0(net3459),
    .S1(net3579),
    .Z(_08085_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13731_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S0(net3639),
    .S1(net3596),
    .Z(_08086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13732_ (.A1(net3639),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .Z(_08087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13733_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .S(net3639),
    .Z(_08088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13734_ (.I0(_08087_),
    .I1(_08088_),
    .S(net3596),
    .Z(_08089_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13735_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S0(net3639),
    .S1(net3596),
    .Z(_08090_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13736_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .S0(net3639),
    .S1(net3596),
    .Z(_08091_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13737_ (.I0(_08086_),
    .I1(_08089_),
    .I2(_08090_),
    .I3(_08091_),
    .S0(net3459),
    .S1(net3579),
    .Z(_08092_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13738_ (.A1(net3577),
    .A2(_08092_),
    .Z(_08093_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13739_ (.A1(_06290_),
    .A2(_08085_),
    .B(_08093_),
    .ZN(_08094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13740_ (.A1(_06310_),
    .A2(net3341),
    .ZN(_08095_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13741_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(_06313_),
    .Z(_08096_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13742_ (.A1(_08080_),
    .A2(_08095_),
    .A3(_08096_),
    .Z(_11622_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _13743_ (.I(_11622_[0]),
    .ZN(_11618_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13744_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(_07017_),
    .Z(_08097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13745_ (.I0(_11622_[0]),
    .I1(_08097_),
    .S(net3371),
    .Z(_11127_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13746_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S0(net3569),
    .S1(net3538),
    .Z(_08098_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13747_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .S0(net3569),
    .S1(net3537),
    .Z(_08099_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13748_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S0(net3569),
    .S1(net3537),
    .Z(_08100_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13749_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .S0(net3569),
    .S1(net3537),
    .Z(_08101_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13750_ (.I0(_08098_),
    .I1(_08099_),
    .I2(_08100_),
    .I3(_08101_),
    .S0(net3427),
    .S1(net3492),
    .Z(_08102_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13751_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S0(net3569),
    .S1(net3538),
    .Z(_08103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13752_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .S(net3534),
    .Z(_08104_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13753_ (.A1(net3534),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .Z(_08105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13754_ (.I0(_08104_),
    .I1(_08105_),
    .S(net3446),
    .Z(_08106_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13755_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S0(net3569),
    .S1(net3538),
    .Z(_08107_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13756_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .S0(net3569),
    .S1(net3538),
    .Z(_08108_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13757_ (.I0(_08103_),
    .I1(_08106_),
    .I2(_08107_),
    .I3(_08108_),
    .S0(net3427),
    .S1(net3492),
    .Z(_08109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13758_ (.I0(_08102_),
    .I1(_08109_),
    .S(net3421),
    .Z(_08110_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13760_ (.A1(net3479),
    .A2(_07736_),
    .Z(_08112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13761_ (.I0(net3483),
    .I1(_08112_),
    .S(_06396_),
    .Z(_08113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _13762_ (.A1(net3380),
    .A2(net530),
    .B1(_08113_),
    .B2(net3379),
    .ZN(_11617_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13763_ (.I(_11617_[0]),
    .ZN(_11621_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13764_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[29] ),
    .ZN(_08114_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13765_ (.A1(net3353),
    .A2(_08114_),
    .B(net3352),
    .ZN(_08115_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13766_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08116_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13767_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08117_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13768_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08118_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13769_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08119_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13770_ (.I0(_08116_),
    .I1(_08117_),
    .I2(_08118_),
    .I3(_08119_),
    .S0(net3459),
    .S1(net3579),
    .Z(_08120_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13771_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S0(net3638),
    .S1(net3596),
    .Z(_08121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13772_ (.A1(net3638),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .Z(_08122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13773_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net3634),
    .Z(_08123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13774_ (.I0(_08122_),
    .I1(_08123_),
    .S(net3596),
    .Z(_08124_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13775_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S0(net3638),
    .S1(net3596),
    .Z(_08125_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13776_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .S0(net3636),
    .S1(net3596),
    .Z(_08126_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13777_ (.I0(_08121_),
    .I1(_08124_),
    .I2(_08125_),
    .I3(_08126_),
    .S0(net3459),
    .S1(net3579),
    .Z(_08127_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13778_ (.A1(net3577),
    .A2(_08127_),
    .Z(_08128_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13779_ (.A1(_06290_),
    .A2(_08120_),
    .B(_08128_),
    .ZN(_08129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13780_ (.A1(_06310_),
    .A2(net3340),
    .ZN(_08130_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13781_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(_06313_),
    .Z(_08131_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13782_ (.A1(_08115_),
    .A2(_08130_),
    .A3(_08131_),
    .Z(_11630_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _13783_ (.I(_11630_[0]),
    .ZN(_11626_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13784_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(_07017_),
    .Z(_08132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13785_ (.I0(_11630_[0]),
    .I1(_08132_),
    .S(net3371),
    .Z(_11131_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13786_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S0(net3566),
    .S1(net3537),
    .Z(_08133_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13787_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .S0(net3566),
    .S1(net3537),
    .Z(_08134_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13788_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S0(net3566),
    .S1(net3537),
    .Z(_08135_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13789_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S0(net3566),
    .S1(net3537),
    .Z(_08136_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13790_ (.I0(_08133_),
    .I1(_08134_),
    .I2(_08135_),
    .I3(_08136_),
    .S0(net3427),
    .S1(net3492),
    .Z(_08137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13791_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S0(net3566),
    .S1(net3537),
    .Z(_08138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13792_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net3534),
    .Z(_08139_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13793_ (.A1(net3534),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .Z(_08140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13794_ (.I0(_08139_),
    .I1(_08140_),
    .S(net3446),
    .Z(_08141_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13795_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S0(net3566),
    .S1(net3537),
    .Z(_08142_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13796_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .S0(net3566),
    .S1(net3537),
    .Z(_08143_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13797_ (.I0(_08138_),
    .I1(_08141_),
    .I2(_08142_),
    .I3(_08143_),
    .S0(net3427),
    .S1(net3492),
    .Z(_08144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13798_ (.I0(_08137_),
    .I1(_08144_),
    .S(net3421),
    .Z(_08145_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13800_ (.I0(net3482),
    .I1(_08112_),
    .S(_06396_),
    .Z(_08147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _13801_ (.A1(net3380),
    .A2(_08145_),
    .B1(_08147_),
    .B2(net3379),
    .ZN(_11625_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13802_ (.I(_11625_[0]),
    .ZN(_11629_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13803_ (.A1(_11125_[0]),
    .A2(_11129_[0]),
    .A3(_08066_),
    .ZN(_08148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13804_ (.I(_08148_),
    .ZN(_08149_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13805_ (.A1(_08065_),
    .A2(_08149_),
    .Z(_08150_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13806_ (.A1(_11129_[0]),
    .A2(_11124_[0]),
    .Z(_08151_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13807_ (.A1(_08150_),
    .A2(_11128_[0]),
    .A3(_08151_),
    .Z(_08152_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _13808_ (.A1(_11133_[0]),
    .A2(_08152_),
    .Z(net170));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13809_ (.A1(_11121_[0]),
    .A2(_11125_[0]),
    .A3(_08060_),
    .ZN(_08153_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _13810_ (.A1(_07795_),
    .A2(_11129_[0]),
    .A3(_07797_),
    .A4(_08153_),
    .Z(_08154_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13811_ (.A1(_07981_),
    .A2(_07984_),
    .B(_08070_),
    .ZN(_08155_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13812_ (.A1(_11117_[0]),
    .A2(_08155_),
    .B(_11116_[0]),
    .ZN(_08156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13813_ (.A1(_11121_[0]),
    .A2(_11125_[0]),
    .ZN(_08157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13814_ (.A1(_11125_[0]),
    .A2(_11120_[0]),
    .B(_11124_[0]),
    .ZN(_08158_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13815_ (.A1(_08156_),
    .A2(_08157_),
    .B(_08158_),
    .ZN(_08159_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _13816_ (.A1(_07795_),
    .A2(_07797_),
    .A3(_08153_),
    .B1(_08159_),
    .B2(_11129_[0]),
    .ZN(_08160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13817_ (.A1(_11129_[0]),
    .A2(_08159_),
    .Z(_08161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13818_ (.A1(net486),
    .A2(net387),
    .B(_08161_),
    .ZN(net169));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13819_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(net3394),
    .B(\cs_registers_i.pc_id_i[30] ),
    .ZN(_08162_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13820_ (.A1(net3353),
    .A2(_08162_),
    .B(net3352),
    .ZN(_08163_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13821_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S0(net3641),
    .S1(net3596),
    .Z(_08164_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13822_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .S0(net3641),
    .S1(net3596),
    .Z(_08165_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13823_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S0(net3641),
    .S1(net3596),
    .Z(_08166_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13824_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .S0(net3641),
    .S1(net3596),
    .Z(_08167_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _13825_ (.I0(_08164_),
    .I1(_08165_),
    .I2(_08166_),
    .I3(_08167_),
    .S0(net3459),
    .S1(net3579),
    .Z(_08168_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13826_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S0(net3639),
    .S1(net3596),
    .Z(_08169_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13827_ (.A1(net480),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .Z(_08170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13828_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net3634),
    .Z(_08171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13829_ (.I0(_08170_),
    .I1(_08171_),
    .S(net3596),
    .Z(_08172_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13830_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S0(net3639),
    .S1(net3596),
    .Z(_08173_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13831_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S0(net3639),
    .S1(net3596),
    .Z(_08174_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13832_ (.I0(_08169_),
    .I1(_08172_),
    .I2(_08173_),
    .I3(_08174_),
    .S0(net3459),
    .S1(net3579),
    .Z(_08175_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13833_ (.A1(net3577),
    .A2(_08175_),
    .Z(_08176_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13834_ (.A1(_06290_),
    .A2(_08168_),
    .B(_08176_),
    .ZN(_08177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13835_ (.A1(_06310_),
    .A2(net3339),
    .ZN(_08178_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13836_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(_06313_),
    .Z(_08179_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13837_ (.A1(_08163_),
    .A2(_08178_),
    .A3(_08179_),
    .Z(_11638_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _13838_ (.I(_11638_[0]),
    .ZN(_11634_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13839_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(_07017_),
    .Z(_08180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13840_ (.I0(_11638_[0]),
    .I1(_08180_),
    .S(net3371),
    .Z(_11135_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13841_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S0(net3569),
    .S1(net3545),
    .Z(_08181_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13842_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .S0(net3569),
    .S1(net3545),
    .Z(_08182_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13843_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S0(net3569),
    .S1(net3545),
    .Z(_08183_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13844_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .S0(net3569),
    .S1(net3545),
    .Z(_08184_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13845_ (.I0(_08181_),
    .I1(_08182_),
    .I2(_08183_),
    .I3(_08184_),
    .S0(net3428),
    .S1(net3492),
    .Z(_08185_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13846_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S0(net3572),
    .S1(net3539),
    .Z(_08186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13847_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net3539),
    .Z(_08187_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13848_ (.A1(net3539),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .Z(_08188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13849_ (.I0(_08187_),
    .I1(_08188_),
    .S(net3447),
    .Z(_08189_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13850_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S0(net3572),
    .S1(net3539),
    .Z(_08190_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13851_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S0(net3572),
    .S1(net3539),
    .Z(_08191_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13852_ (.I0(_08186_),
    .I1(_08189_),
    .I2(_08190_),
    .I3(_08191_),
    .S0(net3428),
    .S1(net3492),
    .Z(_08192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13853_ (.I0(_08185_),
    .I1(_08192_),
    .S(net3422),
    .Z(_08193_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3616 (.I(net449),
    .Z(net3616));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13855_ (.A1(net3480),
    .A2(_07734_),
    .B(_07737_),
    .ZN(_08195_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13856_ (.I(_08195_),
    .ZN(_08196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13857_ (.A1(net3380),
    .A2(_08193_),
    .B1(_08196_),
    .B2(net3379),
    .ZN(_11633_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13858_ (.I(_11633_[0]),
    .ZN(_11637_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13859_ (.A1(_06217_),
    .A2(_06223_),
    .Z(_08197_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13860_ (.A1(_06884_),
    .A2(_08197_),
    .A3(_06228_),
    .B(_06354_),
    .ZN(_08198_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13861_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(net3394),
    .Z(_08199_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13862_ (.A1(\cs_registers_i.pc_id_i[31] ),
    .A2(_08199_),
    .Z(_08200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13863_ (.A1(_08198_),
    .A2(_08200_),
    .B(_07625_),
    .ZN(_08201_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13864_ (.A1(_06208_),
    .A2(_06256_),
    .A3(_06236_),
    .ZN(_08202_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13865_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_08203_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13866_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .S0(net3622),
    .S1(net3597),
    .Z(_08204_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13867_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S0(net3623),
    .S1(net3598),
    .Z(_08205_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13868_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .S0(net3623),
    .S1(net3598),
    .Z(_08206_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13869_ (.I0(_08203_),
    .I1(_08204_),
    .I2(_08205_),
    .I3(_08206_),
    .S0(net3454),
    .S1(_07416_),
    .Z(_08207_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13870_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S0(net3623),
    .S1(net3598),
    .Z(_08208_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13871_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .S0(net3623),
    .S1(net3598),
    .Z(_08209_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13872_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S0(net3623),
    .S1(net3598),
    .Z(_08210_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13873_ (.A1(net3623),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .Z(_08211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13874_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .S(net3623),
    .Z(_08212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13875_ (.I0(_08211_),
    .I1(_08212_),
    .S(net3598),
    .Z(_08213_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13876_ (.I0(_08208_),
    .I1(_08209_),
    .I2(_08210_),
    .I3(_08213_),
    .S0(net3454),
    .S1(_07416_),
    .Z(_08214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13877_ (.I0(_08207_),
    .I1(_08214_),
    .S(_06290_),
    .Z(_08215_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _13878_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(_06313_),
    .B1(_08202_),
    .B2(net3356),
    .ZN(_08216_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13879_ (.A1(_08201_),
    .A2(_08216_),
    .ZN(_11143_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _13880_ (.I(_11143_[0]),
    .ZN(_11139_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13881_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .S0(net3568),
    .S1(net3548),
    .Z(_08217_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13882_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .S0(net3568),
    .S1(net3548),
    .Z(_08218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13883_ (.I0(_08217_),
    .I1(_08218_),
    .S(net3433),
    .Z(_08219_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13884_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S0(net3547),
    .S1(net3510),
    .Z(_08220_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13885_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .S0(net3547),
    .S1(net3510),
    .Z(_08221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13886_ (.I0(_08220_),
    .I1(_08221_),
    .S(net3448),
    .Z(_08222_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13887_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S0(net3574),
    .S1(net3542),
    .Z(_08223_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13888_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .S0(net3569),
    .S1(net3542),
    .Z(_08224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13889_ (.I0(_08223_),
    .I1(_08224_),
    .S(net3433),
    .Z(_08225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13890_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .S(net3547),
    .Z(_08226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13891_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S(net3542),
    .Z(_08227_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13892_ (.A1(net3542),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .Z(_08228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13893_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .S(net3542),
    .Z(_08229_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13894_ (.I0(_08226_),
    .I1(_08227_),
    .I2(_08228_),
    .I3(_08229_),
    .S0(net3568),
    .S1(net3433),
    .Z(_08230_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _13895_ (.I0(_08219_),
    .I1(_08222_),
    .I2(_08225_),
    .I3(_08230_),
    .S0(net3425),
    .S1(net3421),
    .Z(_08231_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3255 (.I(_08616_),
    .Z(net3255));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13897_ (.I0(_08112_),
    .I1(net431),
    .S(net3380),
    .Z(_11142_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13898_ (.I(_11142_[0]),
    .ZN(_11138_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _13899_ (.A1(_06777_),
    .A2(net327),
    .A3(_07011_),
    .ZN(_08233_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13900_ (.A1(net305),
    .A2(_08233_),
    .A3(_11142_[0]),
    .Z(_08234_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _13901_ (.I(net3356),
    .ZN(_08235_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13902_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net432),
    .ZN(_08236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13903_ (.A1(net3655),
    .A2(_08235_),
    .B(_08236_),
    .ZN(_08237_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _13904_ (.A1(net305),
    .A2(_11142_[0]),
    .B1(_08237_),
    .B2(net3374),
    .ZN(_08238_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13905_ (.A1(net3370),
    .A2(_08201_),
    .A3(_08216_),
    .Z(_08239_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _13906_ (.I(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .ZN(_08240_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13907_ (.A1(_08240_),
    .A2(_08233_),
    .A3(_07029_),
    .Z(_08241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13908_ (.A1(_08239_),
    .A2(_08241_),
    .Z(_08242_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13909_ (.A1(_08234_),
    .A2(_08238_),
    .B(_08242_),
    .ZN(_08243_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13910_ (.A1(_08234_),
    .A2(_08238_),
    .A3(_08242_),
    .Z(_08244_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13911_ (.A1(_11128_[0]),
    .A2(_08151_),
    .ZN(_08245_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13912_ (.A1(_11136_[0]),
    .A2(_11132_[0]),
    .ZN(_08246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13913_ (.A1(_08245_),
    .A2(_08246_),
    .ZN(_08247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13914_ (.A1(_08065_),
    .A2(_08149_),
    .B(_08247_),
    .ZN(_08248_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13915_ (.A1(_11133_[0]),
    .A2(_11132_[0]),
    .Z(_08249_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13916_ (.A1(_11137_[0]),
    .A2(_08249_),
    .B(_11136_[0]),
    .ZN(_08250_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13917_ (.A1(_08248_),
    .A2(_08250_),
    .ZN(_08251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13918_ (.A1(_08243_),
    .A2(_08244_),
    .B(_08251_),
    .ZN(_08252_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13919_ (.A1(_08251_),
    .A2(_08243_),
    .A3(_08244_),
    .Z(_08253_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13920_ (.A1(_08252_),
    .A2(_08253_),
    .ZN(_08254_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _13921_ (.I(net3094),
    .ZN(net173));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13922_ (.A1(_11133_[0]),
    .A2(_11132_[0]),
    .ZN(_08255_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13923_ (.I(_11129_[0]),
    .ZN(_08256_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13924_ (.A1(_08256_),
    .A2(_08158_),
    .ZN(_08257_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13925_ (.A1(_11128_[0]),
    .A2(_11132_[0]),
    .A3(_08257_),
    .Z(_08258_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _13926_ (.A1(_08258_),
    .A2(_08075_),
    .A3(_08073_),
    .ZN(_08259_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13927_ (.A1(_08256_),
    .A2(_08157_),
    .ZN(_08260_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13928_ (.A1(_08260_),
    .A2(_08258_),
    .ZN(_08261_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13929_ (.A1(_08255_),
    .A2(_08259_),
    .A3(_08261_),
    .B(_11137_[0]),
    .ZN(_08262_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _13930_ (.A1(_08259_),
    .A2(_08255_),
    .A3(_11137_[0]),
    .A4(_08261_),
    .Z(_08263_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13931_ (.A1(_08262_),
    .A2(_08263_),
    .ZN(net172));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3254 (.I(_08685_),
    .Z(net3254));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13933_ (.A1(_06206_),
    .A2(net3397),
    .ZN(_08265_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13934_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .A2(_06322_),
    .A3(_06331_),
    .ZN(_08266_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13935_ (.A1(_06316_),
    .A2(_06321_),
    .Z(_08267_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13936_ (.A1(_06224_),
    .A2(_06406_),
    .B1(_06328_),
    .B2(_06329_),
    .ZN(_08268_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13937_ (.A1(_06234_),
    .A2(_08267_),
    .A3(_08268_),
    .B(net3560),
    .ZN(_08269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13938_ (.A1(_06343_),
    .A2(_06352_),
    .ZN(_08270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13939_ (.A1(_08266_),
    .A2(_08269_),
    .B(_08270_),
    .ZN(_08271_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13940_ (.A1(_06355_),
    .A2(_06384_),
    .Z(_08272_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13941_ (.A1(_08271_),
    .A2(_08272_),
    .B(_06783_),
    .ZN(_08273_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13942_ (.A1(net485),
    .A2(_08273_),
    .ZN(_08274_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _13943_ (.A1(_06614_),
    .A2(_06594_),
    .A3(_06605_),
    .A4(_06586_),
    .ZN(_08275_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3445 (.I(_06334_),
    .Z(net3445));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13945_ (.A1(_08275_),
    .A2(_06653_),
    .Z(_08277_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13946_ (.A1(net3484),
    .A2(net3485),
    .Z(_08278_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13947_ (.A1(_06441_),
    .A2(_06533_),
    .A3(_08278_),
    .Z(_08279_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13948_ (.A1(_06355_),
    .A2(_08277_),
    .B(_08279_),
    .ZN(_08280_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13949_ (.A1(_06355_),
    .A2(net412),
    .A3(net407),
    .Z(_08281_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13950_ (.A1(_06621_),
    .A2(_06719_),
    .ZN(_08282_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13951_ (.A1(net3378),
    .A2(net3389),
    .Z(_08283_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13952_ (.A1(_06762_),
    .A2(_06621_),
    .B1(_08281_),
    .B2(_08282_),
    .C1(_08283_),
    .C2(_06441_),
    .ZN(_08284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13953_ (.A1(_06718_),
    .A2(_06782_),
    .ZN(_08285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13954_ (.A1(_06811_),
    .A2(_06843_),
    .B(_08284_),
    .C(_08285_),
    .ZN(_08286_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _13955_ (.A1(net3287),
    .A2(_11438_[0]),
    .A3(_08280_),
    .A4(_08286_),
    .Z(_08287_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13956_ (.A1(_11410_[0]),
    .A2(_08274_),
    .A3(_08287_),
    .Z(_08288_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13957_ (.A1(_06322_),
    .A2(_06331_),
    .ZN(_08289_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13958_ (.A1(net3560),
    .A2(_06338_),
    .A3(_06342_),
    .Z(_08290_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _13959_ (.I(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .ZN(_08291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13960_ (.A1(_06338_),
    .A2(_06342_),
    .B(_08291_),
    .ZN(_08292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13961_ (.I0(_08290_),
    .I1(_08292_),
    .S(_06465_),
    .Z(_08293_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13962_ (.A1(net3479),
    .A2(_06343_),
    .A3(_06465_),
    .Z(_08294_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13963_ (.A1(_08289_),
    .A2(_08293_),
    .B(_08294_),
    .C(_06355_),
    .ZN(_08295_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13964_ (.A1(net3380),
    .A2(net412),
    .A3(net407),
    .ZN(_08296_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13965_ (.A1(_06621_),
    .A2(_06719_),
    .Z(_08297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13966_ (.A1(_08296_),
    .A2(_08297_),
    .B(_11474_[0]),
    .ZN(_08298_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _13967_ (.A1(_08295_),
    .A2(_06842_),
    .B(_08298_),
    .C(_06783_),
    .ZN(_08299_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13968_ (.A1(_06773_),
    .A2(net3485),
    .Z(_08300_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13969_ (.A1(net341),
    .A2(_06615_),
    .ZN(_08301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13970_ (.A1(_06534_),
    .A2(_08300_),
    .B1(_08301_),
    .B2(_06355_),
    .ZN(_08302_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13971_ (.A1(_11450_[0]),
    .A2(_08302_),
    .Z(_08303_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13972_ (.A1(_06530_),
    .A2(_08299_),
    .A3(_08303_),
    .Z(_08304_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13973_ (.A1(_08295_),
    .A2(_06842_),
    .B(_06783_),
    .ZN(_08305_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13974_ (.A1(_06530_),
    .A2(_11454_[0]),
    .A3(_08302_),
    .Z(_08306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13975_ (.A1(net412),
    .A2(net407),
    .ZN(_08307_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13976_ (.A1(net3482),
    .A2(net3483),
    .Z(_08308_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _13977_ (.A1(net3480),
    .A2(_06441_),
    .A3(_06533_),
    .A4(_08308_),
    .ZN(_08309_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13978_ (.A1(_06441_),
    .A2(_08283_),
    .A3(_08307_),
    .B(_08309_),
    .ZN(_08310_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13979_ (.A1(_06399_),
    .A2(net329),
    .A3(_08310_),
    .ZN(_08311_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13980_ (.A1(_08305_),
    .A2(_08306_),
    .A3(_08311_),
    .Z(_08312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13981_ (.A1(_06743_),
    .A2(_06751_),
    .B(_08265_),
    .C(_06768_),
    .ZN(_08313_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _13982_ (.A1(_08295_),
    .A2(_06842_),
    .B(_08313_),
    .C(_08298_),
    .ZN(_08314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13983_ (.A1(_06396_),
    .A2(_06397_),
    .Z(_08315_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13984_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A2(_06465_),
    .A3(net3379),
    .A4(_08315_),
    .Z(_08316_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13985_ (.A1(_06528_),
    .A2(_06622_),
    .A3(_06654_),
    .Z(_08317_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _13986_ (.A1(_06527_),
    .A2(_08316_),
    .A3(_08302_),
    .A4(_08317_),
    .Z(_08318_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13987_ (.A1(_06388_),
    .A2(net485),
    .A3(_08314_),
    .A4(_08318_),
    .Z(_08319_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13988_ (.A1(_08304_),
    .A2(_08312_),
    .B1(_08319_),
    .B2(_11410_[0]),
    .ZN(_08320_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13989_ (.A1(_06620_),
    .A2(net3485),
    .ZN(_08321_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13990_ (.A1(net3486),
    .A2(_06441_),
    .A3(_06533_),
    .A4(_08321_),
    .Z(_08322_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13991_ (.A1(_06355_),
    .A2(net341),
    .A3(_06615_),
    .A4(_06653_),
    .Z(_08323_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13992_ (.A1(_08322_),
    .A2(_08323_),
    .Z(_08324_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13993_ (.A1(_11414_[0]),
    .A2(_08324_),
    .A3(_08286_),
    .Z(_08325_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13994_ (.A1(_08288_),
    .A2(_08320_),
    .A3(_08325_),
    .B(net3288),
    .ZN(_08326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13995_ (.A1(_11414_[0]),
    .A2(net3288),
    .ZN(_08327_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13996_ (.A1(_06388_),
    .A2(net485),
    .A3(_08327_),
    .B(_06783_),
    .ZN(_08328_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13997_ (.A1(net485),
    .A2(_08327_),
    .A3(_08273_),
    .B(_11438_[0]),
    .ZN(_08329_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13998_ (.A1(_06388_),
    .A2(net485),
    .A3(_11418_[0]),
    .B(_06783_),
    .ZN(_08330_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13999_ (.A1(net3287),
    .A2(_08280_),
    .A3(_08286_),
    .Z(_08331_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _14000_ (.A1(_11438_[0]),
    .A2(_08328_),
    .B1(_08329_),
    .B2(_08330_),
    .C(_08331_),
    .ZN(_08332_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _14001_ (.A1(net485),
    .A2(_08327_),
    .A3(_08273_),
    .Z(_08333_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14002_ (.A1(_06355_),
    .A2(_06615_),
    .A3(_06653_),
    .Z(_08334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14003_ (.A1(_06534_),
    .A2(_08321_),
    .B(_08334_),
    .ZN(_08335_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14004_ (.A1(_08285_),
    .A2(_08335_),
    .ZN(_08336_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14005_ (.A1(_08280_),
    .A2(_08336_),
    .Z(_08337_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14006_ (.A1(net341),
    .A2(_06841_),
    .Z(_08338_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _14007_ (.A1(net3486),
    .A2(_06534_),
    .B1(_08338_),
    .B2(_06355_),
    .ZN(_08339_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14008_ (.A1(_06783_),
    .A2(_06811_),
    .A3(_08298_),
    .A4(_08339_),
    .Z(_08340_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _14009_ (.A1(_06530_),
    .A2(_08333_),
    .B(_08337_),
    .C(_08340_),
    .ZN(_08341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14010_ (.A1(_06388_),
    .A2(net485),
    .B(_06530_),
    .C(_08327_),
    .ZN(_08342_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14011_ (.I(net341),
    .ZN(_08343_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14012_ (.A1(_06533_),
    .A2(_08278_),
    .Z(_08344_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _14013_ (.A1(_06441_),
    .A2(_08343_),
    .A3(_08277_),
    .B1(_08344_),
    .B2(_06535_),
    .ZN(_08345_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14014_ (.A1(_06530_),
    .A2(_08324_),
    .B(_08345_),
    .ZN(_08346_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _14015_ (.A1(_08299_),
    .A2(_08342_),
    .A3(_08346_),
    .Z(_08347_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14016_ (.A1(_11414_[0]),
    .A2(_11418_[0]),
    .ZN(_08348_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14017_ (.A1(_06353_),
    .A2(_06386_),
    .A3(_06783_),
    .Z(_08349_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14018_ (.A1(net263),
    .A2(_08348_),
    .A3(_08349_),
    .Z(_08350_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14019_ (.A1(_06530_),
    .A2(_06783_),
    .A3(_08310_),
    .Z(_08351_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14020_ (.A1(_06811_),
    .A2(_08280_),
    .A3(_08339_),
    .Z(_08352_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14021_ (.A1(_08351_),
    .A2(_08352_),
    .Z(_08353_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14022_ (.A1(_08295_),
    .A2(_06842_),
    .B(_08324_),
    .ZN(_08354_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14023_ (.A1(_06530_),
    .A2(_06783_),
    .A3(_08310_),
    .ZN(_08355_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _14024_ (.A1(_06783_),
    .A2(_08327_),
    .B(_08354_),
    .C(_08355_),
    .ZN(_08356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14025_ (.A1(_08350_),
    .A2(_08353_),
    .B(_08356_),
    .ZN(_08357_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14026_ (.A1(_08332_),
    .A2(_08341_),
    .A3(_08347_),
    .A4(_08357_),
    .Z(_08358_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14027_ (.A1(_11478_[0]),
    .A2(_11486_[0]),
    .Z(_08359_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _14028_ (.I(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .ZN(_08360_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14029_ (.I(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .ZN(_08361_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14030_ (.A1(_08361_),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Z(_08362_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _14031_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_08360_),
    .A3(_08362_),
    .ZN(_08363_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _14032_ (.A1(_06345_),
    .A2(\id_stage_i.controller_i.instr_fetch_err_i ),
    .A3(_08363_),
    .Z(_08364_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _14033_ (.A1(_11154_[0]),
    .A2(_08285_),
    .A3(_08359_),
    .A4(_08364_),
    .Z(_08365_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14034_ (.I(_08365_),
    .ZN(_08366_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14035_ (.I(_11161_[0]),
    .ZN(_08367_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14036_ (.A1(_11159_[0]),
    .A2(_08367_),
    .B(_11158_[0]),
    .ZN(_08368_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14037_ (.A1(_11159_[0]),
    .A2(_11162_[0]),
    .B(_08368_),
    .ZN(_08369_));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 _14038_ (.I(\cs_registers_i.debug_mode_i ),
    .ZN(_08370_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3498 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(net3498));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14040_ (.A1(_08370_),
    .A2(_08356_),
    .Z(_08372_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14041_ (.A1(_08369_),
    .A2(_08372_),
    .Z(_08373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14042_ (.A1(_08326_),
    .A2(_08358_),
    .B(_08366_),
    .C(_08373_),
    .ZN(_08374_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3669 (.I(net140),
    .Z(net3669));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14044_ (.A1(_08265_),
    .A2(_08374_),
    .B(_06782_),
    .ZN(_08376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14045_ (.A1(net3473),
    .A2(_08376_),
    .ZN(_08377_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _14046_ (.A1(net3485),
    .A2(net3479),
    .A3(_06731_),
    .ZN(_08378_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14047_ (.A1(net3473),
    .A2(_06206_),
    .A3(_06244_),
    .A4(_06720_),
    .Z(_08379_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14048_ (.A1(_08378_),
    .A2(_08379_),
    .Z(_08380_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14049_ (.A1(\cs_registers_i.priv_mode_id_o[1] ),
    .A2(\cs_registers_i.priv_mode_id_o[0] ),
    .Z(_08381_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14050_ (.A1(net3473),
    .A2(net3560),
    .A3(net3499),
    .A4(net3483),
    .Z(_08382_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14051_ (.A1(_06206_),
    .A2(_06244_),
    .A3(_06726_),
    .A4(_08382_),
    .Z(_08383_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14052_ (.A1(_06722_),
    .A2(_06724_),
    .ZN(_08384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14053_ (.A1(_08384_),
    .A2(_08379_),
    .Z(_08385_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14054_ (.A1(\cs_registers_i.csr_mstatus_tw_o ),
    .A2(_08383_),
    .B(_08385_),
    .ZN(_08386_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14055_ (.A1(_08381_),
    .A2(_08386_),
    .ZN(_08387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14056_ (.A1(_08370_),
    .A2(_08380_),
    .B(_08387_),
    .ZN(_08388_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _14057_ (.I(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .ZN(_08389_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14058_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_08361_),
    .A3(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Z(_08390_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14059_ (.A1(_08389_),
    .A2(_08390_),
    .Z(_08391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14060_ (.A1(_08377_),
    .A2(_08388_),
    .B(_08391_),
    .ZN(\id_stage_i.controller_i.illegal_insn_d ));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14061_ (.A1(_06206_),
    .A2(_06244_),
    .A3(_06726_),
    .A4(_06727_),
    .Z(_08392_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14062_ (.A1(net3473),
    .A2(_08392_),
    .Z(_08393_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _14063_ (.A1(\id_stage_i.controller_i.instr_fetch_err_i ),
    .A2(_08376_),
    .A3(_08393_),
    .B(net3473),
    .ZN(_08394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14064_ (.A1(_08388_),
    .A2(_08394_),
    .B(_08391_),
    .ZN(\id_stage_i.controller_i.exc_req_d ));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14065_ (.A1(_06232_),
    .A2(_06229_),
    .Z(_08395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14066_ (.A1(net59),
    .A2(_08395_),
    .ZN(_08396_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14067_ (.I(net25),
    .ZN(_08397_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14068_ (.I(\load_store_unit_i.lsu_err_q ),
    .ZN(_08398_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14069_ (.A1(_08397_),
    .A2(_08398_),
    .Z(_08399_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14070_ (.A1(_08396_),
    .A2(_08399_),
    .ZN(_08400_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14071_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_08400_),
    .Z(\id_stage_i.controller_i.store_err_i ));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _14072_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_08396_),
    .A3(_08399_),
    .ZN(\id_stage_i.controller_i.load_err_i ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _14073_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .ZN(_08401_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14074_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .ZN(_08402_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14075_ (.A1(_11177_[0]),
    .A2(_08402_),
    .Z(_08403_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _14076_ (.A1(_06345_),
    .A2(\id_stage_i.controller_i.instr_fetch_err_i ),
    .A3(_08363_),
    .ZN(_08404_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14077_ (.A1(_06782_),
    .A2(_08404_),
    .Z(_08405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14078_ (.A1(net3647),
    .A2(net3373),
    .Z(_08406_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14079_ (.A1(_08405_),
    .A2(_08406_),
    .Z(_08407_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3615 (.I(net415),
    .Z(net3615));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14081_ (.A1(_08403_),
    .A2(_08407_),
    .Z(_08409_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14082_ (.A1(_08401_),
    .A2(_08409_),
    .B(_07015_),
    .ZN(_08410_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14083_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A2(_08407_),
    .Z(_08411_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_44_clk_i_regs (.I(clknet_6_55__leaf_clk_i_regs),
    .Z(clknet_leaf_44_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14085_ (.A1(_08410_),
    .A2(_08411_),
    .Z(_00005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3253 (.I(net302),
    .Z(net3253));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14087_ (.I(net3655),
    .ZN(_08414_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3257 (.I(_08581_),
    .Z(net3257));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14089_ (.I(_07192_),
    .ZN(_08416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14090_ (.A1(_11017_[0]),
    .A2(net382),
    .ZN(_08417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14091_ (.A1(net305),
    .A2(_08233_),
    .B(_08417_),
    .ZN(_08418_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14092_ (.A1(_08416_),
    .A2(_08418_),
    .B(net308),
    .ZN(_08419_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _14093_ (.A1(net308),
    .A2(_08416_),
    .A3(_08418_),
    .Z(_08420_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14094_ (.A1(net292),
    .A2(_07187_),
    .Z(_08421_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14095_ (.A1(_07190_),
    .A2(net305),
    .A3(_08233_),
    .A4(net278),
    .Z(_08422_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14096_ (.A1(net292),
    .A2(_07187_),
    .ZN(_08423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14097_ (.I0(_11033_[0]),
    .I1(_08423_),
    .S(net272),
    .Z(_08424_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _14098_ (.A1(net260),
    .A2(_08421_),
    .B(_08422_),
    .C(_08424_),
    .ZN(net175));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _14099_ (.I(_11658_[0]),
    .ZN(_08425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14100_ (.A1(_07245_),
    .A2(net374),
    .B(_11028_[0]),
    .ZN(_08426_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14101_ (.A1(_07190_),
    .A2(_08426_),
    .B(_07196_),
    .ZN(_08427_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14102_ (.A1(net455),
    .A2(_08427_),
    .Z(net176));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14103_ (.A1(net475),
    .A2(_11021_[0]),
    .B(_11020_[0]),
    .ZN(_08428_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14104_ (.A1(net351),
    .A2(_08428_),
    .B(_07193_),
    .ZN(_08429_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _14105_ (.A1(_11029_[0]),
    .A2(_08429_),
    .Z(net174));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14106_ (.A1(_08425_),
    .A2(net178),
    .A3(net176),
    .A4(net174),
    .Z(_08430_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14107_ (.A1(net152),
    .A2(_08430_),
    .ZN(_08431_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _14108_ (.A1(_07202_),
    .A2(_07203_),
    .B(_07254_),
    .C(_08431_),
    .ZN(_08432_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14109_ (.A1(_08419_),
    .A2(_08420_),
    .B(net175),
    .C(_08432_),
    .ZN(_08433_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14110_ (.A1(_07261_),
    .A2(_07262_),
    .B(net154),
    .C(net157),
    .ZN(_08434_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _14111_ (.A1(_07308_),
    .A2(_07309_),
    .A3(net153),
    .A4(net156),
    .ZN(_08435_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14112_ (.I(net158),
    .ZN(_08436_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14113_ (.A1(_08436_),
    .A2(_07798_),
    .A3(_07799_),
    .Z(_08437_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14114_ (.A1(_08433_),
    .A2(_08434_),
    .A3(_08435_),
    .A4(_08437_),
    .Z(_08438_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14115_ (.A1(net155),
    .A2(net169),
    .ZN(_08439_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _14116_ (.A1(net160),
    .A2(net159),
    .A3(net163),
    .A4(net165),
    .ZN(_08440_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14117_ (.A1(_08076_),
    .A2(_08077_),
    .B(net162),
    .C(net164),
    .ZN(_08441_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14118_ (.A1(_08438_),
    .A2(_08439_),
    .A3(_08440_),
    .A4(_08441_),
    .Z(_08442_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _14119_ (.A1(net166),
    .A2(net367),
    .A3(net170),
    .ZN(_08443_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14120_ (.A1(net297),
    .A2(_08262_),
    .A3(net396),
    .A4(_08443_),
    .Z(_08444_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14121_ (.A1(_08442_),
    .A2(_08444_),
    .Z(_08445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14122_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_08407_),
    .ZN(_08446_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14123_ (.A1(_08414_),
    .A2(_08407_),
    .B1(_08445_),
    .B2(_08446_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3252 (.I(_11425_[0]),
    .Z(net3252));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3256 (.I(net3255),
    .Z(net3256));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14126_ (.A1(_06717_),
    .A2(_07020_),
    .ZN(_08449_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14127_ (.A1(net3659),
    .A2(net3338),
    .Z(_08450_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14128_ (.A1(net3657),
    .A2(_08450_),
    .Z(_08451_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _14129_ (.A1(net3658),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A3(_07017_),
    .Z(_08452_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14130_ (.A1(net320),
    .A2(_06243_),
    .ZN(_08453_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14131_ (.A1(net3373),
    .A2(_08453_),
    .Z(_08454_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14132_ (.A1(net3356),
    .A2(_08454_),
    .ZN(_08455_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14133_ (.A1(_06744_),
    .A2(_08406_),
    .Z(_08456_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14134_ (.A1(_08455_),
    .A2(_08456_),
    .B(net3658),
    .ZN(_08457_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14135_ (.A1(net3356),
    .A2(_08454_),
    .Z(_08458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14136_ (.A1(_06744_),
    .A2(_08406_),
    .ZN(_08459_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14137_ (.A1(net320),
    .A2(net3416),
    .B(_06344_),
    .ZN(_08460_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14138_ (.A1(net3373),
    .A2(_08460_),
    .Z(_08461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14139_ (.A1(net432),
    .A2(_08461_),
    .ZN(_08462_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _14140_ (.A1(_08458_),
    .A2(_08459_),
    .A3(_08462_),
    .Z(_08463_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3250 (.I(net3249),
    .Z(net3250));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14142_ (.A1(_08458_),
    .A2(_08462_),
    .ZN(_08465_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14143_ (.A1(_08463_),
    .A2(_08465_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .ZN(_08466_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14144_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_08452_),
    .B1(_08457_),
    .B2(_08466_),
    .ZN(_08467_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14145_ (.A1(net3647),
    .A2(_08467_),
    .ZN(_08468_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _14146_ (.A1(net3373),
    .A2(_08405_),
    .A3(_08468_),
    .ZN(_08469_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14147_ (.A1(_08406_),
    .A2(_08469_),
    .Z(_08470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14148_ (.I0(_08451_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .S(_08470_),
    .Z(_00000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14149_ (.A1(net3397),
    .A2(net3373),
    .Z(_08471_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14150_ (.A1(net3659),
    .A2(_08471_),
    .Z(_08472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14151_ (.I0(_08472_),
    .I1(net3657),
    .S(_08470_),
    .Z(_00001_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3497 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(net3497));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3247 (.I(_08517_),
    .Z(net3247));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3248 (.I(_08517_),
    .Z(net3248));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14155_ (.A1(net3654),
    .A2(_08401_),
    .A3(_08403_),
    .Z(_08476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14156_ (.I0(net3656),
    .I1(_08476_),
    .S(_08407_),
    .Z(_00002_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3244 (.I(_08529_),
    .Z(net3244));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14158_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_08445_),
    .ZN(_08478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14159_ (.A1(_07027_),
    .A2(_08478_),
    .ZN(_08479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14160_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .I1(_08479_),
    .S(_08407_),
    .Z(_00003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14161_ (.I(\cs_registers_i.pc_if_i[2] ),
    .ZN(_10997_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _14162_ (.I(_09748_[0]),
    .ZN(\alu_adder_result_ex[0] ));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14163_ (.A1(_08419_),
    .A2(_08420_),
    .Z(net171));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14164_ (.I0(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .S(net3338),
    .Z(_08480_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14165_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .Z(_08481_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3259 (.I(net3257),
    .Z(net3259));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14167_ (.A1(net3659),
    .A2(_08480_),
    .B1(net3407),
    .B2(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .ZN(_08483_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14168_ (.I(_08483_),
    .ZN(_11181_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14169_ (.I0(net334),
    .I1(_07544_),
    .S(_08481_),
    .Z(_08484_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3240 (.I(_08549_),
    .Z(net3240));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14171_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Z(_08486_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3241 (.I(net3240),
    .Z(net3241));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14173_ (.I0(_06916_),
    .I1(_07525_),
    .S(_08486_),
    .Z(_08488_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14174_ (.A1(net3337),
    .A2(net3334),
    .Z(_11182_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3655 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .Z(net3655));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3243 (.I(_08529_),
    .Z(net3243));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14177_ (.I0(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .S(net3338),
    .Z(_08491_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3238 (.I(_08556_),
    .Z(net3238));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14179_ (.A1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .A2(net3407),
    .B1(_08491_),
    .B2(net3659),
    .ZN(_09750_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14180_ (.I0(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .S(net3338),
    .Z(_08493_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14181_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(net3407),
    .B1(_08493_),
    .B2(net3659),
    .ZN(_09755_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3614 (.I(net333),
    .Z(net3614));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3236 (.I(net3235),
    .Z(net3236));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14184_ (.I0(_06457_),
    .I1(_07641_),
    .S(_08481_),
    .Z(_08496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14185_ (.A1(net3334),
    .A2(net529),
    .Z(_09760_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14186_ (.I0(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .S(net3338),
    .Z(_08497_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14187_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(net3407),
    .B1(_08497_),
    .B2(net3659),
    .ZN(_09766_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14188_ (.I0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .S(net3338),
    .Z(_08498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14189_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(net3407),
    .B1(_08498_),
    .B2(net3659),
    .ZN(_09774_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3496 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(net3496));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14191_ (.I0(_07060_),
    .I1(_07624_),
    .S(_08486_),
    .Z(_08500_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14192_ (.A1(net529),
    .A2(net3330),
    .Z(_09779_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14193_ (.I0(_06487_),
    .I1(_07676_),
    .S(_08481_),
    .Z(_08501_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3234 (.I(net3232),
    .Z(net3234));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14195_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .ZN(_08503_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3251 (.I(net3249),
    .Z(net3251));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14197_ (.I0(_06933_),
    .I1(_06926_),
    .S(_06290_),
    .Z(_08505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14198_ (.A1(_08505_),
    .A2(_08503_),
    .ZN(_08506_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14199_ (.A1(_07566_),
    .A2(_08503_),
    .B(_08506_),
    .ZN(_08507_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14200_ (.A1(net3328),
    .A2(net3285),
    .Z(_09778_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14201_ (.I0(net330),
    .I1(_07732_),
    .S(_08481_),
    .Z(_08508_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14202_ (.A1(net3334),
    .A2(net3325),
    .Z(_09777_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14203_ (.I0(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .S(net3338),
    .Z(_08509_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14204_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(net3407),
    .B1(_08509_),
    .B2(net3659),
    .ZN(_09792_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14205_ (.I0(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .S(net3338),
    .Z(_08510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14206_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(net3407),
    .B1(_08510_),
    .B2(net3659),
    .ZN(_09807_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14207_ (.I0(_07105_),
    .I1(_07711_),
    .S(_08486_),
    .Z(_08511_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14208_ (.A1(net529),
    .A2(net3321),
    .Z(_09812_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14209_ (.I(_07659_),
    .ZN(_08512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14210_ (.I0(_07087_),
    .I1(_08512_),
    .S(_08486_),
    .Z(_08513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14211_ (.A1(net3328),
    .A2(net3251),
    .Z(_09811_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14212_ (.A1(net3330),
    .A2(net3324),
    .Z(_09810_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14213_ (.I0(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .S(net3338),
    .Z(_08514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14214_ (.A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .A2(net3407),
    .B1(_08514_),
    .B2(net3659),
    .ZN(_09826_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _14215_ (.I(_07132_),
    .ZN(_08515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14216_ (.A1(_08515_),
    .A2(_08503_),
    .ZN(_08516_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14217_ (.A1(_07756_),
    .A2(_08503_),
    .B(_08516_),
    .ZN(_08517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14218_ (.A1(net529),
    .A2(net3247),
    .Z(_09833_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14219_ (.A1(net3328),
    .A2(net3321),
    .Z(_09832_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3227 (.I(_10255_[0]),
    .Z(net3227));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14221_ (.A1(net3324),
    .A2(net3251),
    .Z(_09831_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3648 (.I(net304),
    .Z(net3648));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14223_ (.I0(net341),
    .I1(_07776_),
    .S(_08481_),
    .Z(_08520_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3532 (.I(net3531),
    .Z(net3532));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14225_ (.A1(net3330),
    .A2(net3318),
    .ZN(_09841_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14226_ (.I0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .S(net3338),
    .Z(_08522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14227_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(net3407),
    .B1(_08522_),
    .B2(net3659),
    .ZN(_09863_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14228_ (.A1(net858),
    .A2(_08486_),
    .Z(_08523_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14229_ (.A1(_07817_),
    .A2(_08503_),
    .B(_08523_),
    .ZN(_08524_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14230_ (.A1(net529),
    .A2(net3279),
    .Z(_09868_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14231_ (.A1(net3328),
    .A2(net3247),
    .Z(_09867_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14232_ (.A1(net3324),
    .A2(net3321),
    .Z(_09866_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3230 (.I(_08577_),
    .Z(net3230));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14234_ (.A1(net3251),
    .A2(net3318),
    .ZN(_09876_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14235_ (.I0(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .S(net3338),
    .Z(_08526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14236_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(net3407),
    .B1(_08526_),
    .B2(net3659),
    .ZN(_09891_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _14237_ (.I(_07172_),
    .ZN(_08527_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _14238_ (.I(_07859_),
    .ZN(_08528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14239_ (.I0(_08527_),
    .I1(_08528_),
    .S(_08486_),
    .Z(_08529_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14240_ (.A1(net529),
    .A2(net3243),
    .Z(_09896_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14241_ (.A1(net3328),
    .A2(net3279),
    .Z(_09895_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14242_ (.A1(net3324),
    .A2(net3247),
    .Z(_09894_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3232 (.I(net476),
    .Z(net3232));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14244_ (.A1(net3321),
    .A2(net3318),
    .ZN(_09904_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14245_ (.I0(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .S(net3338),
    .Z(_08531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14246_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(net3407),
    .B1(_08531_),
    .B2(net3659),
    .ZN(_09924_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14247_ (.A1(_07220_),
    .A2(_08486_),
    .Z(_08532_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14248_ (.A1(_08503_),
    .A2(_07920_),
    .B(_08532_),
    .ZN(_08533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14249_ (.A1(net529),
    .A2(net3274),
    .Z(_09929_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14250_ (.A1(net3328),
    .A2(net3243),
    .Z(_09928_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14251_ (.A1(net3324),
    .A2(net3279),
    .Z(_09927_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3225 (.I(_10545_[0]),
    .Z(net3225));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14253_ (.A1(net3247),
    .A2(net3318),
    .ZN(_09937_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14254_ (.I0(net412),
    .I1(_07936_),
    .S(_08481_),
    .Z(_08535_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place3228 (.I(net3227),
    .Z(net3228));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_clk_i_regs (.I(clknet_6_29__leaf_clk_i_regs),
    .Z(clknet_leaf_4_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14257_ (.A1(net3330),
    .A2(net3314),
    .ZN(_09947_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14258_ (.I0(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .S(net3338),
    .Z(_08538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14259_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(net3407),
    .B1(_08538_),
    .B2(net3659),
    .ZN(_09960_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14260_ (.A1(net443),
    .A2(_08486_),
    .Z(_08539_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14261_ (.A1(_07957_),
    .A2(_08503_),
    .B(_08539_),
    .ZN(_08540_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14262_ (.A1(net3332),
    .A2(net3272),
    .Z(_09965_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14263_ (.A1(_08501_),
    .A2(_08533_),
    .Z(_09964_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14264_ (.A1(net3326),
    .A2(_08529_),
    .Z(_09963_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3221 (.I(_08676_),
    .Z(net3221));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3613 (.I(net416),
    .Z(net3613));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14267_ (.A1(net3317),
    .A2(net437),
    .ZN(_09973_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14268_ (.A1(net3251),
    .A2(net3314),
    .ZN(_09983_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _14269_ (.A1(_06831_),
    .A2(_06821_),
    .A3(_06817_),
    .A4(_06840_),
    .ZN(_08543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14270_ (.I0(_08543_),
    .I1(_08055_),
    .S(_08481_),
    .Z(_08544_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3231 (.I(net3230),
    .Z(net3231));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14272_ (.A1(net3334),
    .A2(net3313),
    .Z(_09986_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14273_ (.I0(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .S(_08449_),
    .Z(_08546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14274_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(net3407),
    .B1(_08546_),
    .B2(net3659),
    .ZN(_10005_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14275_ (.I(_07278_),
    .ZN(_08547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14276_ (.A1(_08547_),
    .A2(_08503_),
    .ZN(_08548_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14277_ (.A1(_08001_),
    .A2(_08503_),
    .B(_08548_),
    .ZN(_08549_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14278_ (.A1(_08496_),
    .A2(_08549_),
    .Z(_10010_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14279_ (.A1(_08501_),
    .A2(_08540_),
    .Z(_10009_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14280_ (.A1(_08508_),
    .A2(_08533_),
    .Z(_10008_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3233 (.I(net3232),
    .Z(net3233));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14282_ (.A1(net3317),
    .A2(net3244),
    .ZN(_10018_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14283_ (.A1(net3323),
    .A2(net3314),
    .ZN(_10028_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14284_ (.I0(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .S(_08449_),
    .Z(_08551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14285_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(_08481_),
    .B1(_08551_),
    .B2(net3659),
    .ZN(_10044_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14286_ (.A1(_06880_),
    .A2(_08503_),
    .Z(_08552_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14287_ (.A1(_08038_),
    .A2(_08486_),
    .B(_08552_),
    .ZN(_08553_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14288_ (.A1(_08496_),
    .A2(_08553_),
    .Z(_10047_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14289_ (.A1(_08501_),
    .A2(_08549_),
    .Z(_10049_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14290_ (.A1(_08540_),
    .A2(_08508_),
    .Z(_10048_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3224 (.I(net3223),
    .Z(net3224));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14292_ (.A1(_08520_),
    .A2(_08533_),
    .ZN(_10057_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14293_ (.A1(_08517_),
    .A2(_08535_),
    .ZN(_10067_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14294_ (.A1(_08500_),
    .A2(_08544_),
    .Z(_10072_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3220 (.I(_02535_),
    .Z(net3220));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14296_ (.I0(_07346_),
    .I1(_08110_),
    .S(_08481_),
    .Z(_08556_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3226 (.I(_10493_[0]),
    .Z(net3226));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14298_ (.A1(_08507_),
    .A2(_08556_),
    .Z(_10071_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14299_ (.I0(_07389_),
    .I1(_08145_),
    .S(_08481_),
    .Z(_08558_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3219 (.I(_02558_),
    .Z(net3219));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14301_ (.A1(_08488_),
    .A2(_08558_),
    .Z(_10070_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14302_ (.I0(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .S(_08449_),
    .Z(_08560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14303_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(net3407),
    .B1(_08560_),
    .B2(net3659),
    .ZN(_10091_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14304_ (.A1(_06309_),
    .A2(_08486_),
    .Z(_08561_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14305_ (.A1(_08094_),
    .A2(_08503_),
    .B(_08561_),
    .ZN(_08562_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3216 (.I(_10433_[0]),
    .Z(net3216));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14307_ (.A1(_08496_),
    .A2(_08562_),
    .ZN(_10096_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3222 (.I(_08676_),
    .Z(net3222));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14309_ (.A1(_08520_),
    .A2(_08540_),
    .ZN(_10103_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14310_ (.A1(_08524_),
    .A2(_08535_),
    .ZN(_10113_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14311_ (.A1(_08513_),
    .A2(_08544_),
    .Z(_10118_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14312_ (.A1(_08500_),
    .A2(_08556_),
    .Z(_10117_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14313_ (.A1(_08507_),
    .A2(_08558_),
    .Z(_10116_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14314_ (.I0(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .S(_08449_),
    .Z(_08565_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14315_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net3407),
    .B1(_08565_),
    .B2(net3659),
    .ZN(_10141_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14316_ (.I(_08129_),
    .ZN(_08566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14317_ (.I0(_07368_),
    .I1(_08566_),
    .S(_08486_),
    .Z(_08567_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14318_ (.A1(_08496_),
    .A2(_08567_),
    .Z(_10147_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14319_ (.A1(_08501_),
    .A2(_08562_),
    .Z(_10146_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14320_ (.A1(net3326),
    .A2(_08553_),
    .Z(_10145_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3214 (.I(_10436_[0]),
    .Z(net3214));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14322_ (.A1(net3317),
    .A2(net3240),
    .ZN(_10155_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14323_ (.A1(net3244),
    .A2(net3314),
    .ZN(_10164_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14324_ (.A1(net3322),
    .A2(net3313),
    .Z(_10169_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14325_ (.A1(net3249),
    .A2(net3238),
    .Z(_10168_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14326_ (.A1(net3329),
    .A2(net3310),
    .Z(_10167_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14327_ (.A1(_07066_),
    .A2(_08453_),
    .Z(_08569_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14328_ (.A1(_08215_),
    .A2(_08569_),
    .A3(_08486_),
    .Z(_08570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14329_ (.A1(net3335),
    .A2(_08570_),
    .Z(_10187_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14330_ (.I0(_07470_),
    .I1(_08215_),
    .S(_08486_),
    .Z(_08571_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3218 (.I(_02922_),
    .Z(net3218));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14332_ (.I0(net276),
    .I1(_07582_),
    .S(_08481_),
    .Z(_08573_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3223 (.I(_08669_),
    .Z(net3223));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14334_ (.A1(_08571_),
    .A2(net3307),
    .Z(_10194_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _14335_ (.I(_07426_),
    .ZN(_08575_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14336_ (.I(_08177_),
    .ZN(_08576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14337_ (.I0(_08575_),
    .I1(_08576_),
    .S(_08486_),
    .Z(_08577_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14338_ (.A1(net3332),
    .A2(net3230),
    .Z(_10193_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14339_ (.A1(net3327),
    .A2(net3235),
    .Z(_10192_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14340_ (.A1(net3324),
    .A2(net3268),
    .ZN(_10203_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14341_ (.I0(_06653_),
    .I1(_07875_),
    .S(_08481_),
    .Z(_08578_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3210 (.I(_08897_),
    .Z(net3210));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3208 (.I(_08959_),
    .Z(net3208));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14344_ (.A1(net3273),
    .A2(net3306),
    .ZN(_10213_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14345_ (.I0(_06805_),
    .I1(_08017_),
    .S(_08481_),
    .Z(_08581_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14347_ (.A1(net3281),
    .A2(net3259),
    .Z(_10218_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14348_ (.A1(net3248),
    .A2(net3313),
    .Z(_10217_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14349_ (.A1(net3323),
    .A2(net3238),
    .Z(_10216_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14350_ (.A1(net3250),
    .A2(net3310),
    .ZN(_10230_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14351_ (.A1(net3659),
    .A2(_06717_),
    .A3(_07066_),
    .Z(_08583_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3212 (.I(_10497_[0]),
    .Z(net3212));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14353_ (.A1(net3657),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .B1(_08583_),
    .B2(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .ZN(_08585_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _14354_ (.I(_08585_),
    .ZN(_10256_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14355_ (.A1(_08570_),
    .A2(net3307),
    .Z(_10255_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14356_ (.A1(net3332),
    .A2(_08571_),
    .Z(_10261_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14357_ (.A1(net3327),
    .A2(net3230),
    .Z(_10260_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14358_ (.A1(net3324),
    .A2(net3235),
    .Z(_10259_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14359_ (.A1(net3319),
    .A2(net3268),
    .ZN(_10271_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14360_ (.A1(net3315),
    .A2(net3273),
    .ZN(_10281_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14361_ (.A1(net3281),
    .A2(net3313),
    .Z(_10286_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14362_ (.A1(net3248),
    .A2(net3239),
    .Z(_10285_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14363_ (.A1(net3323),
    .A2(net3310),
    .Z(_10284_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14364_ (.I0(_07449_),
    .I1(_08193_),
    .S(_08481_),
    .Z(_08586_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3207 (.I(_03099_),
    .Z(net3207));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_43_clk_i_regs (.I(clknet_6_55__leaf_clk_i_regs),
    .Z(clknet_leaf_43_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14367_ (.A1(net3250),
    .A2(net3301),
    .ZN(_10298_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _14368_ (.A1(net3657),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .A3(_08569_),
    .ZN(_08589_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3203 (.I(_10651_[0]),
    .Z(net3203));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3453 (.I(_06334_),
    .Z(net3453));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14371_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(_08583_),
    .ZN(_08592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14372_ (.A1(_08589_),
    .A2(_08592_),
    .ZN(_10312_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3202 (.I(_10652_[0]),
    .Z(net3202));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14374_ (.A1(net3332),
    .A2(net3265),
    .Z(_10317_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14375_ (.A1(net3327),
    .A2(net3263),
    .Z(_10316_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14376_ (.A1(net3324),
    .A2(net3230),
    .Z(_10315_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_101_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_101_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14378_ (.A1(net3319),
    .A2(net3236),
    .ZN(_10327_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14379_ (.A1(net3315),
    .A2(net3242),
    .ZN(_10337_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14380_ (.A1(net3244),
    .A2(net3313),
    .Z(_10342_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14381_ (.A1(net3281),
    .A2(net3239),
    .Z(_10341_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14382_ (.A1(net3248),
    .A2(net3311),
    .Z(_10340_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14383_ (.A1(net3323),
    .A2(net3302),
    .ZN(_10354_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14384_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(_08583_),
    .ZN(_08595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14385_ (.A1(_08589_),
    .A2(_08595_),
    .ZN(_10370_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14386_ (.A1(net3327),
    .A2(net3265),
    .Z(_10374_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14387_ (.A1(net3324),
    .A2(net3263),
    .Z(_10373_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_100_clk_i_regs (.I(clknet_6_60__leaf_clk_i_regs),
    .Z(clknet_leaf_100_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14389_ (.A1(net3319),
    .A2(net3231),
    .ZN(_10384_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_98_clk_i_regs (.I(clknet_6_60__leaf_clk_i_regs),
    .Z(clknet_leaf_98_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14391_ (.A1(net3315),
    .A2(net3271),
    .ZN(_10393_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14392_ (.A1(net3276),
    .A2(net3313),
    .Z(_10399_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14393_ (.A1(net3245),
    .A2(net3239),
    .Z(_10398_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14394_ (.A1(net3281),
    .A2(net3311),
    .Z(_10397_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14395_ (.A1(net3248),
    .A2(net3302),
    .ZN(_10411_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14396_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(_08583_),
    .ZN(_08598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14397_ (.A1(_08589_),
    .A2(_08598_),
    .ZN(_10428_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14398_ (.A1(net3324),
    .A2(net3265),
    .Z(_10431_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14399_ (.A1(net3319),
    .A2(net3264),
    .ZN(_10439_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14400_ (.A1(net3315),
    .A2(net3269),
    .ZN(_10450_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14401_ (.A1(net3273),
    .A2(net3313),
    .Z(_10454_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14402_ (.A1(net3276),
    .A2(net3239),
    .Z(_10453_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14403_ (.A1(net3245),
    .A2(net3311),
    .Z(_10455_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14404_ (.A1(net3282),
    .A2(net3302),
    .ZN(_10467_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14405_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(net3303),
    .ZN(_08599_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14406_ (.A1(_08589_),
    .A2(_08599_),
    .ZN(_10484_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14407_ (.A1(net3319),
    .A2(net3265),
    .Z(_10493_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14408_ (.I0(_08275_),
    .I1(_07838_),
    .S(_08481_),
    .Z(_08600_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3201 (.I(_08910_),
    .Z(net3201));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14410_ (.A1(net3264),
    .A2(net3300),
    .Z(_10492_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14411_ (.A1(net3231),
    .A2(net3306),
    .Z(_10491_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14412_ (.A1(net3315),
    .A2(net3237),
    .ZN(_10505_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14413_ (.A1(net3313),
    .A2(net3242),
    .Z(_10510_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14414_ (.A1(net3273),
    .A2(net3239),
    .Z(_10509_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14415_ (.A1(net479),
    .A2(net3311),
    .Z(_10508_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14416_ (.A1(net3246),
    .A2(net3302),
    .ZN(_10522_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14417_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(net3303),
    .ZN(_08602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14418_ (.A1(_08589_),
    .A2(_08602_),
    .ZN(_10539_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14419_ (.A1(net3265),
    .A2(net3300),
    .Z(_10545_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14420_ (.A1(net3264),
    .A2(net3306),
    .Z(_10544_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14421_ (.A1(net3315),
    .A2(net3231),
    .ZN(_10557_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14422_ (.A1(net3313),
    .A2(net3271),
    .Z(_10562_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14423_ (.A1(net3242),
    .A2(net3239),
    .Z(_10561_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14424_ (.A1(net3273),
    .A2(net3311),
    .Z(_10560_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14425_ (.A1(net479),
    .A2(net3302),
    .ZN(_10574_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14426_ (.A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .A2(net3303),
    .ZN(_08603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14427_ (.A1(_08589_),
    .A2(_08603_),
    .ZN(_10591_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14428_ (.A1(net3265),
    .A2(net3306),
    .Z(_10598_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14429_ (.A1(net3315),
    .A2(net3264),
    .ZN(_10610_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14430_ (.A1(net3313),
    .A2(net3269),
    .Z(_10615_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14431_ (.A1(net3271),
    .A2(net3239),
    .Z(_10614_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14432_ (.A1(net3242),
    .A2(net3311),
    .Z(_10613_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14433_ (.A1(net3273),
    .A2(net3302),
    .ZN(_10627_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14434_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(net3303),
    .ZN(_08604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14435_ (.A1(_08589_),
    .A2(_08604_),
    .ZN(_10644_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14436_ (.A1(net3315),
    .A2(net3266),
    .Z(_10658_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14437_ (.I0(net407),
    .I1(_07973_),
    .S(_08481_),
    .Z(_08605_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14439_ (.A1(net3264),
    .A2(net3297),
    .Z(_10657_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14440_ (.A1(net3231),
    .A2(net3260),
    .Z(_10656_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14441_ (.A1(net3313),
    .A2(net3237),
    .Z(_10663_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14442_ (.A1(net3239),
    .A2(net3269),
    .Z(_10662_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14443_ (.A1(net3271),
    .A2(net3311),
    .Z(_10661_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14444_ (.A1(net3242),
    .A2(net3302),
    .ZN(_10677_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14445_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(net3303),
    .ZN(_08607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14446_ (.A1(_08589_),
    .A2(_08607_),
    .ZN(_10694_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14447_ (.A1(net3266),
    .A2(net3297),
    .Z(_10704_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14448_ (.A1(net3264),
    .A2(net3260),
    .Z(_10703_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14449_ (.A1(net3313),
    .A2(net3231),
    .Z(_10708_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14450_ (.A1(net3239),
    .A2(net3237),
    .Z(_10707_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14451_ (.A1(net3311),
    .A2(net3269),
    .Z(_10709_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14452_ (.A1(net3271),
    .A2(net3302),
    .ZN(_10724_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14453_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(net3303),
    .ZN(_08608_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14454_ (.A1(_08589_),
    .A2(_08608_),
    .ZN(_10741_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14455_ (.A1(net3266),
    .A2(net3260),
    .Z(_10748_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14456_ (.A1(net3313),
    .A2(net3264),
    .Z(_10753_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14457_ (.A1(net3239),
    .A2(net3231),
    .Z(_10752_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14458_ (.A1(net3311),
    .A2(net3237),
    .Z(_10751_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14459_ (.A1(net3269),
    .A2(net3302),
    .ZN(_10768_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14460_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(net3303),
    .ZN(_08609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14461_ (.A1(_08589_),
    .A2(_08609_),
    .ZN(_10785_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14462_ (.A1(net3313),
    .A2(net3266),
    .Z(_10794_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14463_ (.A1(net3239),
    .A2(net3264),
    .Z(_10793_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14464_ (.A1(net3311),
    .A2(net3231),
    .Z(_10792_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14465_ (.A1(net3237),
    .A2(net3302),
    .ZN(_10809_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14466_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(net3303),
    .ZN(_08610_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14467_ (.A1(_08589_),
    .A2(_08610_),
    .ZN(_10826_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14468_ (.A1(net3239),
    .A2(net3266),
    .Z(_10834_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14469_ (.A1(net3311),
    .A2(net3264),
    .Z(_10833_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14470_ (.A1(net3231),
    .A2(net3302),
    .ZN(_10848_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14471_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(net3303),
    .ZN(_08611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14472_ (.A1(_08589_),
    .A2(_08611_),
    .ZN(_10865_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14473_ (.A1(net3311),
    .A2(net3266),
    .Z(_10872_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14474_ (.A1(net3264),
    .A2(net3302),
    .ZN(_10886_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14475_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(net3303),
    .ZN(_08612_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14476_ (.A1(_08589_),
    .A2(_08612_),
    .ZN(_10903_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14477_ (.A1(net3266),
    .A2(net3302),
    .Z(_10921_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14478_ (.I0(_07486_),
    .I1(_08231_),
    .S(_08481_),
    .Z(_08613_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14480_ (.A1(net3264),
    .A2(net3294),
    .Z(_10920_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14481_ (.A1(_07066_),
    .A2(net431),
    .A3(_08460_),
    .Z(_08615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14482_ (.A1(_08615_),
    .A2(_08481_),
    .ZN(_08616_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_97_clk_i_regs (.I(clknet_6_60__leaf_clk_i_regs),
    .Z(clknet_leaf_97_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14484_ (.A1(net3231),
    .A2(net3256),
    .ZN(_10919_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14485_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net3303),
    .ZN(_08618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14486_ (.A1(_08589_),
    .A2(_08618_),
    .ZN(_10940_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14487_ (.A1(net3266),
    .A2(net3294),
    .Z(_10952_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14488_ (.A1(net3264),
    .A2(net3256),
    .ZN(_10951_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14489_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A2(net3303),
    .ZN(_08619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14490_ (.A1(_08589_),
    .A2(_08619_),
    .ZN(_10971_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14491_ (.A1(net3266),
    .A2(net3256),
    .ZN(_10982_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14492_ (.I(net3216),
    .ZN(_10436_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14493_ (.I(_10914_[0]),
    .ZN(_10915_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14494_ (.A1(_06241_),
    .A2(_06344_),
    .B(_06245_),
    .ZN(_08620_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14495_ (.A1(_06246_),
    .A2(_06224_),
    .A3(_08404_),
    .A4(_08620_),
    .Z(_08621_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14496_ (.A1(_06782_),
    .A2(_08621_),
    .B(\id_stage_i.branch_set ),
    .ZN(_08622_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3662 (.I(net3661),
    .Z(net3662));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14498_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_08360_),
    .A3(_08362_),
    .Z(_08624_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_95_clk_i_regs (.I(clknet_6_62__leaf_clk_i_regs),
    .Z(clknet_leaf_95_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14500_ (.A1(net3473),
    .A2(\id_stage_i.controller_i.instr_fetch_err_i ),
    .ZN(_08626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14501_ (.A1(_08624_),
    .A2(_08626_),
    .ZN(_08627_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _14502_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.exc_req_q ),
    .A3(\id_stage_i.controller_i.load_err_q ),
    .Z(_08628_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14503_ (.A1(_08391_),
    .A2(_08628_),
    .ZN(_08629_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14504_ (.I(\cs_registers_i.priv_mode_id_o[1] ),
    .ZN(_11156_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14505_ (.A1(\cs_registers_i.dcsr_q[12] ),
    .A2(_11156_[0]),
    .ZN(_08630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14506_ (.A1(\cs_registers_i.dcsr_q[15] ),
    .A2(_08381_),
    .ZN(_08631_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14507_ (.A1(\cs_registers_i.priv_mode_id_o[0] ),
    .A2(_08630_),
    .B(_08631_),
    .ZN(_08632_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14508_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_08632_),
    .Z(_08633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14509_ (.A1(net3473),
    .A2(\id_stage_i.controller_i.instr_fetch_err_i ),
    .Z(_08634_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14510_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_08634_),
    .ZN(_08635_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14511_ (.A1(net3560),
    .A2(_08393_),
    .A3(_08635_),
    .Z(_08636_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14512_ (.A1(_08633_),
    .A2(_08636_),
    .Z(_08637_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14513_ (.I(\cs_registers_i.nmi_mode_i ),
    .ZN(_08638_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14514_ (.A1(net145),
    .A2(\cs_registers_i.csr_mstatus_mie_o ),
    .Z(_08639_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14515_ (.A1(_08370_),
    .A2(_08638_),
    .A3(_08639_),
    .Z(_08640_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _14516_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_08390_),
    .A3(_08640_),
    .ZN(_08641_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14517_ (.I(_08641_),
    .ZN(_08642_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14518_ (.A1(\cs_registers_i.mie_q[14] ),
    .A2(net135),
    .ZN(_08643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14519_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net141),
    .B1(\cs_registers_i.mie_q[7] ),
    .B2(net142),
    .ZN(_08644_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14520_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net139),
    .B1(\cs_registers_i.mie_q[5] ),
    .B2(net140),
    .ZN(_08645_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14521_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net137),
    .B1(\cs_registers_i.mie_q[3] ),
    .B2(net138),
    .ZN(_08646_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14522_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(net130),
    .B1(\cs_registers_i.mie_q[1] ),
    .B2(net136),
    .ZN(_08647_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _14523_ (.A1(_08644_),
    .A2(_08645_),
    .A3(_08646_),
    .A4(_08647_),
    .Z(_08648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14524_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(net133),
    .B1(\cs_registers_i.mie_q[13] ),
    .B2(net134),
    .ZN(_08649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14525_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net131),
    .B1(\cs_registers_i.mie_q[11] ),
    .B2(net132),
    .ZN(_08650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14526_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net143),
    .B1(\cs_registers_i.mie_q[9] ),
    .B2(net144),
    .ZN(_08651_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14527_ (.A1(_08649_),
    .A2(_08650_),
    .A3(_08651_),
    .Z(_08652_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14528_ (.A1(_08643_),
    .A2(_08648_),
    .A3(_08652_),
    .Z(_08653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14529_ (.A1(\cs_registers_i.mie_q[16] ),
    .A2(net147),
    .B(net145),
    .ZN(_08654_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _14530_ (.A1(net129),
    .A2(\cs_registers_i.mie_q[15] ),
    .B1(\cs_registers_i.mie_q[17] ),
    .B2(net146),
    .ZN(_08655_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _14531_ (.A1(_08653_),
    .A2(_08654_),
    .A3(_08655_),
    .ZN(_08656_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14532_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(net60),
    .Z(_08657_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _14533_ (.I(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .ZN(_08658_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14534_ (.A1(_08360_),
    .A2(_08658_),
    .Z(_08659_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14535_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_08659_),
    .Z(_08660_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14536_ (.A1(_08389_),
    .A2(_08660_),
    .Z(_08661_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _14537_ (.A1(_08642_),
    .A2(net3354),
    .B1(_08657_),
    .B2(_08661_),
    .ZN(_08662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14538_ (.A1(_08389_),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .ZN(_08663_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _14539_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.exc_req_q ),
    .A3(\id_stage_i.controller_i.load_err_q ),
    .ZN(_08664_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14540_ (.A1(_08391_),
    .A2(_08664_),
    .Z(_08665_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14541_ (.A1(_06733_),
    .A2(_08379_),
    .Z(_08666_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14542_ (.A1(_08659_),
    .A2(_08663_),
    .B1(_08665_),
    .B2(_08666_),
    .ZN(_08667_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14543_ (.A1(_08662_),
    .A2(_08667_),
    .Z(_08668_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _14544_ (.A1(_08622_),
    .A2(_08627_),
    .B1(_08629_),
    .B2(_08637_),
    .C(_08668_),
    .ZN(_08669_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3199 (.I(_08928_),
    .Z(net3199));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3091 (.I(_01951_),
    .Z(net3091));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3194 (.I(_01984_),
    .Z(net3194));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14548_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .A2(_08669_),
    .Z(_08673_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14549_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_08673_),
    .Z(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14550_ (.A1(_08622_),
    .A2(_08627_),
    .ZN(_08674_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14551_ (.A1(_08629_),
    .A2(_08637_),
    .B(_08668_),
    .ZN(_08675_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14552_ (.A1(_08674_),
    .A2(_08675_),
    .ZN(_08676_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place3195 (.I(_07013_),
    .Z(net3195));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3191 (.I(_02669_),
    .Z(net3191));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3092 (.I(_03750_),
    .Z(net3092));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14556_ (.I0(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .I1(_08385_),
    .S(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .Z(_08680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14557_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_08659_),
    .ZN(_08681_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14558_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_08628_),
    .B(_08390_),
    .ZN(_08682_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14559_ (.A1(_08681_),
    .A2(_08682_),
    .ZN(_08683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14560_ (.A1(_08380_),
    .A2(_08665_),
    .Z(_08684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _14561_ (.A1(_08362_),
    .A2(_08680_),
    .B(_08683_),
    .C(_08684_),
    .ZN(_08685_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3643 (.I(net449),
    .Z(net3643));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3100 (.I(_03521_),
    .Z(net3100));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer572 (.I(_07153_),
    .Z(net858));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3120 (.I(_11279_[0]),
    .Z(net3120));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14566_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(net3674),
    .Z(_08690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14567_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net3666),
    .ZN(_08691_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14568_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net3668),
    .Z(_08692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14569_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net3672),
    .ZN(_08693_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14570_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(net3673),
    .A3(_08693_),
    .Z(_08694_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14571_ (.A1(\cs_registers_i.mie_q[3] ),
    .A2(net3671),
    .B(_08694_),
    .ZN(_08695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14572_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net3670),
    .B(_08695_),
    .ZN(_08696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14573_ (.A1(\cs_registers_i.mie_q[5] ),
    .A2(net3669),
    .B(_08696_),
    .ZN(_08697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14574_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(net3667),
    .ZN(_08698_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14575_ (.A1(_08692_),
    .A2(_08697_),
    .B(_08698_),
    .ZN(_08699_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14576_ (.A1(\cs_registers_i.mie_q[9] ),
    .A2(net3665),
    .B1(_08691_),
    .B2(_08699_),
    .ZN(_08700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14577_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net3677),
    .B(_08700_),
    .ZN(_08701_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14578_ (.A1(\cs_registers_i.mie_q[11] ),
    .A2(net3676),
    .B(_08701_),
    .ZN(_08702_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14579_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(net3675),
    .B(_08702_),
    .ZN(_08703_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _14580_ (.A1(_08690_),
    .A2(_08703_),
    .B(_08643_),
    .ZN(_08704_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14581_ (.A1(_08638_),
    .A2(net145),
    .B(net3382),
    .ZN(_08705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14582_ (.A1(_08642_),
    .A2(net3354),
    .ZN(_08706_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14583_ (.A1(_08704_),
    .A2(_08705_),
    .B(_08706_),
    .ZN(_08707_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3518 (.I(net3516),
    .Z(net3518));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14585_ (.A1(_08385_),
    .A2(_08665_),
    .Z(_08709_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14586_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(_08684_),
    .B1(_08709_),
    .B2(\cs_registers_i.csr_mepc_o[2] ),
    .ZN(_08710_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14587_ (.I(_08710_),
    .ZN(_08711_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14588_ (.A1(_08624_),
    .A2(net171),
    .B(_08707_),
    .C(_08711_),
    .ZN(_08712_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _14589_ (.A1(_08676_),
    .A2(net3254),
    .A3(_08712_),
    .Z(_08713_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14590_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .A2(_08676_),
    .ZN(_08714_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14591_ (.A1(_08713_),
    .A2(_08714_),
    .ZN(_11660_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14592_ (.I(net3405),
    .ZN(_08715_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14593_ (.A1(_08715_),
    .A2(net3404),
    .B(net3406),
    .ZN(_08716_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14594_ (.A1(net3401),
    .A2(_08716_),
    .ZN(_08717_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14595_ (.A1(net3402),
    .A2(_08717_),
    .ZN(_08718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14596_ (.A1(_08638_),
    .A2(net145),
    .ZN(_08719_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14597_ (.A1(_08643_),
    .A2(_08719_),
    .Z(_08720_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14598_ (.I(_08720_),
    .ZN(_08721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14599_ (.A1(net3403),
    .A2(_08718_),
    .B(_08721_),
    .C(net3382),
    .ZN(_08722_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14600_ (.A1(_08706_),
    .A2(_08722_),
    .Z(_08723_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14601_ (.A1(_08391_),
    .A2(_08628_),
    .Z(_08724_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14602_ (.A1(_08624_),
    .A2(net174),
    .B1(_08724_),
    .B2(\cs_registers_i.debug_mode_i ),
    .ZN(_08725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14603_ (.A1(\cs_registers_i.csr_depc_o[3] ),
    .A2(_08684_),
    .B1(_08709_),
    .B2(\cs_registers_i.csr_mepc_o[3] ),
    .ZN(_08726_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14604_ (.A1(_08723_),
    .A2(_08725_),
    .A3(_08726_),
    .Z(_08727_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _14605_ (.A1(_08676_),
    .A2(net3254),
    .A3(_08727_),
    .Z(_08728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14606_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .A2(_08676_),
    .ZN(_08729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14607_ (.A1(_08728_),
    .A2(_08729_),
    .ZN(_11663_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _14608_ (.I(\cs_registers_i.pc_if_i[1] ),
    .ZN(_08730_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3517 (.I(net559),
    .Z(net3517));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3136 (.I(_11337_[0]),
    .Z(net3136));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14611_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .ZN(_08733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14612_ (.A1(net107),
    .A2(net96),
    .B(net94),
    .ZN(_08734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3190 (.I(_03218_),
    .Z(net3190));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _14614_ (.I(net3652),
    .ZN(_08736_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3137 (.I(net3136),
    .Z(net3137));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14616_ (.I0(_08733_),
    .I1(_08734_),
    .S(_08736_),
    .Z(_08738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14617_ (.A1(_08730_),
    .A2(_08738_),
    .ZN(_08739_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3134 (.I(_11343_[0]),
    .Z(net3134));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14619_ (.A1(net3652),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .Z(_08741_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14620_ (.A1(_08736_),
    .A2(net104),
    .A3(net103),
    .Z(_08742_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14621_ (.A1(_08741_),
    .A2(_08742_),
    .Z(_08743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14622_ (.I0(net94),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_08744_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _14623_ (.A1(_08743_),
    .A2(_08744_),
    .Z(_08745_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14624_ (.I(_08745_),
    .ZN(_08746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14625_ (.A1(net3653),
    .A2(_08746_),
    .ZN(_10998_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14626_ (.A1(_08739_),
    .A2(_10998_[0]),
    .Z(_11388_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14627_ (.I(_11388_[0]),
    .ZN(_10999_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14628_ (.I(net149),
    .ZN(_08747_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _14629_ (.A1(net60),
    .A2(core_busy_q),
    .A3(_08656_),
    .B(fetch_enable_q),
    .ZN(net150));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14630_ (.A1(_08747_),
    .A2(net150),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3452 (.I(net3450),
    .Z(net3452));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14632_ (.A1(net3334),
    .A2(net3309),
    .ZN(_09749_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3145 (.I(_11318_[0]),
    .Z(net3145));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14634_ (.A1(net3337),
    .A2(net3330),
    .ZN(_09754_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14635_ (.A1(net3330),
    .A2(net3309),
    .ZN(_09764_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14636_ (.A1(net3251),
    .A2(net3309),
    .ZN(_09772_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14637_ (.A1(net3321),
    .A2(net481),
    .ZN(_09790_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14638_ (.A1(net3285),
    .A2(net3325),
    .ZN(_09795_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14639_ (.A1(net3247),
    .A2(net481),
    .ZN(_09805_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14640_ (.A1(net3333),
    .A2(net3305),
    .ZN(_09839_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14641_ (.I(_11220_[0]),
    .ZN(_09856_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14642_ (.A1(net3243),
    .A2(net481),
    .ZN(_09861_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14643_ (.A1(net3285),
    .A2(net3305),
    .ZN(_09874_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14644_ (.A1(net3274),
    .A2(net3307),
    .ZN(_09889_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14645_ (.A1(net3330),
    .A2(net3305),
    .ZN(_09902_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14646_ (.A1(net3272),
    .A2(net478),
    .ZN(_09922_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14647_ (.A1(net3251),
    .A2(net3305),
    .ZN(_09935_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3146 (.I(_11313_[0]),
    .Z(net3146));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14649_ (.A1(net3334),
    .A2(net3258),
    .ZN(_09945_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14650_ (.A1(net3241),
    .A2(net3307),
    .ZN(_09958_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14651_ (.A1(net3321),
    .A2(net3304),
    .ZN(_09971_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14652_ (.A1(net3284),
    .A2(net3258),
    .ZN(_09981_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14653_ (.A1(net3270),
    .A2(net482),
    .ZN(_10003_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14654_ (.A1(net3247),
    .A2(net3304),
    .ZN(_10016_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14655_ (.A1(net3329),
    .A2(net3257),
    .ZN(_10026_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14656_ (.A1(_08562_),
    .A2(_08573_),
    .ZN(_10042_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14657_ (.A1(net3278),
    .A2(_08578_),
    .ZN(_10055_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14658_ (.A1(net3249),
    .A2(_08581_),
    .ZN(_10065_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14659_ (.A1(_08567_),
    .A2(_08573_),
    .ZN(_10089_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14660_ (.A1(_08508_),
    .A2(_08549_),
    .ZN(_10094_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14661_ (.A1(_08529_),
    .A2(_08578_),
    .ZN(_10101_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14662_ (.A1(_08511_),
    .A2(_08581_),
    .ZN(_10111_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14663_ (.A1(net3335),
    .A2(_08571_),
    .ZN(_10140_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14664_ (.A1(net3275),
    .A2(net3304),
    .ZN(_10153_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14665_ (.A1(net3248),
    .A2(net3257),
    .ZN(_10162_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3151 (.I(_11264_[0]),
    .Z(net3151));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14667_ (.A1(net3242),
    .A2(net3300),
    .ZN(_10201_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3161 (.I(_11220_[0]),
    .Z(net3161));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14669_ (.A1(net3244),
    .A2(net3297),
    .ZN(_10211_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3162 (.I(_04319_),
    .Z(net3162));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14671_ (.A1(net3284),
    .A2(_08613_),
    .ZN(_10228_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14672_ (.A1(net3333),
    .A2(net3255),
    .Z(_10237_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14673_ (.A1(net3242),
    .A2(net3306),
    .ZN(_10269_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14674_ (.A1(net3244),
    .A2(net3259),
    .ZN(_10279_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14675_ (.A1(net3284),
    .A2(_08616_),
    .Z(_10296_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14676_ (.A1(net3271),
    .A2(net3306),
    .ZN(_10325_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14677_ (.A1(net3276),
    .A2(net3259),
    .ZN(_10335_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14678_ (.A1(net3329),
    .A2(net3255),
    .Z(_10352_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14679_ (.A1(net3269),
    .A2(net3306),
    .ZN(_10382_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14680_ (.A1(net3242),
    .A2(net3297),
    .ZN(_10392_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14681_ (.A1(net3250),
    .A2(net3255),
    .Z(_10409_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14682_ (.A1(net3236),
    .A2(net3306),
    .ZN(_10437_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14683_ (.A1(net3242),
    .A2(net3260),
    .ZN(_10448_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14684_ (.A1(net3323),
    .A2(net3255),
    .Z(_10465_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14685_ (.A1(net3271),
    .A2(net3260),
    .ZN(_10503_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14686_ (.A1(net3248),
    .A2(net3255),
    .Z(_10520_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14687_ (.A1(net3269),
    .A2(net3260),
    .ZN(_10555_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14688_ (.A1(net3282),
    .A2(net3256),
    .Z(_10572_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14689_ (.A1(net3237),
    .A2(net3260),
    .ZN(_10608_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14690_ (.A1(net3246),
    .A2(net3256),
    .Z(_10625_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14691_ (.A1(net479),
    .A2(net3256),
    .Z(_10675_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14692_ (.A1(net3273),
    .A2(net3256),
    .Z(_10722_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14693_ (.A1(net3242),
    .A2(net3256),
    .Z(_10766_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14694_ (.A1(net3271),
    .A2(net3256),
    .Z(_10807_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14695_ (.A1(net3269),
    .A2(net3256),
    .Z(_10846_[0]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14696_ (.A1(net3237),
    .A2(net3256),
    .Z(_10884_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14697_ (.A1(net3337),
    .A2(net3251),
    .ZN(_09765_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14698_ (.A1(net3337),
    .A2(net3321),
    .ZN(_09773_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14699_ (.A1(net3336),
    .A2(net3247),
    .ZN(_09791_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14700_ (.A1(net3330),
    .A2(net3328),
    .ZN(_09796_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14701_ (.A1(net3336),
    .A2(net3279),
    .ZN(_09806_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14702_ (.A1(net3279),
    .A2(net481),
    .ZN(_09827_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14703_ (.A1(net3285),
    .A2(net3299),
    .ZN(_09840_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14704_ (.I(_11218_[0]),
    .ZN(_09857_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14705_ (.A1(net3336),
    .A2(net3274),
    .ZN(_09862_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14706_ (.A1(net3330),
    .A2(net3299),
    .ZN(_09875_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14707_ (.A1(net3336),
    .A2(net446),
    .ZN(_09890_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14708_ (.A1(net3251),
    .A2(net3299),
    .ZN(_09903_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14709_ (.A1(net3336),
    .A2(net3241),
    .ZN(_09923_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14710_ (.A1(net3321),
    .A2(net3299),
    .ZN(_09936_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14711_ (.A1(net3284),
    .A2(net3295),
    .ZN(_09946_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14712_ (.A1(net3336),
    .A2(net3270),
    .ZN(_09959_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14713_ (.A1(net3247),
    .A2(net3298),
    .ZN(_09972_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14714_ (.A1(net3330),
    .A2(net3296),
    .ZN(_09982_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14715_ (.A1(net577),
    .A2(net3268),
    .ZN(_10004_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14716_ (.A1(net3280),
    .A2(net3298),
    .ZN(_10017_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14717_ (.A1(net3251),
    .A2(net3296),
    .ZN(_10027_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14718_ (.A1(_08484_),
    .A2(_08567_),
    .ZN(_10043_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14719_ (.A1(_08529_),
    .A2(_08600_),
    .ZN(_10056_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14720_ (.A1(_08511_),
    .A2(_08605_),
    .ZN(_10066_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14721_ (.A1(_08484_),
    .A2(_08577_),
    .ZN(_10090_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14722_ (.A1(_08501_),
    .A2(_08553_),
    .ZN(_10095_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14723_ (.A1(_08533_),
    .A2(_08600_),
    .ZN(_10102_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14724_ (.A1(_08517_),
    .A2(_08605_),
    .ZN(_10112_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14725_ (.A1(net3272),
    .A2(net3298),
    .ZN(_10154_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14726_ (.A1(net3280),
    .A2(net3296),
    .ZN(_10163_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14727_ (.A1(net3319),
    .A2(net3270),
    .ZN(_10202_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14728_ (.A1(net3276),
    .A2(net3315),
    .ZN(_10212_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14729_ (.A1(net3329),
    .A2(_08586_),
    .ZN(_10229_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14730_ (.I(_11283_[0]),
    .ZN(_10238_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14731_ (.A1(net3270),
    .A2(net3300),
    .ZN(_10270_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14732_ (.A1(net3276),
    .A2(net3297),
    .ZN(_10280_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14733_ (.A1(net3329),
    .A2(net3293),
    .ZN(_10297_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14734_ (.A1(net3269),
    .A2(net3300),
    .ZN(_10326_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14735_ (.A1(net3273),
    .A2(net3297),
    .ZN(_10336_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14736_ (.A1(net3250),
    .A2(net3294),
    .ZN(_10353_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14737_ (.A1(net3236),
    .A2(net3300),
    .ZN(_10383_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14738_ (.A1(net3323),
    .A2(net3294),
    .ZN(_10410_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14739_ (.A1(net3231),
    .A2(net3300),
    .ZN(_10438_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14740_ (.A1(net3271),
    .A2(net3297),
    .ZN(_10449_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14741_ (.A1(net3248),
    .A2(net3294),
    .ZN(_10466_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14742_ (.A1(net3269),
    .A2(net3297),
    .ZN(_10504_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14743_ (.A1(net3282),
    .A2(net3294),
    .ZN(_10521_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14744_ (.A1(net3237),
    .A2(net3297),
    .ZN(_10556_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14745_ (.A1(net3246),
    .A2(net3294),
    .ZN(_10573_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14746_ (.A1(net3231),
    .A2(net3297),
    .ZN(_10609_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14747_ (.A1(net479),
    .A2(net3294),
    .ZN(_10626_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14748_ (.A1(net3273),
    .A2(net3294),
    .ZN(_10676_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14749_ (.A1(net3242),
    .A2(net3294),
    .ZN(_10723_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14750_ (.A1(net3271),
    .A2(net3294),
    .ZN(_10767_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14751_ (.A1(net3269),
    .A2(net3294),
    .ZN(_10808_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14752_ (.A1(net3237),
    .A2(net3294),
    .ZN(_10847_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14753_ (.A1(net3231),
    .A2(net3294),
    .ZN(_10885_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14754_ (.A1(net3337),
    .A2(net3285),
    .ZN(_09751_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14755_ (.A1(net3285),
    .A2(net3309),
    .ZN(_09756_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14756_ (.A1(net529),
    .A2(net3251),
    .ZN(_09797_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14757_ (.A1(net3336),
    .A2(net3243),
    .ZN(_09828_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14758_ (.A1(net3307),
    .A2(net3230),
    .ZN(_10142_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14759_ (.A1(net3273),
    .A2(net3260),
    .ZN(_10394_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14760_ (.I(_09882_[0]),
    .ZN(_09883_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14761_ (.I(_09910_[0]),
    .ZN(_09911_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14762_ (.I(_10082_[0]),
    .ZN(_10083_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14763_ (.I(_10128_[0]),
    .ZN(_10129_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14764_ (.I(_09781_[0]),
    .ZN(_09782_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14765_ (.I(_09814_[0]),
    .ZN(_09815_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14766_ (.I(_09835_[0]),
    .ZN(_09836_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14767_ (.I(_09847_[0]),
    .ZN(_09848_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14768_ (.I(_09870_[0]),
    .ZN(_09871_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14769_ (.I(_09898_[0]),
    .ZN(_09899_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14770_ (.I(_09931_[0]),
    .ZN(_09932_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14771_ (.I(_09967_[0]),
    .ZN(_09968_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14772_ (.I(_09994_[0]),
    .ZN(_09995_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14773_ (.I(_10012_[0]),
    .ZN(_10013_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14774_ (.I(_10051_[0]),
    .ZN(_10052_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14775_ (.I(_10074_[0]),
    .ZN(_10075_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14776_ (.I(_10120_[0]),
    .ZN(_10121_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14777_ (.I(_10149_[0]),
    .ZN(_10150_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14778_ (.I(_10171_[0]),
    .ZN(_10172_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14779_ (.I(_10191_[0]),
    .ZN(_10198_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14780_ (.I(_10196_[0]),
    .ZN(_10197_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14781_ (.I(_10220_[0]),
    .ZN(_10221_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14782_ (.I(_10236_[0]),
    .ZN(_10239_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14783_ (.I(_10246_[0]),
    .ZN(_10247_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14784_ (.I(_10258_[0]),
    .ZN(_10266_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14785_ (.I(_10263_[0]),
    .ZN(_10264_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14786_ (.I(_10288_[0]),
    .ZN(_10289_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14787_ (.I(_10314_[0]),
    .ZN(_10322_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14788_ (.I(_10319_[0]),
    .ZN(_10320_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14789_ (.I(_10344_[0]),
    .ZN(_10345_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14790_ (.I(_10364_[0]),
    .ZN(_10365_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14791_ (.I(_10372_[0]),
    .ZN(_10379_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14792_ (.I(_10376_[0]),
    .ZN(_10377_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14793_ (.I(_10401_[0]),
    .ZN(_10402_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14794_ (.I(_10421_[0]),
    .ZN(_10422_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14795_ (.I(_10435_[0]),
    .ZN(_10445_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14796_ (.I(_10457_[0]),
    .ZN(_10458_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14797_ (.I(_10477_[0]),
    .ZN(_10478_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14798_ (.I(_10486_[0]),
    .ZN(_10488_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14799_ (.I(_10495_[0]),
    .ZN(_10496_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14800_ (.I(_10512_[0]),
    .ZN(_10513_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14801_ (.I(_10532_[0]),
    .ZN(_10533_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14802_ (.I(_10543_[0]),
    .ZN(_10552_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14803_ (.I(_10547_[0]),
    .ZN(_10549_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14804_ (.I(_10564_[0]),
    .ZN(_10565_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14805_ (.I(_10584_[0]),
    .ZN(_10585_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14806_ (.I(_10593_[0]),
    .ZN(_10595_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14807_ (.I(_10600_[0]),
    .ZN(_10602_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14808_ (.I(_10617_[0]),
    .ZN(_10618_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14809_ (.I(_10637_[0]),
    .ZN(_10638_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14810_ (.I(_10655_[0]),
    .ZN(_10672_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14811_ (.I(_10660_[0]),
    .ZN(_10667_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14812_ (.I(_10665_[0]),
    .ZN(_10666_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14813_ (.I(_10687_[0]),
    .ZN(_10688_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14814_ (.I(_10698_[0]),
    .ZN(_10700_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14815_ (.I(_10706_[0]),
    .ZN(_10713_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14816_ (.I(_10711_[0]),
    .ZN(_10714_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14817_ (.I(_10734_[0]),
    .ZN(_10735_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14818_ (.I(_10747_[0]),
    .ZN(_10763_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14819_ (.I(_10750_[0]),
    .ZN(_10758_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14820_ (.I(_10755_[0]),
    .ZN(_10756_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14821_ (.I(_10778_[0]),
    .ZN(_10779_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14822_ (.I(_10791_[0]),
    .ZN(_10804_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14823_ (.I(_10796_[0]),
    .ZN(_10797_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14824_ (.I(_10819_[0]),
    .ZN(_10820_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14825_ (.I(_10832_[0]),
    .ZN(_10843_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14826_ (.I(_10836_[0]),
    .ZN(_10837_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14827_ (.I(_10858_[0]),
    .ZN(_10859_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14828_ (.I(_10871_[0]),
    .ZN(_10881_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14829_ (.I(_10874_[0]),
    .ZN(_10875_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14830_ (.I(_10896_[0]),
    .ZN(_10897_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14831_ (.I(_10905_[0]),
    .ZN(_10907_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14832_ (.I(_10918_[0]),
    .ZN(_10934_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14833_ (.I(_10923_[0]),
    .ZN(_10924_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14834_ (.I(_10932_[0]),
    .ZN(_10933_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14835_ (.I(_10942_[0]),
    .ZN(_10944_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14836_ (.I(_10954_[0]),
    .ZN(_10956_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14837_ (.I(_10963_[0]),
    .ZN(_10964_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14838_ (.I(_10973_[0]),
    .ZN(_10975_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14839_ (.I(_10990_[0]),
    .ZN(_10991_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14840_ (.I(_09798_[0]),
    .ZN(_11214_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14841_ (.I(_09897_[0]),
    .ZN(_09940_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14842_ (.I(_09930_[0]),
    .ZN(_09976_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14843_ (.I(_09966_[0]),
    .ZN(_10021_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14844_ (.I(_09989_[0]),
    .ZN(_10034_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14845_ (.I(_09993_[0]),
    .ZN(_10039_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14846_ (.I(_10011_[0]),
    .ZN(_10060_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14847_ (.I(_10050_[0]),
    .ZN(_10106_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14848_ (.I(_10148_[0]),
    .ZN(_10206_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14849_ (.I(_10190_[0]),
    .ZN(_10265_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14850_ (.I(_10195_[0]),
    .ZN(_10274_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14851_ (.I(_10219_[0]),
    .ZN(_10301_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14852_ (.I(_10245_[0]),
    .ZN(_10309_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14853_ (.I(_10257_[0]),
    .ZN(_10321_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14854_ (.I(_10262_[0]),
    .ZN(_10330_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14855_ (.I(_10287_[0]),
    .ZN(_10357_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14856_ (.I(_10313_[0]),
    .ZN(_10378_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14857_ (.I(_10318_[0]),
    .ZN(_10387_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14858_ (.I(_10343_[0]),
    .ZN(_10414_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14859_ (.I(_10363_[0]),
    .ZN(_10425_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14860_ (.I(_10375_[0]),
    .ZN(_10442_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14861_ (.I(_10400_[0]),
    .ZN(_10470_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14862_ (.I(_10420_[0]),
    .ZN(_10481_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14863_ (.I(_10429_[0]),
    .ZN(_10487_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14864_ (.I(_10432_[0]),
    .ZN(_10497_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14865_ (.I(_10434_[0]),
    .ZN(_10500_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14866_ (.I(_10456_[0]),
    .ZN(_10525_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14867_ (.I(_10476_[0]),
    .ZN(_10536_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14868_ (.I(_10494_[0]),
    .ZN(_10548_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14869_ (.I(_10511_[0]),
    .ZN(_10577_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14870_ (.I(_10531_[0]),
    .ZN(_10588_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14871_ (.I(_10540_[0]),
    .ZN(_10594_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14872_ (.I(_10542_[0]),
    .ZN(_10605_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14873_ (.I(_10546_[0]),
    .ZN(_10601_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14874_ (.I(_10563_[0]),
    .ZN(_10630_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14875_ (.I(_10583_[0]),
    .ZN(_10641_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14876_ (.I(_10599_[0]),
    .ZN(_10649_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14877_ (.I(_10616_[0]),
    .ZN(_10680_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14878_ (.I(_10636_[0]),
    .ZN(_10691_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14879_ (.I(_10647_[0]),
    .ZN(_10699_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14880_ (.I(_10654_[0]),
    .ZN(_10719_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14881_ (.I(_10659_[0]),
    .ZN(_10712_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14882_ (.I(_10664_[0]),
    .ZN(_10727_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14883_ (.I(_10686_[0]),
    .ZN(_10738_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14884_ (.I(_10705_[0]),
    .ZN(_10757_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14885_ (.I(_10710_[0]),
    .ZN(_10771_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14886_ (.I(_10733_[0]),
    .ZN(_10782_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14887_ (.I(_10746_[0]),
    .ZN(_10803_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14888_ (.I(_10749_[0]),
    .ZN(_10798_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14889_ (.I(_10754_[0]),
    .ZN(_10812_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14890_ (.I(_10777_[0]),
    .ZN(_10823_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14891_ (.I(_10790_[0]),
    .ZN(_10842_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14892_ (.I(_10795_[0]),
    .ZN(_10851_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14893_ (.I(_10818_[0]),
    .ZN(_10862_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14894_ (.I(_10831_[0]),
    .ZN(_10880_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14895_ (.I(_10835_[0]),
    .ZN(_10889_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14896_ (.I(_10857_[0]),
    .ZN(_10900_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14897_ (.I(_10866_[0]),
    .ZN(_10906_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14898_ (.I(_10868_[0]),
    .ZN(_10910_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14899_ (.I(_10873_[0]),
    .ZN(_10925_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14900_ (.I(_10895_[0]),
    .ZN(_10937_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14901_ (.I(_10904_[0]),
    .ZN(_10943_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14902_ (.I(_10917_[0]),
    .ZN(_10965_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14903_ (.I(_10922_[0]),
    .ZN(_10955_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14904_ (.I(_10931_[0]),
    .ZN(_10968_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14905_ (.I(_10941_[0]),
    .ZN(_10974_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14906_ (.I(_10962_[0]),
    .ZN(_10994_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3165 (.I(_04304_),
    .Z(net3165));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3166 (.I(_04298_),
    .Z(net3166));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14909_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[1] ),
    .B2(_07029_),
    .ZN(_08756_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3167 (.I(_04293_),
    .Z(net3167));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14911_ (.A1(net276),
    .A2(_07031_),
    .ZN(_08758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14912_ (.A1(net3655),
    .A2(_06935_),
    .B(_08756_),
    .C(_08758_),
    .ZN(_08759_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3170 (.I(_04271_),
    .Z(net3170));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3169 (.I(_04281_),
    .Z(net3169));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14915_ (.I0(net3196),
    .I1(_07013_),
    .S(_06440_),
    .Z(_08762_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14916_ (.A1(net3374),
    .A2(_08759_),
    .B(_08762_),
    .ZN(_11018_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14917_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[2] ),
    .B2(_07029_),
    .ZN(_08763_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14918_ (.A1(net557),
    .A2(_07031_),
    .ZN(_08764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14919_ (.A1(net3655),
    .A2(_07061_),
    .B(_08763_),
    .C(_08764_),
    .ZN(_08765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14920_ (.I0(net3196),
    .I1(net267),
    .S(_11410_[0]),
    .Z(_08766_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14921_ (.A1(net3374),
    .A2(_08765_),
    .B(_08766_),
    .ZN(_11022_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14922_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[3] ),
    .B2(_07029_),
    .ZN(_08767_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14923_ (.A1(net436),
    .A2(_07031_),
    .ZN(_08768_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14924_ (.A1(net3655),
    .A2(_07088_),
    .B(_08767_),
    .C(_08768_),
    .ZN(_08769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14925_ (.I0(net3196),
    .I1(net267),
    .S(_11418_[0]),
    .Z(_08770_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14926_ (.A1(net3374),
    .A2(_08769_),
    .B(_08770_),
    .ZN(_11026_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3168 (.I(_04288_),
    .Z(net3168));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14928_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[4] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net331),
    .ZN(_08772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14929_ (.A1(net3655),
    .A2(_07106_),
    .B(_08772_),
    .ZN(_08773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14930_ (.I0(net3196),
    .I1(_07013_),
    .S(_06530_),
    .Z(_08774_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14931_ (.A1(net3374),
    .A2(_08773_),
    .B(_08774_),
    .ZN(_11030_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14932_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[5] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net341),
    .ZN(_08775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14933_ (.A1(net3655),
    .A2(net3367),
    .B(_08775_),
    .ZN(_08776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14934_ (.I0(net3196),
    .I1(_07013_),
    .S(_11434_[0]),
    .Z(_08777_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14935_ (.A1(net3374),
    .A2(_08776_),
    .B(_08777_),
    .ZN(_11034_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14936_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[6] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net428),
    .ZN(_08778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14937_ (.A1(net3655),
    .A2(net3366),
    .B(_08778_),
    .ZN(_08779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14938_ (.I0(net3196),
    .I1(net267),
    .S(_11442_[0]),
    .Z(_08780_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14939_ (.A1(net3374),
    .A2(_08779_),
    .B(_08780_),
    .ZN(_11038_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14940_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[7] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net426),
    .ZN(_08781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14941_ (.A1(net3655),
    .A2(net3365),
    .B(_08781_),
    .ZN(_08782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14942_ (.I0(net3196),
    .I1(_07013_),
    .S(_11450_[0]),
    .Z(_08783_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14943_ (.A1(net3374),
    .A2(_08782_),
    .B(_08783_),
    .ZN(_11042_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14944_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[8] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net412),
    .ZN(_08784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14945_ (.A1(net3655),
    .A2(net3364),
    .B(_08784_),
    .ZN(_08785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14946_ (.I0(net3196),
    .I1(net267),
    .S(_11458_[0]),
    .Z(_08786_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14947_ (.A1(net3374),
    .A2(_08785_),
    .B(_08786_),
    .ZN(_11046_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3171 (.I(_04240_),
    .Z(net3171));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14949_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[9] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net408),
    .ZN(_08788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14950_ (.A1(net3655),
    .A2(net3363),
    .B(_08788_),
    .ZN(_08789_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3188 (.I(_02690_),
    .Z(net3188));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14952_ (.I0(net3196),
    .I1(_07013_),
    .S(_11466_[0]),
    .Z(_08791_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14953_ (.A1(net3374),
    .A2(_08789_),
    .B(_08791_),
    .ZN(_11050_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14954_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[10] ),
    .B2(_07029_),
    .ZN(_08792_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14955_ (.A1(net425),
    .A2(_07031_),
    .ZN(_08793_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14956_ (.A1(net3655),
    .A2(net3362),
    .B(_08792_),
    .C(_08793_),
    .ZN(_08794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14957_ (.I0(net3196),
    .I1(_07013_),
    .S(_11474_[0]),
    .Z(_08795_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14958_ (.A1(net3374),
    .A2(_08794_),
    .B(_08795_),
    .ZN(_11054_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3172 (.I(_04236_),
    .Z(net3172));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3173 (.I(_04232_),
    .Z(net3173));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14961_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[11] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net422),
    .ZN(_08798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14962_ (.A1(net3655),
    .A2(net3377),
    .B(_08798_),
    .ZN(_08799_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3175 (.I(_04221_),
    .Z(net3175));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14964_ (.I0(net305),
    .I1(net267),
    .S(_11482_[0]),
    .Z(_08801_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14965_ (.A1(net3374),
    .A2(_08799_),
    .B(_08801_),
    .ZN(_11058_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14966_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[12] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net420),
    .ZN(_08802_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14967_ (.A1(net3655),
    .A2(net3381),
    .B(_08802_),
    .ZN(_08803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14968_ (.I0(net3197),
    .I1(net309),
    .S(_11493_[0]),
    .Z(_08804_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14969_ (.A1(net3374),
    .A2(_08803_),
    .B(_08804_),
    .ZN(_11062_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14970_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[13] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net424),
    .ZN(_08805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14971_ (.A1(net3655),
    .A2(_07369_),
    .B(_08805_),
    .ZN(_08806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14972_ (.I0(net3196),
    .I1(net3195),
    .S(_11501_[0]),
    .Z(_08807_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14973_ (.A1(net3374),
    .A2(_08806_),
    .B(_08807_),
    .ZN(_11066_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3176 (.I(_04216_),
    .Z(net3176));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14975_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[14] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_07449_),
    .ZN(_08809_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14976_ (.A1(net3655),
    .A2(net3351),
    .B(_08809_),
    .ZN(_08810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14977_ (.I0(net3196),
    .I1(net3195),
    .S(_11509_[0]),
    .Z(_08811_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14978_ (.A1(net3374),
    .A2(_08810_),
    .B(_08811_),
    .ZN(_11070_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _14979_ (.I(net3350),
    .ZN(_08812_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3177 (.I(_04210_),
    .Z(net3177));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14981_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[15] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_07486_),
    .ZN(_08814_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14982_ (.A1(net3655),
    .A2(_08812_),
    .B(_08814_),
    .ZN(_08815_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14983_ (.I0(net305),
    .I1(net3195),
    .S(_11517_[0]),
    .Z(_08816_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14984_ (.A1(net3374),
    .A2(_08815_),
    .B(_08816_),
    .ZN(_11074_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14985_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[16] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_07544_),
    .ZN(_08817_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14986_ (.A1(net3655),
    .A2(_07526_),
    .B(_08817_),
    .ZN(_08818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14987_ (.I0(net305),
    .I1(net3195),
    .S(_11525_[0]),
    .Z(_08819_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14988_ (.A1(net3374),
    .A2(_08818_),
    .B(_08819_),
    .ZN(_11078_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14989_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[17] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_07582_),
    .ZN(_08820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14990_ (.A1(net3655),
    .A2(net3349),
    .B(_08820_),
    .ZN(_08821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14991_ (.I0(net3197),
    .I1(net282),
    .S(_11533_[0]),
    .Z(_08822_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14992_ (.A1(net3374),
    .A2(_08821_),
    .B(_08822_),
    .ZN(_11082_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14993_ (.I(net3359),
    .ZN(_08823_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14994_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[18] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net414),
    .ZN(_08824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14995_ (.A1(net3655),
    .A2(_08823_),
    .B(_08824_),
    .ZN(_08825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14996_ (.I0(net3197),
    .I1(net282),
    .S(_11541_[0]),
    .Z(_08826_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14997_ (.A1(net3375),
    .A2(_08825_),
    .B(_08826_),
    .ZN(_11086_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14998_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[19] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net441),
    .ZN(_08827_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14999_ (.A1(net3655),
    .A2(net3348),
    .B(_08827_),
    .ZN(_08828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15000_ (.I0(net305),
    .I1(net282),
    .S(_11549_[0]),
    .Z(_08829_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15001_ (.A1(net3374),
    .A2(_08828_),
    .B(_08829_),
    .ZN(_11090_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3183 (.I(_04030_),
    .Z(net3183));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15003_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[20] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net410),
    .ZN(_08831_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15004_ (.A1(net3655),
    .A2(_07712_),
    .B(_08831_),
    .ZN(_08832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15005_ (.I0(net309),
    .I1(net305),
    .S(_11553_[0]),
    .Z(_08833_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15006_ (.A1(net3374),
    .A2(_08832_),
    .B(_08833_),
    .ZN(_11094_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3192 (.I(_02529_),
    .Z(net3192));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3447 (.I(net3446),
    .Z(net3447));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15009_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[21] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net442),
    .ZN(_08836_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15010_ (.A1(net3655),
    .A2(net3347),
    .B(_08836_),
    .ZN(_08837_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3178 (.I(_04156_),
    .Z(net3178));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15012_ (.I0(net309),
    .I1(net305),
    .S(_11561_[0]),
    .Z(_08839_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15013_ (.A1(net3374),
    .A2(_08837_),
    .B(_08839_),
    .ZN(_11098_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15014_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[22] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_07838_),
    .ZN(_08840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15015_ (.A1(net3655),
    .A2(net3346),
    .B(_08840_),
    .ZN(_08841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15016_ (.I0(net282),
    .I1(net3197),
    .S(_11569_[0]),
    .Z(_08842_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15017_ (.A1(net3375),
    .A2(_08841_),
    .B(_08842_),
    .ZN(_11102_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15018_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[23] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_07875_),
    .ZN(_08843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15019_ (.A1(net3655),
    .A2(net3345),
    .B(_08843_),
    .ZN(_08844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15020_ (.I0(net282),
    .I1(net305),
    .S(_11577_[0]),
    .Z(_08845_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15021_ (.A1(net3375),
    .A2(_08844_),
    .B(_08845_),
    .ZN(_11106_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15022_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[24] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_07936_),
    .ZN(_08846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15023_ (.A1(net3655),
    .A2(net3344),
    .B(_08846_),
    .ZN(_08847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15024_ (.I0(net3195),
    .I1(net305),
    .S(_11585_[0]),
    .Z(_08848_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15025_ (.A1(net3375),
    .A2(_08847_),
    .B(_08848_),
    .ZN(_11110_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15026_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[25] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_07973_),
    .ZN(_08849_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15027_ (.A1(net3655),
    .A2(net3343),
    .B(_08849_),
    .ZN(_08850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15028_ (.I0(net309),
    .I1(net3197),
    .S(_11593_[0]),
    .Z(_08851_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15029_ (.A1(net3375),
    .A2(_08850_),
    .B(_08851_),
    .ZN(_11114_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15030_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[26] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_08017_),
    .ZN(_08852_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15031_ (.A1(net3655),
    .A2(net3342),
    .B(_08852_),
    .ZN(_08853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15032_ (.I0(net282),
    .I1(net3197),
    .S(_11601_[0]),
    .Z(_08854_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15033_ (.A1(net3375),
    .A2(_08853_),
    .B(_08854_),
    .ZN(_11118_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15034_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[27] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_08055_),
    .ZN(_08855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15035_ (.A1(net3655),
    .A2(net3357),
    .B(_08855_),
    .ZN(_08856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15036_ (.I0(net282),
    .I1(net3197),
    .S(_11609_[0]),
    .Z(_08857_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15037_ (.A1(net3375),
    .A2(_08856_),
    .B(_08857_),
    .ZN(_11122_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15038_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[28] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(net530),
    .ZN(_08858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15039_ (.A1(net3655),
    .A2(net3341),
    .B(_08858_),
    .ZN(_08859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15040_ (.I0(net282),
    .I1(net3197),
    .S(_11617_[0]),
    .Z(_08860_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15041_ (.A1(net3374),
    .A2(_08859_),
    .B(_08860_),
    .ZN(_11126_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15042_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[29] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_08145_),
    .ZN(_08861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15043_ (.A1(net3655),
    .A2(net3340),
    .B(_08861_),
    .ZN(_08862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15044_ (.I0(net282),
    .I1(net3197),
    .S(_11625_[0]),
    .Z(_08863_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15045_ (.A1(net3375),
    .A2(_08862_),
    .B(_08863_),
    .ZN(_11130_[0]));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15046_ (.A1(_07027_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[30] ),
    .B2(_07029_),
    .C1(_07031_),
    .C2(_08193_),
    .ZN(_08864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15047_ (.A1(net3655),
    .A2(net3339),
    .B(_08864_),
    .ZN(_08865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15048_ (.I0(net282),
    .I1(net3197),
    .S(_11633_[0]),
    .Z(_08866_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15049_ (.A1(net3375),
    .A2(_08865_),
    .B(_08866_),
    .ZN(_11134_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _15050_ (.I(_06849_),
    .ZN(_11146_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3451 (.I(net3450),
    .Z(net3451));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _15052_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .ZN(_11169_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15053_ (.I(_09758_[0]),
    .ZN(_09759_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15054_ (.A1(net3334),
    .A2(net3328),
    .Z(_11190_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15055_ (.I(_09770_[0]),
    .ZN(_09786_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15056_ (.A1(net3334),
    .A2(net3318),
    .Z(_11202_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15057_ (.I(_09804_[0]),
    .ZN(_11204_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15058_ (.A1(net3334),
    .A2(net3299),
    .Z(_11211_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15059_ (.I(_09803_[0]),
    .ZN(_09822_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15060_ (.I(_09843_[0]),
    .ZN(_09845_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15061_ (.I(_09819_[0]),
    .ZN(_09852_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15062_ (.I(_09878_[0]),
    .ZN(_09880_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15063_ (.I(_09842_[0]),
    .ZN(_09879_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15064_ (.A1(net3334),
    .A2(net3314),
    .Z(_11228_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15065_ (.I(_09906_[0]),
    .ZN(_09908_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15066_ (.I(_09877_[0]),
    .ZN(_09907_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15067_ (.A1(net3334),
    .A2(net3295),
    .Z(_11237_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15068_ (.I(_09887_[0]),
    .ZN(_09918_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15069_ (.I(_09915_[0]),
    .ZN(_09954_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15070_ (.I(_09948_[0]),
    .ZN(_09987_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15071_ (.I(_09951_[0]),
    .ZN(_09999_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15072_ (.A1(net3333),
    .A2(net3238),
    .Z(_11257_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15073_ (.I(_10077_[0]),
    .ZN(_10079_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15074_ (.I(_10032_[0]),
    .ZN(_10078_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15075_ (.I(_10040_[0]),
    .ZN(_11268_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15076_ (.I(_10123_[0]),
    .ZN(_10125_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15077_ (.I(_10076_[0]),
    .ZN(_10124_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15078_ (.A1(net3333),
    .A2(net3301),
    .Z(_11274_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15079_ (.I(_10087_[0]),
    .ZN(_10136_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15080_ (.A1(net3333),
    .A2(net3293),
    .Z(_11280_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15081_ (.I(_10133_[0]),
    .ZN(_10183_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15082_ (.I(_08616_),
    .ZN(_10188_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15083_ (.I(_10232_[0]),
    .ZN(_10234_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15084_ (.I(_10175_[0]),
    .ZN(_10242_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15085_ (.I(_10180_[0]),
    .ZN(_10251_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15086_ (.I(_10302_[0]),
    .ZN(_11296_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15087_ (.I(_10292_[0]),
    .ZN(_10360_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15088_ (.I(_10310_[0]),
    .ZN(_11298_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15089_ (.I(_10358_[0]),
    .ZN(_11302_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15090_ (.I(_10368_[0]),
    .ZN(_11304_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15091_ (.I(_10415_[0]),
    .ZN(_11308_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15092_ (.I(_10426_[0]),
    .ZN(_11310_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15093_ (.I(_10471_[0]),
    .ZN(_11314_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15094_ (.I(_10482_[0]),
    .ZN(_11316_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15095_ (.I(_10526_[0]),
    .ZN(_11320_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15096_ (.I(_10537_[0]),
    .ZN(_11322_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15097_ (.I(_10578_[0]),
    .ZN(_11326_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15098_ (.I(_10589_[0]),
    .ZN(_11328_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15099_ (.I(_10596_[0]),
    .ZN(_10653_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15100_ (.I(_10631_[0]),
    .ZN(_11332_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15101_ (.I(_10642_[0]),
    .ZN(_11334_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15102_ (.I(_10681_[0]),
    .ZN(_11338_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15103_ (.I(_10692_[0]),
    .ZN(_11340_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15104_ (.I(_10728_[0]),
    .ZN(_11344_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15105_ (.I(_10739_[0]),
    .ZN(_11346_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15106_ (.I(_10772_[0]),
    .ZN(_11350_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15107_ (.I(_10783_[0]),
    .ZN(_11352_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15108_ (.I(_10651_[0]),
    .ZN(_10652_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15109_ (.I(_10813_[0]),
    .ZN(_11356_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15110_ (.I(_10824_[0]),
    .ZN(_11358_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15111_ (.I(_10852_[0]),
    .ZN(_11362_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15112_ (.I(_10863_[0]),
    .ZN(_11364_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15113_ (.I(_10890_[0]),
    .ZN(_11368_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15114_ (.I(_10901_[0]),
    .ZN(_11370_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15115_ (.I(_10926_[0]),
    .ZN(_11374_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15116_ (.I(_10938_[0]),
    .ZN(_11376_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15117_ (.I(_10957_[0]),
    .ZN(_11382_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15118_ (.I(_10969_[0]),
    .ZN(_11384_[0]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15119_ (.A1(_11458_[0]),
    .A2(_06783_),
    .ZN(_11160_[0]));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _15120_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .ZN(_11170_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15121_ (.I(_09753_[0]),
    .ZN(_11185_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15122_ (.I(_09752_[0]),
    .ZN(_09761_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15123_ (.A1(net529),
    .A2(net3285),
    .Z(_11191_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15124_ (.I(_09771_[0]),
    .ZN(_11193_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15125_ (.I(_09784_[0]),
    .ZN(_09787_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15126_ (.A1(net3285),
    .A2(net3318),
    .Z(_11212_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15127_ (.I(_09820_[0]),
    .ZN(_09823_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15128_ (.I(_09850_[0]),
    .ZN(_09853_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15129_ (.I(_09888_[0]),
    .ZN(_11230_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15130_ (.A1(net3285),
    .A2(net3314),
    .Z(_11238_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15131_ (.I(_09916_[0]),
    .ZN(_09919_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15132_ (.I(_09949_[0]),
    .ZN(_11246_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15133_ (.I(_09952_[0]),
    .ZN(_09955_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15134_ (.I(_09985_[0]),
    .ZN(_09988_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15135_ (.I(_09941_[0]),
    .ZN(_09992_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15136_ (.I(_09997_[0]),
    .ZN(_10000_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15137_ (.A1(net3284),
    .A2(net3313),
    .Z(_11258_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15138_ (.I(_10041_[0]),
    .ZN(_11261_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15139_ (.I(_10022_[0]),
    .ZN(_10080_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15140_ (.I(_10035_[0]),
    .ZN(_11266_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15141_ (.I(_10088_[0]),
    .ZN(_11269_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15142_ (.I(_10061_[0]),
    .ZN(_10126_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15143_ (.I(_10134_[0]),
    .ZN(_10137_[0]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15144_ (.A1(net3284),
    .A2(net3301),
    .Z(_11281_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15145_ (.I(_10181_[0]),
    .ZN(_10184_[0]));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15146_ (.A1(net3657),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .B1(_08583_),
    .B2(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .ZN(_08868_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15147_ (.I(_08868_),
    .ZN(_10189_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15148_ (.I(_10241_[0]),
    .ZN(_10244_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15149_ (.I(_10249_[0]),
    .ZN(_10252_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15150_ (.I(_10303_[0]),
    .ZN(_11291_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15151_ (.I(_10311_[0]),
    .ZN(_11293_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15152_ (.I(_10359_[0]),
    .ZN(_11297_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15153_ (.I(_10369_[0]),
    .ZN(_11299_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15154_ (.I(_10416_[0]),
    .ZN(_11303_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15155_ (.I(_10348_[0]),
    .ZN(_10419_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15156_ (.I(_10427_[0]),
    .ZN(_11305_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15157_ (.I(_10472_[0]),
    .ZN(_11309_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15158_ (.I(_10405_[0]),
    .ZN(_10475_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15159_ (.I(_10483_[0]),
    .ZN(_11311_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15160_ (.I(_10527_[0]),
    .ZN(_11315_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15161_ (.I(_10461_[0]),
    .ZN(_10530_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15162_ (.I(_10538_[0]),
    .ZN(_11317_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15163_ (.I(_10579_[0]),
    .ZN(_11321_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15164_ (.I(_10516_[0]),
    .ZN(_10582_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15165_ (.I(_10590_[0]),
    .ZN(_11323_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15166_ (.I(_10632_[0]),
    .ZN(_11327_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15167_ (.I(_10568_[0]),
    .ZN(_10635_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15168_ (.I(_10643_[0]),
    .ZN(_11329_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15169_ (.I(_10682_[0]),
    .ZN(_11333_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15170_ (.I(_10621_[0]),
    .ZN(_10685_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15171_ (.I(_10693_[0]),
    .ZN(_11335_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15172_ (.I(_10729_[0]),
    .ZN(_11339_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15173_ (.I(_10670_[0]),
    .ZN(_10732_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15174_ (.I(_10740_[0]),
    .ZN(_11341_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15175_ (.I(_10773_[0]),
    .ZN(_11345_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15176_ (.I(_10717_[0]),
    .ZN(_10775_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15177_ (.I(_10784_[0]),
    .ZN(_11347_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15178_ (.I(_10814_[0]),
    .ZN(_11351_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15179_ (.I(_10761_[0]),
    .ZN(_10817_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15180_ (.I(_10825_[0]),
    .ZN(_11353_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15181_ (.I(_10853_[0]),
    .ZN(_11357_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15182_ (.I(_10801_[0]),
    .ZN(_10856_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15183_ (.I(_10864_[0]),
    .ZN(_11359_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15184_ (.I(_10891_[0]),
    .ZN(_11363_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15185_ (.I(_10840_[0]),
    .ZN(_10894_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15186_ (.I(_10902_[0]),
    .ZN(_11365_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15187_ (.I(_10912_[0]),
    .ZN(_10916_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15188_ (.I(_10927_[0]),
    .ZN(_11369_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15189_ (.I(_10878_[0]),
    .ZN(_10930_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15190_ (.I(_10939_[0]),
    .ZN(_11371_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15191_ (.I(_10958_[0]),
    .ZN(_11375_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15192_ (.I(_10913_[0]),
    .ZN(_10961_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15193_ (.I(_10970_[0]),
    .ZN(_11377_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15194_ (.I(_10996_[0]),
    .ZN(_11385_[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3179 (.I(_04151_),
    .Z(net3179));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 _15196_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .ZN(_08869_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15197_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .ZN(_08870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15198_ (.A1(_08360_),
    .A2(_08658_),
    .ZN(_08871_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15199_ (.A1(_08389_),
    .A2(_08361_),
    .Z(_08872_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15200_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_08658_),
    .B1(_08871_),
    .B2(_08872_),
    .ZN(_08873_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3450 (.I(_06334_),
    .Z(net3450));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3180 (.I(_04133_),
    .Z(net3180));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15203_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .B(_08676_),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .ZN(_08876_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15204_ (.A1(_08870_),
    .A2(_08873_),
    .A3(_08876_),
    .Z(_08877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15205_ (.A1(_08869_),
    .A2(_08877_),
    .ZN(_08878_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _15206_ (.I(_08878_),
    .ZN(_11661_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15207_ (.I(_11215_[0]),
    .ZN(_09818_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15208_ (.I(_11225_[0]),
    .ZN(_09858_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15209_ (.I(_11241_[0]),
    .ZN(_09914_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15210_ (.I(_11248_[0]),
    .ZN(_09950_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15211_ (.I(_11267_[0]),
    .ZN(_10086_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15212_ (.I(_11277_[0]),
    .ZN(_10132_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15213_ (.I(_11286_[0]),
    .ZN(_10179_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15214_ (.I(_11192_[0]),
    .ZN(_09769_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15215_ (.I(_11203_[0]),
    .ZN(_09802_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15216_ (.I(_11229_[0]),
    .ZN(_09886_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15217_ (.I(_11260_[0]),
    .ZN(_10031_[0]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15218_ (.I(_11292_[0]),
    .ZN(_10304_[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15219_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .S(_08470_),
    .Z(_00007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15220_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .I1(net3659),
    .S(_08470_),
    .Z(_00008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3449 (.I(net3448),
    .Z(net3449));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15222_ (.I0(net3658),
    .I1(net3656),
    .S(_08407_),
    .Z(_00009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15223_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .I1(net3655),
    .S(_08407_),
    .Z(_00010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15224_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .S(_08407_),
    .Z(_00011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15225_ (.A1(_06317_),
    .A2(_06757_),
    .Z(_08880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15226_ (.A1(_06761_),
    .A2(_08880_),
    .Z(_08881_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3181 (.I(_04122_),
    .Z(net3181));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15228_ (.A1(_06953_),
    .A2(_08880_),
    .A3(_08405_),
    .Z(_08883_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15229_ (.A1(_06340_),
    .A2(_08883_),
    .Z(_08884_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15230_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_08884_),
    .Z(_08885_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15231_ (.A1(_06232_),
    .A2(net26),
    .Z(_08886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15232_ (.A1(_08885_),
    .A2(_08886_),
    .ZN(_08887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15233_ (.I0(_08881_),
    .I1(\load_store_unit_i.data_type_q[2] ),
    .S(_08887_),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _15234_ (.A1(_06746_),
    .A2(_06758_),
    .ZN(_08888_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3446 (.I(_06334_),
    .Z(net3446));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15236_ (.I0(_08888_),
    .I1(\load_store_unit_i.data_type_q[1] ),
    .S(_08887_),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15237_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11395_[0]),
    .Z(_08890_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15238_ (.A1(_11148_[0]),
    .A2(_08890_),
    .Z(_08891_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _15239_ (.A1(_08354_),
    .A2(_08355_),
    .ZN(_08892_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15240_ (.A1(_08892_),
    .A2(_08328_),
    .Z(_08893_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3182 (.I(_04115_),
    .Z(net3182));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15242_ (.A1(_06783_),
    .A2(_08327_),
    .ZN(_08895_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _15243_ (.A1(_06530_),
    .A2(_08299_),
    .A3(_08303_),
    .ZN(_08896_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15244_ (.A1(net485),
    .A2(_08349_),
    .Z(_08897_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15245_ (.A1(_08895_),
    .A2(_08896_),
    .A3(_08897_),
    .Z(_08898_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15246_ (.A1(_08328_),
    .A2(_08896_),
    .Z(_08899_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3205 (.I(_10650_[0]),
    .Z(net3205));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15248_ (.A1(\cs_registers_i.dcsr_q[0] ),
    .A2(_08893_),
    .B1(_08898_),
    .B2(\cs_registers_i.mcause_q[0] ),
    .C1(_08899_),
    .C2(\cs_registers_i.mscratch_q[0] ),
    .ZN(_08901_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3184 (.I(_03629_),
    .Z(net3184));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3200 (.I(_08912_),
    .Z(net3200));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3189 (.I(_02593_),
    .Z(net3189));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15252_ (.A1(_06530_),
    .A2(_06783_),
    .ZN(_08905_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15253_ (.A1(_08895_),
    .A2(_08905_),
    .Z(_08906_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3197 (.I(net3196),
    .Z(net3197));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15255_ (.I(\cs_registers_i.mhpmcounter[1888] ),
    .ZN(_08908_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _15256_ (.A1(net301),
    .A2(net485),
    .A3(_06530_),
    .A4(_08327_),
    .Z(_08909_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _15257_ (.A1(_08336_),
    .A2(_08340_),
    .A3(_08909_),
    .ZN(_08910_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3186 (.I(_11073_[0]),
    .Z(net3186));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _15259_ (.A1(_06530_),
    .A2(_08333_),
    .B(_08340_),
    .C(_08280_),
    .ZN(_08912_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3187 (.I(_11065_[0]),
    .Z(net3187));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15261_ (.I(\cs_registers_i.mhpmcounter[1856] ),
    .ZN(_08914_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15262_ (.A1(_08908_),
    .A2(_08910_),
    .B1(_08912_),
    .B2(_08914_),
    .ZN(_08915_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15263_ (.A1(_08897_),
    .A2(_08906_),
    .A3(_08915_),
    .ZN(_08916_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15264_ (.A1(_08905_),
    .A2(_08328_),
    .Z(_08917_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _15265_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .ZN(_08918_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15266_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .ZN(_08919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15267_ (.A1(_08286_),
    .A2(_08345_),
    .ZN(_08920_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15268_ (.A1(_08342_),
    .A2(_08920_),
    .Z(_08921_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _15269_ (.A1(_08918_),
    .A2(_08910_),
    .B1(_08912_),
    .B2(_08919_),
    .C(_08921_),
    .ZN(_08922_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15270_ (.A1(_08917_),
    .A2(_08922_),
    .ZN(_08923_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15271_ (.A1(_11434_[0]),
    .A2(_08331_),
    .A3(_08328_),
    .Z(_08924_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3193 (.I(_02515_),
    .Z(net3193));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15273_ (.A1(_08274_),
    .A2(_08348_),
    .A3(_08287_),
    .Z(_08926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15274_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_08924_),
    .B(_08926_),
    .ZN(_08927_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15275_ (.A1(_08356_),
    .A2(_08897_),
    .Z(_08928_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3196 (.I(_07009_),
    .Z(net3196));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15277_ (.A1(_11414_[0]),
    .A2(net3288),
    .Z(_08930_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15278_ (.A1(_06388_),
    .A2(net263),
    .A3(_06783_),
    .A4(_08930_),
    .Z(_08931_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15279_ (.A1(_08931_),
    .A2(_08896_),
    .Z(_08932_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3198 (.I(_05562_),
    .Z(net3198));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15281_ (.A1(\cs_registers_i.dscratch0_q[0] ),
    .A2(net3199),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[0] ),
    .ZN(_08934_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15282_ (.A1(_08350_),
    .A2(_08353_),
    .Z(_08935_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3209 (.I(_08959_),
    .Z(net3209));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15284_ (.A1(_06388_),
    .A2(net485),
    .A3(_06783_),
    .A4(_08930_),
    .Z(_08937_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15285_ (.A1(_08896_),
    .A2(_08937_),
    .Z(_08938_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3206 (.I(_03181_),
    .Z(net3206));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15287_ (.A1(_08892_),
    .A2(_08937_),
    .Z(_08940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15288_ (.A1(net62),
    .A2(_08935_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[0] ),
    .C1(\cs_registers_i.dscratch1_q[0] ),
    .C2(_08940_),
    .ZN(_08941_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15289_ (.A1(_08927_),
    .A2(_08934_),
    .A3(_08941_),
    .Z(_08942_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15290_ (.A1(_08901_),
    .A2(_08916_),
    .A3(_08923_),
    .A4(_08942_),
    .Z(_08943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15291_ (.A1(_11399_[0]),
    .A2(_08943_),
    .ZN(_08944_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15292_ (.A1(_08891_),
    .A2(_08944_),
    .Z(_08945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15293_ (.A1(_08326_),
    .A2(_08358_),
    .ZN(_08946_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3213 (.I(_10602_[0]),
    .Z(net3213));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15295_ (.I(_11154_[0]),
    .ZN(_08948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15296_ (.A1(_06783_),
    .A2(_08404_),
    .Z(_08949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15297_ (.A1(_08370_),
    .A2(_08356_),
    .B(_08369_),
    .ZN(_08950_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15298_ (.A1(_08948_),
    .A2(_08359_),
    .A3(_08949_),
    .A4(_08950_),
    .Z(_08951_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3237 (.I(net3236),
    .Z(net3237));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15300_ (.A1(_08946_),
    .A2(_08924_),
    .A3(_08951_),
    .ZN(_08953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15301_ (.I0(_08945_),
    .I1(\cs_registers_i.mcountinhibit_q[0] ),
    .S(_08953_),
    .Z(_00014_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3239 (.I(net3238),
    .Z(net3239));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15303_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11409_[0]),
    .Z(_08955_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15304_ (.A1(_11148_[0]),
    .A2(_08955_),
    .Z(_08956_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3448 (.I(_06334_),
    .Z(net3448));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3249 (.I(_08513_),
    .Z(net3249));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _15307_ (.A1(_06388_),
    .A2(net485),
    .B(_06783_),
    .ZN(_08959_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3262 (.I(_08575_),
    .Z(net3262));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15309_ (.A1(\cs_registers_i.mhpmcounter[1858] ),
    .A2(_08897_),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .ZN(_08961_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15310_ (.A1(_08912_),
    .A2(_08961_),
    .ZN(_08962_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15311_ (.A1(_08336_),
    .A2(_08340_),
    .A3(_08909_),
    .Z(_08963_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3281 (.I(net3280),
    .Z(net3281));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15313_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A2(_08963_),
    .A3(_08959_),
    .Z(_08965_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15314_ (.I(\cs_registers_i.mhpmcounter[1890] ),
    .ZN(_08966_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3432 (.I(net3427),
    .Z(net3432));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15316_ (.A1(_08966_),
    .A2(_08910_),
    .B(_08921_),
    .ZN(_08968_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15317_ (.A1(_08897_),
    .A2(_08968_),
    .Z(_08969_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _15318_ (.A1(_08962_),
    .A2(_08965_),
    .A3(_08969_),
    .B(_08906_),
    .ZN(_08970_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15319_ (.A1(\cs_registers_i.csr_mepc_o[2] ),
    .A2(_08896_),
    .Z(_08971_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15320_ (.A1(_08287_),
    .A2(_08971_),
    .Z(_08972_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15321_ (.A1(\cs_registers_i.mcountinhibit_q[2] ),
    .A2(_08924_),
    .B1(_08972_),
    .B2(_08931_),
    .ZN(_08973_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3278 (.I(_08524_),
    .Z(net3278));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15323_ (.A1(\cs_registers_i.mcause_q[2] ),
    .A2(_08898_),
    .B1(_08899_),
    .B2(\cs_registers_i.mscratch_q[2] ),
    .C1(_08938_),
    .C2(\cs_registers_i.mtval_q[2] ),
    .ZN(_08975_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3288 (.I(_11422_[0]),
    .Z(net3288));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15325_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_08328_),
    .ZN(_08977_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15326_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(_08931_),
    .B1(_08937_),
    .B2(\cs_registers_i.dscratch1_q[2] ),
    .ZN(_08978_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15327_ (.A1(_08977_),
    .A2(_08978_),
    .ZN(_08979_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3299 (.I(net3298),
    .Z(net3299));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15329_ (.A1(net84),
    .A2(_08935_),
    .B1(_08979_),
    .B2(_08892_),
    .C1(_08928_),
    .C2(\cs_registers_i.dscratch0_q[2] ),
    .ZN(_08981_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15330_ (.A1(_08970_),
    .A2(_08973_),
    .A3(_08975_),
    .A4(_08981_),
    .ZN(_08982_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15331_ (.A1(_11409_[0]),
    .A2(_08982_),
    .Z(_08983_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15332_ (.A1(_08956_),
    .A2(_08983_),
    .Z(_08984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15333_ (.I0(_08984_),
    .I1(\cs_registers_i.mcountinhibit_q[2] ),
    .S(_08953_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15334_ (.A1(_08891_),
    .A2(_08944_),
    .ZN(_08985_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3284 (.I(_08507_),
    .Z(net3284));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15336_ (.A1(net3287),
    .A2(_08931_),
    .ZN(_08987_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15337_ (.A1(_08987_),
    .A2(_08337_),
    .A3(_08340_),
    .Z(_08988_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15338_ (.A1(_08951_),
    .A2(_08917_),
    .Z(_08989_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15339_ (.A1(_08988_),
    .A2(_08989_),
    .Z(_08990_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3305 (.I(net3304),
    .Z(net3305));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15341_ (.A1(_08910_),
    .A2(_08990_),
    .ZN(_08992_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3332 (.I(_08496_),
    .Z(net3332));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3335 (.I(_08484_),
    .Z(net3335));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _15344_ (.I(\cs_registers_i.mcountinhibit_q[0] ),
    .ZN(_08995_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3338 (.I(_08449_),
    .Z(net3338));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15346_ (.A1(_08988_),
    .A2(_08989_),
    .ZN(_08997_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3385 (.I(_06840_),
    .Z(net3385));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15348_ (.A1(_08995_),
    .A2(_08997_),
    .ZN(_08999_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15349_ (.A1(_08963_),
    .A2(_08990_),
    .Z(_09000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15350_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_08997_),
    .B(_09000_),
    .ZN(_09001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15351_ (.I0(_08999_),
    .I1(_09001_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .Z(_09002_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15352_ (.A1(_08985_),
    .A2(_08992_),
    .B(_09002_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15353_ (.A1(_08910_),
    .A2(_08990_),
    .Z(_09003_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3373 (.I(_07020_),
    .Z(net3373));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3399 (.I(_06490_),
    .Z(net3399));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk_i_regs (.I(clknet_6_31__leaf_clk_i_regs),
    .Z(clknet_leaf_7_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_42_clk_i_regs (.I(clknet_6_55__leaf_clk_i_regs),
    .Z(clknet_leaf_42_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_40_clk_i_regs (.I(clknet_6_54__leaf_clk_i_regs),
    .Z(clknet_leaf_40_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3590 (.I(net3589),
    .Z(net3590));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15360_ (.A1(\cs_registers_i.mhpmcounter[1866] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .ZN(_09010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15361_ (.A1(\cs_registers_i.mhpmcounter[1898] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .ZN(_09011_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15362_ (.A1(_08912_),
    .A2(_09010_),
    .B1(_09011_),
    .B2(_08910_),
    .ZN(_09012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15363_ (.A1(\cs_registers_i.csr_mtvec_o[10] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09012_),
    .ZN(_09013_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3589 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .Z(net3589));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3576 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .Z(net3576));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15366_ (.A1(\cs_registers_i.dscratch0_q[10] ),
    .A2(_08928_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[10] ),
    .C1(\cs_registers_i.mscratch_q[10] ),
    .C2(_08899_),
    .ZN(_09016_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3588 (.I(net3583),
    .Z(net3588));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15368_ (.A1(_08892_),
    .A2(_08931_),
    .Z(_09018_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3596 (.I(net3589),
    .Z(net3596));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15370_ (.A1(\cs_registers_i.dscratch1_q[10] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[10] ),
    .C1(net63),
    .C2(_08935_),
    .ZN(_09020_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3580 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .Z(net3580));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15372_ (.A1(\cs_registers_i.mtval_q[10] ),
    .A2(_08938_),
    .B(_08924_),
    .ZN(_09022_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15373_ (.A1(_09013_),
    .A2(_09016_),
    .A3(_09020_),
    .A4(_09022_),
    .Z(_09023_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3595 (.I(net3593),
    .Z(net3595));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3594 (.I(net3593),
    .Z(net3594));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15376_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11473_[0]),
    .Z(_09026_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15377_ (.A1(_11148_[0]),
    .A2(_09026_),
    .ZN(_09027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _15378_ (.A1(_11477_[0]),
    .A2(_09023_),
    .B(_09027_),
    .ZN(_09028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _15379_ (.I(_09028_),
    .ZN(_09029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15380_ (.A1(_08995_),
    .A2(_08997_),
    .Z(_09030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15381_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .A2(_11165_[0]),
    .Z(_09031_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15382_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .Z(_09032_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15383_ (.A1(_09031_),
    .A2(_09032_),
    .Z(_09033_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15384_ (.A1(_09030_),
    .A2(_09033_),
    .Z(_09034_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15385_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .Z(_09035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15386_ (.A1(_09034_),
    .A2(_09035_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .C(_09003_),
    .ZN(_09036_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15387_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .A2(_09034_),
    .A3(_09035_),
    .Z(_09037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15388_ (.A1(_09003_),
    .A2(_09029_),
    .B(_09036_),
    .C(_09037_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3593 (.I(net3589),
    .Z(net3593));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15390_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11481_[0]),
    .Z(_09039_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15391_ (.A1(_11148_[0]),
    .A2(_09039_),
    .Z(_09040_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15392_ (.A1(_08328_),
    .A2(_08287_),
    .Z(_09041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15393_ (.A1(\cs_registers_i.mstatus_q[2] ),
    .A2(_09041_),
    .ZN(_09042_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15394_ (.A1(_08287_),
    .A2(_08350_),
    .Z(_09043_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3592 (.I(net3589),
    .Z(net3592));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3591 (.I(net3589),
    .Z(net3591));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15397_ (.A1(\cs_registers_i.mie_q[15] ),
    .A2(_09043_),
    .ZN(_09046_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place3624 (.I(net3606),
    .Z(net3624));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3623 (.I(net3622),
    .Z(net3623));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3605 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .Z(net3605));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3602 (.I(net3597),
    .Z(net3602));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3604 (.I(net3597),
    .Z(net3604));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15403_ (.A1(\cs_registers_i.dscratch1_q[11] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[11] ),
    .C1(net64),
    .C2(_08935_),
    .ZN(_09052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15404_ (.A1(\cs_registers_i.mhpmcounter[1899] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .ZN(_09053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15405_ (.A1(\cs_registers_i.mhpmcounter[1867] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .ZN(_09054_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15406_ (.A1(_08910_),
    .A2(_09053_),
    .B1(_09054_),
    .B2(_08912_),
    .ZN(_09055_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15407_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09055_),
    .ZN(_09056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15408_ (.A1(\cs_registers_i.dscratch0_q[11] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09057_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15409_ (.A1(\cs_registers_i.dcsr_q[11] ),
    .A2(_08893_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[11] ),
    .C1(_08938_),
    .C2(\cs_registers_i.mtval_q[11] ),
    .ZN(_09058_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3601 (.I(net3597),
    .Z(net3601));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15411_ (.A1(_08896_),
    .A2(_08350_),
    .Z(_09060_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3599 (.I(net3597),
    .Z(net3599));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15413_ (.A1(\cs_registers_i.mscratch_q[11] ),
    .A2(_08899_),
    .B1(_09060_),
    .B2(net129),
    .ZN(_09062_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15414_ (.A1(_09056_),
    .A2(_09057_),
    .A3(_09058_),
    .A4(_09062_),
    .Z(_09063_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15415_ (.A1(_09042_),
    .A2(_09046_),
    .A3(_09052_),
    .A4(_09063_),
    .Z(_09064_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15416_ (.A1(_11485_[0]),
    .A2(_09064_),
    .ZN(_09065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15417_ (.A1(_09040_),
    .A2(_09065_),
    .ZN(_09066_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3164 (.I(_04309_),
    .Z(net3164));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15419_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .A2(_09003_),
    .ZN(_09068_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15420_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(_08995_),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .Z(_09069_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15421_ (.A1(_08997_),
    .A2(_09069_),
    .Z(_09070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15422_ (.A1(_09032_),
    .A2(_09070_),
    .Z(_09071_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15423_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .A2(_09035_),
    .A3(_09071_),
    .Z(_09072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15424_ (.I0(_09068_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .S(_09072_),
    .Z(_09073_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15425_ (.A1(_09003_),
    .A2(_09066_),
    .B(_09073_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15426_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11494_[0]),
    .Z(_09074_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15427_ (.A1(_11148_[0]),
    .A2(_09074_),
    .Z(_09075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3163 (.I(_04314_),
    .Z(net3163));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk_i (.I(clk_i),
    .Z(clknet_0_clk_i));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3174 (.I(_04226_),
    .Z(net3174));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15431_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .ZN(_09079_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15432_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .ZN(_09080_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3158 (.I(_11244_[0]),
    .Z(net3158));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15434_ (.A1(_08910_),
    .A2(_09079_),
    .B1(_09080_),
    .B2(_08912_),
    .ZN(_09082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15435_ (.A1(_08906_),
    .A2(_09082_),
    .ZN(_09083_));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22947__6 (.ZN(net255));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3539 (.I(net3538),
    .Z(net3539));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15438_ (.A1(\cs_registers_i.dscratch0_q[12] ),
    .A2(_08928_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[12] ),
    .C1(\cs_registers_i.mscratch_q[12] ),
    .C2(_08899_),
    .ZN(_09086_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_104_clk_i_regs (.I(clknet_6_54__leaf_clk_i_regs),
    .Z(clknet_leaf_104_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15440_ (.A1(\cs_registers_i.csr_mtvec_o[12] ),
    .A2(_08926_),
    .ZN(_09088_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _15441_ (.A1(_11438_[0]),
    .A2(_08328_),
    .B(_08329_),
    .C(_08331_),
    .ZN(_09089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15442_ (.A1(\cs_registers_i.mstatus_q[3] ),
    .A2(_09041_),
    .ZN(_09090_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15443_ (.A1(\cs_registers_i.dscratch1_q[12] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[12] ),
    .C1(net65),
    .C2(_08935_),
    .ZN(_09091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15444_ (.A1(\cs_registers_i.dcsr_q[12] ),
    .A2(_08893_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[12] ),
    .ZN(_09092_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15445_ (.A1(_09089_),
    .A2(_09090_),
    .A3(_09091_),
    .A4(_09092_),
    .Z(_09093_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15446_ (.A1(_09083_),
    .A2(_09086_),
    .A3(_09088_),
    .A4(_09093_),
    .ZN(_09094_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15447_ (.A1(_11494_[0]),
    .A2(_09094_),
    .Z(_09095_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15448_ (.A1(_09075_),
    .A2(_09095_),
    .ZN(_09096_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15449_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .A3(_09035_),
    .Z(_09097_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15450_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(_09034_),
    .A3(_09097_),
    .Z(_09098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15451_ (.A1(_09034_),
    .A2(_09097_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .C(_09003_),
    .ZN(_09099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15452_ (.A1(_09003_),
    .A2(_09096_),
    .B(_09098_),
    .C(_09099_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15453_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(_09097_),
    .Z(_09100_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15454_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .A2(_09100_),
    .Z(_09101_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_108_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_108_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_106_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_106_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15457_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11502_[0]),
    .Z(_09104_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15458_ (.A1(_11148_[0]),
    .A2(_09104_),
    .ZN(_09105_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_109_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_109_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15460_ (.A1(\cs_registers_i.mhpmcounter[1869] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .ZN(_09107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15461_ (.A1(\cs_registers_i.mhpmcounter[1901] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .ZN(_09108_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15462_ (.A1(_08912_),
    .A2(_09107_),
    .B1(_09108_),
    .B2(_08910_),
    .ZN(_09109_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15463_ (.A1(\cs_registers_i.mscratch_q[13] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[13] ),
    .ZN(_09110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15464_ (.A1(\cs_registers_i.dscratch0_q[13] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15465_ (.A1(\cs_registers_i.dscratch1_q[13] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[13] ),
    .C1(net66),
    .C2(_08935_),
    .ZN(_09112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15466_ (.A1(\cs_registers_i.dcsr_q[13] ),
    .A2(_08893_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[13] ),
    .ZN(_09113_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15467_ (.A1(_09110_),
    .A2(_09111_),
    .A3(_09112_),
    .A4(_09113_),
    .ZN(_09114_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _15468_ (.A1(\cs_registers_i.csr_mtvec_o[13] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09109_),
    .C(_09114_),
    .ZN(_09115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15469_ (.A1(_11498_[0]),
    .A2(_09115_),
    .Z(_09116_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15470_ (.A1(_09105_),
    .A2(_09116_),
    .Z(_09117_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15471_ (.A1(_09003_),
    .A2(_09117_),
    .Z(_09118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15472_ (.A1(_09071_),
    .A2(_09100_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .C(_09003_),
    .ZN(_09119_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15473_ (.A1(_09071_),
    .A2(_09101_),
    .B(_09118_),
    .C(_09119_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_110_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_110_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15475_ (.A1(\cs_registers_i.mhpmcounter[1870] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .ZN(_09121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15476_ (.A1(\cs_registers_i.mhpmcounter[1902] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .ZN(_09122_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_111_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_111_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15478_ (.A1(_08912_),
    .A2(_09121_),
    .B1(_09122_),
    .B2(_08910_),
    .ZN(_09124_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15479_ (.A1(\cs_registers_i.csr_mtvec_o[14] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09124_),
    .ZN(_09125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15480_ (.A1(\cs_registers_i.dscratch0_q[14] ),
    .A2(_08928_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[14] ),
    .C1(\cs_registers_i.mscratch_q[14] ),
    .C2(_08899_),
    .ZN(_09126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15481_ (.A1(\cs_registers_i.dscratch1_q[14] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[14] ),
    .C1(net67),
    .C2(_08935_),
    .ZN(_09127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15482_ (.A1(\cs_registers_i.mtval_q[14] ),
    .A2(_08938_),
    .B(_08924_),
    .ZN(_09128_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15483_ (.A1(_09125_),
    .A2(_09126_),
    .A3(_09127_),
    .A4(_09128_),
    .Z(_09129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15484_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11510_[0]),
    .Z(_09130_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15485_ (.A1(_11148_[0]),
    .A2(_09130_),
    .ZN(_09131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _15486_ (.A1(_11506_[0]),
    .A2(_09129_),
    .B(_09131_),
    .ZN(_09132_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _15487_ (.I(_09132_),
    .ZN(_09133_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15488_ (.A1(_09034_),
    .A2(_09101_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .C(_09003_),
    .ZN(_09134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15489_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .A2(_09034_),
    .A3(_09101_),
    .Z(_09135_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15490_ (.A1(_09003_),
    .A2(_09133_),
    .B(_09134_),
    .C(_09135_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_112_clk_i_regs (.I(clknet_6_56__leaf_clk_i_regs),
    .Z(clknet_leaf_112_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_113_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_113_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15493_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11518_[0]),
    .Z(_09138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15494_ (.A1(\cs_registers_i.mhpmcounter[1871] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .ZN(_09139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15495_ (.A1(\cs_registers_i.mhpmcounter[1903] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .ZN(_09140_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15496_ (.A1(_08912_),
    .A2(_09139_),
    .B1(_09140_),
    .B2(_08910_),
    .ZN(_09141_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15497_ (.A1(\cs_registers_i.mscratch_q[15] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[15] ),
    .ZN(_09142_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15498_ (.A1(\cs_registers_i.dscratch0_q[15] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09143_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15499_ (.A1(\cs_registers_i.dscratch1_q[15] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[15] ),
    .C1(net68),
    .C2(_08935_),
    .ZN(_09144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15500_ (.A1(\cs_registers_i.dcsr_q[15] ),
    .A2(_08893_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[15] ),
    .ZN(_09145_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15501_ (.A1(_09142_),
    .A2(_09143_),
    .A3(_09144_),
    .A4(_09145_),
    .ZN(_09146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _15502_ (.A1(\cs_registers_i.csr_mtvec_o[15] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09141_),
    .C(_09146_),
    .ZN(_09147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15503_ (.A1(_11514_[0]),
    .A2(_09147_),
    .ZN(_09148_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _15504_ (.A1(_11148_[0]),
    .A2(_09138_),
    .B(_09148_),
    .ZN(_09149_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_119_clk_i_regs (.I(clknet_6_59__leaf_clk_i_regs),
    .Z(clknet_leaf_119_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15506_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .A4(_09032_),
    .Z(_09151_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15507_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .A2(_09151_),
    .A3(_09101_),
    .Z(_09152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15508_ (.A1(_08995_),
    .A2(_09152_),
    .ZN(_09153_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_122_clk_i_regs (.I(clknet_6_59__leaf_clk_i_regs),
    .Z(clknet_leaf_122_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15510_ (.A1(_08997_),
    .A2(_09153_),
    .B(_09000_),
    .ZN(_09155_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15511_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(_09155_),
    .ZN(_09156_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15512_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(_09152_),
    .Z(_09157_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15513_ (.A1(_09030_),
    .A2(_09157_),
    .Z(_09158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15514_ (.A1(_09003_),
    .A2(_09149_),
    .B(_09156_),
    .C(_09158_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_124_clk_i_regs (.I(clknet_6_59__leaf_clk_i_regs),
    .Z(clknet_leaf_124_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15516_ (.I0(_06849_),
    .I1(_11151_[0]),
    .S(_11522_[0]),
    .Z(_09160_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15517_ (.A1(\cs_registers_i.mscratch_q[16] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[16] ),
    .ZN(_09161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15518_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(_09043_),
    .ZN(_09162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15519_ (.A1(\cs_registers_i.dscratch1_q[16] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .C1(net69),
    .C2(_08935_),
    .ZN(_09163_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_125_clk_i_regs (.I(clknet_6_59__leaf_clk_i_regs),
    .Z(clknet_leaf_125_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3159 (.I(net3158),
    .Z(net3159));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15522_ (.A1(\cs_registers_i.mhpmcounter[1872] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .ZN(_09166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15523_ (.A1(\cs_registers_i.mhpmcounter[1904] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .ZN(_09167_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15524_ (.A1(_08912_),
    .A2(_09166_),
    .B1(_09167_),
    .B2(_08910_),
    .ZN(_09168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15525_ (.A1(\cs_registers_i.dscratch0_q[16] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15526_ (.A1(\cs_registers_i.mtval_q[16] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net130),
    .ZN(_09170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15527_ (.A1(_09169_),
    .A2(_09170_),
    .ZN(_09171_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15528_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09168_),
    .C(_09171_),
    .ZN(_09172_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15529_ (.A1(_09161_),
    .A2(_09162_),
    .A3(_09163_),
    .A4(_09172_),
    .ZN(_09173_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15530_ (.A1(_11148_[0]),
    .A2(_09160_),
    .B1(_09173_),
    .B2(_11526_[0]),
    .ZN(_09174_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_126_clk_i_regs (.I(clknet_6_59__leaf_clk_i_regs),
    .Z(clknet_leaf_126_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15532_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A3(_09033_),
    .A4(_09101_),
    .Z(_09176_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15533_ (.A1(_08995_),
    .A2(_09176_),
    .Z(_09177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15534_ (.A1(_08963_),
    .A2(_08990_),
    .ZN(_09178_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15535_ (.A1(_08990_),
    .A2(_09177_),
    .B(_09178_),
    .ZN(_09179_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15536_ (.A1(_08997_),
    .A2(_09177_),
    .Z(_09180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15537_ (.I0(_09179_),
    .I1(_09180_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .Z(_09181_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15538_ (.A1(_09003_),
    .A2(_09174_),
    .B(_09181_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15539_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11534_[0]),
    .Z(_09182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15540_ (.A1(\cs_registers_i.csr_mepc_o[17] ),
    .A2(_08932_),
    .B(_08924_),
    .ZN(_09183_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15541_ (.A1(\cs_registers_i.dscratch1_q[17] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[17] ),
    .C1(net70),
    .C2(_08935_),
    .ZN(_09184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15542_ (.A1(\cs_registers_i.mstatus_q[1] ),
    .A2(_09041_),
    .B1(_09043_),
    .B2(\cs_registers_i.mie_q[1] ),
    .ZN(_09185_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15543_ (.A1(\cs_registers_i.mhpmcounter[1873] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .ZN(_09186_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15544_ (.A1(\cs_registers_i.mhpmcounter[1905] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .ZN(_09187_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15545_ (.A1(_08912_),
    .A2(_09186_),
    .B1(_09187_),
    .B2(_08910_),
    .ZN(_09188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15546_ (.A1(\cs_registers_i.dscratch0_q[17] ),
    .A2(_08928_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[17] ),
    .ZN(_09189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15547_ (.A1(\cs_registers_i.mscratch_q[17] ),
    .A2(_08899_),
    .B1(_09060_),
    .B2(net3673),
    .ZN(_09190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15548_ (.A1(_09189_),
    .A2(_09190_),
    .ZN(_09191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15549_ (.A1(\cs_registers_i.csr_mtvec_o[17] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09188_),
    .C(_09191_),
    .ZN(_09192_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15550_ (.A1(_09183_),
    .A2(_09184_),
    .A3(_09185_),
    .A4(_09192_),
    .ZN(_09193_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15551_ (.A1(_11148_[0]),
    .A2(_09182_),
    .B1(_09193_),
    .B2(_11534_[0]),
    .ZN(_09194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15552_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A2(_08992_),
    .ZN(_09195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15553_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A2(_09158_),
    .ZN(_09196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15554_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .I1(_09195_),
    .S(_09196_),
    .Z(_09197_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15555_ (.A1(_08992_),
    .A2(_09194_),
    .B(_09197_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15556_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11542_[0]),
    .Z(_09198_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15557_ (.A1(\cs_registers_i.mscratch_q[18] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[18] ),
    .ZN(_09199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15558_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(_09043_),
    .ZN(_09200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15559_ (.A1(\cs_registers_i.dscratch1_q[18] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[18] ),
    .C1(net71),
    .C2(_08935_),
    .ZN(_09201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15560_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .ZN(_09202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15561_ (.A1(\cs_registers_i.mhpmcounter[1906] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .ZN(_09203_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15562_ (.A1(net3200),
    .A2(_09202_),
    .B1(_09203_),
    .B2(net3201),
    .ZN(_09204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15563_ (.A1(\cs_registers_i.dscratch0_q[18] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15564_ (.A1(\cs_registers_i.mtval_q[18] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3672),
    .ZN(_09206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15565_ (.A1(_09205_),
    .A2(_09206_),
    .ZN(_09207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15566_ (.A1(\cs_registers_i.csr_mtvec_o[18] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09204_),
    .C(_09207_),
    .ZN(_09208_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15567_ (.A1(_09199_),
    .A2(_09200_),
    .A3(_09201_),
    .A4(_09208_),
    .ZN(_09209_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15568_ (.A1(_11148_[0]),
    .A2(_09198_),
    .B1(_09209_),
    .B2(_11542_[0]),
    .ZN(_09210_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15569_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A3(_09177_),
    .Z(_09211_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15570_ (.A1(_08990_),
    .A2(_09211_),
    .B(_09178_),
    .ZN(_09212_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15571_ (.A1(_08997_),
    .A2(_09211_),
    .Z(_09213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15572_ (.I0(_09212_),
    .I1(_09213_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .Z(_09214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15573_ (.A1(_09003_),
    .A2(_09210_),
    .B(_09214_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15574_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11550_[0]),
    .Z(_09215_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15575_ (.A1(_11148_[0]),
    .A2(_09215_),
    .ZN(_09216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15576_ (.A1(\cs_registers_i.mscratch_q[19] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[19] ),
    .ZN(_09217_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15577_ (.A1(\cs_registers_i.mie_q[3] ),
    .A2(_09043_),
    .ZN(_09218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15578_ (.A1(\cs_registers_i.dscratch1_q[19] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[19] ),
    .C1(net72),
    .C2(_08935_),
    .ZN(_09219_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15579_ (.A1(\cs_registers_i.mhpmcounter[1875] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .ZN(_09220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15580_ (.A1(\cs_registers_i.mhpmcounter[1907] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .ZN(_09221_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15581_ (.A1(net3200),
    .A2(_09220_),
    .B1(_09221_),
    .B2(net3201),
    .ZN(_09222_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15582_ (.A1(\cs_registers_i.dscratch0_q[19] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09223_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15583_ (.A1(\cs_registers_i.mtval_q[19] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3671),
    .ZN(_09224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15584_ (.A1(_09223_),
    .A2(_09224_),
    .ZN(_09225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15585_ (.A1(\cs_registers_i.csr_mtvec_o[19] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09222_),
    .C(_09225_),
    .ZN(_09226_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15586_ (.A1(_09217_),
    .A2(_09218_),
    .A3(_09219_),
    .A4(_09226_),
    .Z(_09227_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15587_ (.A1(_11546_[0]),
    .A2(_09227_),
    .Z(_09228_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15588_ (.A1(_09216_),
    .A2(_09228_),
    .Z(_09229_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15589_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .A2(_09003_),
    .ZN(_09230_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15590_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .A4(_09158_),
    .Z(_09231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15591_ (.I0(_09230_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .S(_09231_),
    .Z(_09232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15592_ (.A1(_09003_),
    .A2(_09229_),
    .B(_09232_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15593_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11402_[0]),
    .Z(_09233_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15594_ (.A1(_11148_[0]),
    .A2(_09233_),
    .Z(_09234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15595_ (.A1(\cs_registers_i.mhpmcounter[1889] ),
    .A2(_08897_),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .ZN(_09235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15596_ (.A1(\cs_registers_i.mhpmcounter[1857] ),
    .A2(_08897_),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .ZN(_09236_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15597_ (.A1(_08910_),
    .A2(_09235_),
    .B1(_09236_),
    .B2(_08912_),
    .ZN(_09237_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15598_ (.A1(\cs_registers_i.dcsr_q[1] ),
    .A2(_08893_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .ZN(_09238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15599_ (.A1(\cs_registers_i.mcause_q[1] ),
    .A2(_08898_),
    .B1(_08899_),
    .B2(\cs_registers_i.mscratch_q[1] ),
    .ZN(_09239_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15600_ (.A1(\cs_registers_i.dscratch1_q[1] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[1] ),
    .C1(net73),
    .C2(_08935_),
    .ZN(_09240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15601_ (.A1(\cs_registers_i.dscratch0_q[1] ),
    .A2(net3199),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[1] ),
    .ZN(_09241_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15602_ (.A1(_09238_),
    .A2(_09239_),
    .A3(_09240_),
    .A4(_09241_),
    .ZN(_09242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _15603_ (.A1(_08906_),
    .A2(_09237_),
    .B(_09242_),
    .ZN(_09243_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15604_ (.A1(_11406_[0]),
    .A2(_09243_),
    .ZN(_09244_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15605_ (.A1(_09234_),
    .A2(_09244_),
    .Z(_09245_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3156 (.I(_11252_[0]),
    .Z(net3156));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15607_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .I1(_11166_[0]),
    .S(_09030_),
    .Z(_09247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15608_ (.I0(_09245_),
    .I1(_09247_),
    .S(_08992_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15609_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .Z(_09248_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15610_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .A2(_09248_),
    .Z(_09249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15611_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11558_[0]),
    .Z(_09250_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15612_ (.A1(\cs_registers_i.mhpmcounter[1908] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .ZN(_09251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15613_ (.A1(\cs_registers_i.mhpmcounter[1876] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .ZN(_09252_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15614_ (.A1(_08910_),
    .A2(_09251_),
    .B1(_09252_),
    .B2(_08912_),
    .ZN(_09253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15615_ (.A1(_08906_),
    .A2(_09253_),
    .ZN(_09254_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15616_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_08926_),
    .ZN(_09255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15617_ (.A1(\cs_registers_i.dscratch1_q[20] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[20] ),
    .C1(net74),
    .C2(_08935_),
    .ZN(_09256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15618_ (.A1(\cs_registers_i.mscratch_q[20] ),
    .A2(_08899_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[20] ),
    .ZN(_09257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15619_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(_09043_),
    .ZN(_09258_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15620_ (.A1(_09089_),
    .A2(_09256_),
    .A3(_09257_),
    .A4(_09258_),
    .Z(_09259_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15621_ (.A1(\cs_registers_i.dscratch0_q[20] ),
    .A2(_08928_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[20] ),
    .C1(_09060_),
    .C2(net3670),
    .ZN(_09260_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15622_ (.A1(_09254_),
    .A2(_09255_),
    .A3(_09259_),
    .A4(_09260_),
    .ZN(_09261_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15623_ (.A1(_11148_[0]),
    .A2(_09250_),
    .B1(_09261_),
    .B2(_11558_[0]),
    .ZN(_09262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15624_ (.A1(_09180_),
    .A2(_09248_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .ZN(_09263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15625_ (.I0(_09262_),
    .I1(_09263_),
    .S(_08992_),
    .Z(_09264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15626_ (.A1(_09180_),
    .A2(_09249_),
    .B(_09264_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15627_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11566_[0]),
    .Z(_09265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15628_ (.A1(\cs_registers_i.dscratch0_q[21] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15629_ (.A1(\cs_registers_i.dscratch1_q[21] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[21] ),
    .C1(net75),
    .C2(_08935_),
    .ZN(_09267_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15630_ (.A1(\cs_registers_i.csr_mstatus_tw_o ),
    .A2(_09041_),
    .B1(_09043_),
    .B2(\cs_registers_i.mie_q[5] ),
    .ZN(_09268_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15631_ (.A1(\cs_registers_i.mhpmcounter[1909] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .ZN(_09269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15632_ (.A1(\cs_registers_i.mhpmcounter[1877] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .ZN(_09270_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15633_ (.A1(_08910_),
    .A2(_09269_),
    .B1(_09270_),
    .B2(_08912_),
    .ZN(_09271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15634_ (.A1(\cs_registers_i.mscratch_q[21] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[21] ),
    .ZN(_09272_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15635_ (.A1(\cs_registers_i.mtval_q[21] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3669),
    .ZN(_09273_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15636_ (.A1(_09272_),
    .A2(_09273_),
    .ZN(_09274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15637_ (.A1(\cs_registers_i.csr_mtvec_o[21] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09271_),
    .C(_09274_),
    .ZN(_09275_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15638_ (.A1(_09266_),
    .A2(_09267_),
    .A3(_09268_),
    .A4(_09275_),
    .ZN(_09276_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15639_ (.A1(_11148_[0]),
    .A2(_09265_),
    .B1(_09276_),
    .B2(_11566_[0]),
    .ZN(_09277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15640_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A2(_08992_),
    .ZN(_09278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15641_ (.A1(_09158_),
    .A2(_09249_),
    .ZN(_09279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15642_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .I1(_09278_),
    .S(_09279_),
    .Z(_09280_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15643_ (.A1(_08992_),
    .A2(_09277_),
    .B(_09280_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15644_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11574_[0]),
    .Z(_09281_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15645_ (.A1(\cs_registers_i.mscratch_q[22] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[22] ),
    .ZN(_09282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15646_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(_09043_),
    .ZN(_09283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15647_ (.A1(\cs_registers_i.dscratch1_q[22] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[22] ),
    .C1(net76),
    .C2(_08935_),
    .ZN(_09284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15648_ (.A1(\cs_registers_i.mhpmcounter[1878] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .ZN(_09285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15649_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .ZN(_09286_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15650_ (.A1(net3200),
    .A2(_09285_),
    .B1(_09286_),
    .B2(net3201),
    .ZN(_09287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15651_ (.A1(\cs_registers_i.dscratch0_q[22] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15652_ (.A1(\cs_registers_i.mtval_q[22] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3668),
    .ZN(_09289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15653_ (.A1(_09288_),
    .A2(_09289_),
    .ZN(_09290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15654_ (.A1(\cs_registers_i.csr_mtvec_o[22] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09287_),
    .C(_09290_),
    .ZN(_09291_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15655_ (.A1(_09282_),
    .A2(_09283_),
    .A3(_09284_),
    .A4(_09291_),
    .ZN(_09292_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15656_ (.A1(_11148_[0]),
    .A2(_09281_),
    .B1(_09292_),
    .B2(_11574_[0]),
    .ZN(_09293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15657_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .A2(_08992_),
    .ZN(_09294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15658_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A2(_09249_),
    .Z(_09295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15659_ (.A1(_09180_),
    .A2(_09295_),
    .ZN(_09296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15660_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .I1(_09294_),
    .S(_09296_),
    .Z(_09297_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15661_ (.A1(_08992_),
    .A2(_09293_),
    .B(_09297_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15662_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11582_[0]),
    .Z(_09298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15663_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(_09043_),
    .ZN(_09299_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15664_ (.A1(\cs_registers_i.dscratch1_q[23] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[23] ),
    .C1(net77),
    .C2(_08935_),
    .ZN(_09300_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15665_ (.A1(\cs_registers_i.csr_mepc_o[23] ),
    .A2(_08932_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[23] ),
    .ZN(_09301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15666_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .ZN(_09302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15667_ (.A1(\cs_registers_i.mhpmcounter[1911] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .ZN(_09303_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15668_ (.A1(net3200),
    .A2(_09302_),
    .B1(_09303_),
    .B2(net3201),
    .ZN(_09304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15669_ (.A1(\cs_registers_i.dscratch0_q[23] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09305_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15670_ (.A1(\cs_registers_i.mscratch_q[23] ),
    .A2(_08899_),
    .B1(_09060_),
    .B2(net3667),
    .ZN(_09306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15671_ (.A1(_09305_),
    .A2(_09306_),
    .ZN(_09307_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15672_ (.A1(\cs_registers_i.csr_mtvec_o[23] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09304_),
    .C(_09307_),
    .ZN(_09308_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15673_ (.A1(_09299_),
    .A2(_09300_),
    .A3(_09301_),
    .A4(_09308_),
    .ZN(_09309_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15674_ (.A1(_11148_[0]),
    .A2(_09298_),
    .B1(_09309_),
    .B2(_11582_[0]),
    .ZN(_09310_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3204 (.I(net3203),
    .Z(net3204));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15676_ (.A1(_08995_),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .A3(_09157_),
    .A4(_09295_),
    .Z(_09312_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15677_ (.A1(_08990_),
    .A2(_09312_),
    .Z(_09313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15678_ (.A1(_09178_),
    .A2(_09313_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .ZN(_09314_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15679_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .A2(_08997_),
    .A3(_09312_),
    .Z(_09315_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15680_ (.A1(_09003_),
    .A2(_09310_),
    .B(_09314_),
    .C(_09315_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15681_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11590_[0]),
    .Z(_09316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15682_ (.A1(\cs_registers_i.mhpmcounter[1880] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .ZN(_09317_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15683_ (.A1(\cs_registers_i.mhpmcounter[1912] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .ZN(_09318_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15684_ (.A1(_08912_),
    .A2(_09317_),
    .B1(_09318_),
    .B2(net3201),
    .ZN(_09319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15685_ (.A1(_08906_),
    .A2(_09319_),
    .Z(_09320_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15686_ (.A1(\cs_registers_i.csr_mtvec_o[24] ),
    .A2(_08926_),
    .Z(_09321_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15687_ (.A1(\cs_registers_i.mscratch_q[24] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[24] ),
    .ZN(_09322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15688_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(_09043_),
    .ZN(_09323_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15689_ (.A1(\cs_registers_i.dscratch1_q[24] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[24] ),
    .C1(net78),
    .C2(_08935_),
    .ZN(_09324_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15690_ (.A1(_09322_),
    .A2(_09323_),
    .A3(_09324_),
    .ZN(_09325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15691_ (.A1(\cs_registers_i.dscratch0_q[24] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15692_ (.A1(\cs_registers_i.mtval_q[24] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3666),
    .ZN(_09327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15693_ (.A1(_09326_),
    .A2(_09327_),
    .ZN(_09328_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _15694_ (.A1(_09320_),
    .A2(_09321_),
    .A3(_09325_),
    .A4(_09328_),
    .Z(_09329_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15695_ (.A1(_11148_[0]),
    .A2(_09316_),
    .B1(_09329_),
    .B2(_11590_[0]),
    .ZN(_09330_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15696_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .A3(_09295_),
    .Z(_09331_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15697_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .A2(_09180_),
    .A3(_09331_),
    .Z(_09332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15698_ (.A1(_09180_),
    .A2(_09331_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .C(_09003_),
    .ZN(_09333_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15699_ (.A1(_09003_),
    .A2(_09330_),
    .B(_09332_),
    .C(_09333_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15700_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11598_[0]),
    .Z(_09334_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15701_ (.A1(_11148_[0]),
    .A2(_09334_),
    .ZN(_09335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15702_ (.A1(\cs_registers_i.mscratch_q[25] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[25] ),
    .ZN(_09336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15703_ (.A1(\cs_registers_i.mie_q[9] ),
    .A2(_09043_),
    .ZN(_09337_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15704_ (.A1(\cs_registers_i.dscratch1_q[25] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[25] ),
    .C1(net79),
    .C2(_08935_),
    .ZN(_09338_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15705_ (.A1(\cs_registers_i.mhpmcounter[1881] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .ZN(_09339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15706_ (.A1(\cs_registers_i.mhpmcounter[1913] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .ZN(_09340_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15707_ (.A1(net3200),
    .A2(_09339_),
    .B1(_09340_),
    .B2(net3201),
    .ZN(_09341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15708_ (.A1(\cs_registers_i.dscratch0_q[25] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09342_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15709_ (.A1(\cs_registers_i.mtval_q[25] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3665),
    .ZN(_09343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15710_ (.A1(_09342_),
    .A2(_09343_),
    .ZN(_09344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15711_ (.A1(\cs_registers_i.csr_mtvec_o[25] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09341_),
    .C(_09344_),
    .ZN(_09345_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15712_ (.A1(_09336_),
    .A2(_09337_),
    .A3(_09338_),
    .A4(_09345_),
    .Z(_09346_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15713_ (.A1(_11594_[0]),
    .A2(_09346_),
    .Z(_09347_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15714_ (.A1(_09335_),
    .A2(_09347_),
    .Z(_09348_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15715_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .A3(_09331_),
    .Z(_09349_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15716_ (.A1(_09030_),
    .A2(_09157_),
    .A3(_09349_),
    .Z(_09350_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15717_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .A2(_09158_),
    .A3(_09331_),
    .Z(_09351_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _15718_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .A2(_09003_),
    .A3(_09351_),
    .ZN(_09352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15719_ (.A1(_09003_),
    .A2(_09348_),
    .B(_09350_),
    .C(_09352_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15720_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11606_[0]),
    .Z(_09353_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15721_ (.A1(\cs_registers_i.mhpmcounter[1882] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .ZN(_09354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15722_ (.A1(\cs_registers_i.mhpmcounter[1914] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .ZN(_09355_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15723_ (.A1(net3200),
    .A2(_09354_),
    .B1(_09355_),
    .B2(net3201),
    .ZN(_09356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15724_ (.A1(_08906_),
    .A2(_09356_),
    .Z(_09357_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15725_ (.A1(\cs_registers_i.csr_mtvec_o[26] ),
    .A2(_08926_),
    .Z(_09358_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15726_ (.A1(\cs_registers_i.mscratch_q[26] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[26] ),
    .ZN(_09359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15727_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(_09043_),
    .ZN(_09360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15728_ (.A1(\cs_registers_i.dscratch1_q[26] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[26] ),
    .C1(net80),
    .C2(_08935_),
    .ZN(_09361_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15729_ (.A1(_09359_),
    .A2(_09360_),
    .A3(_09361_),
    .ZN(_09362_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15730_ (.A1(\cs_registers_i.dscratch0_q[26] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09363_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15731_ (.A1(\cs_registers_i.mtval_q[26] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3677),
    .ZN(_09364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15732_ (.A1(_09363_),
    .A2(_09364_),
    .ZN(_09365_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _15733_ (.A1(_09357_),
    .A2(_09358_),
    .A3(_09362_),
    .A4(_09365_),
    .Z(_09366_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15734_ (.A1(_11148_[0]),
    .A2(_09353_),
    .B1(_09366_),
    .B2(_11606_[0]),
    .ZN(_09367_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15735_ (.A1(_09177_),
    .A2(_09349_),
    .Z(_09368_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15736_ (.A1(_08990_),
    .A2(_09368_),
    .B(_09178_),
    .ZN(_09369_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15737_ (.A1(_08997_),
    .A2(_09368_),
    .Z(_09370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15738_ (.I0(_09369_),
    .I1(_09370_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .Z(_09371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15739_ (.A1(_09003_),
    .A2(_09367_),
    .B(_09371_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15740_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11614_[0]),
    .Z(_09372_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15741_ (.A1(\cs_registers_i.mscratch_q[27] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[27] ),
    .ZN(_09373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15742_ (.A1(\cs_registers_i.mie_q[11] ),
    .A2(_09043_),
    .ZN(_09374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15743_ (.A1(\cs_registers_i.dscratch1_q[27] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[27] ),
    .C1(net81),
    .C2(_08935_),
    .ZN(_09375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15744_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .ZN(_09376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15745_ (.A1(\cs_registers_i.mhpmcounter[1915] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .ZN(_09377_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15746_ (.A1(net3200),
    .A2(_09376_),
    .B1(_09377_),
    .B2(net3201),
    .ZN(_09378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15747_ (.A1(\cs_registers_i.dscratch0_q[27] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15748_ (.A1(\cs_registers_i.mtval_q[27] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3676),
    .ZN(_09380_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15749_ (.A1(_09379_),
    .A2(_09380_),
    .ZN(_09381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15750_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09378_),
    .C(_09381_),
    .ZN(_09382_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15751_ (.A1(_09373_),
    .A2(_09374_),
    .A3(_09375_),
    .A4(_09382_),
    .ZN(_09383_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15752_ (.A1(_11148_[0]),
    .A2(_09372_),
    .B1(_09383_),
    .B2(_11614_[0]),
    .ZN(_09384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15753_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(_09350_),
    .B(_09003_),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .ZN(_09385_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15754_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A3(_09350_),
    .Z(_09386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15755_ (.A1(_09003_),
    .A2(_09384_),
    .B(_09385_),
    .C(_09386_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15756_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11622_[0]),
    .Z(_09387_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _15757_ (.A1(_11148_[0]),
    .A2(_09387_),
    .ZN(_09388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15758_ (.A1(\cs_registers_i.mscratch_q[28] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[28] ),
    .ZN(_09389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15759_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(_09043_),
    .ZN(_09390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15760_ (.A1(\cs_registers_i.dscratch1_q[28] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[28] ),
    .C1(net82),
    .C2(_08935_),
    .ZN(_09391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15761_ (.A1(\cs_registers_i.mhpmcounter[1884] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .ZN(_09392_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15762_ (.A1(\cs_registers_i.mhpmcounter[1916] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .ZN(_09393_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15763_ (.A1(net3200),
    .A2(_09392_),
    .B1(_09393_),
    .B2(net3201),
    .ZN(_09394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15764_ (.A1(\cs_registers_i.dscratch0_q[28] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09395_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15765_ (.A1(\cs_registers_i.mtval_q[28] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3675),
    .ZN(_09396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15766_ (.A1(_09395_),
    .A2(_09396_),
    .ZN(_09397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15767_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09394_),
    .C(_09397_),
    .ZN(_09398_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15768_ (.A1(_09389_),
    .A2(_09390_),
    .A3(_09391_),
    .A4(_09398_),
    .Z(_09399_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15769_ (.A1(_11618_[0]),
    .A2(_09399_),
    .Z(_09400_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15770_ (.A1(_09388_),
    .A2(_09400_),
    .Z(_09401_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15771_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A2(_09003_),
    .ZN(_09402_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15772_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A3(_09370_),
    .Z(_09403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15773_ (.I0(_09402_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .S(_09403_),
    .Z(_09404_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15774_ (.A1(_09003_),
    .A2(_09401_),
    .B(_09404_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15775_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11630_[0]),
    .Z(_09405_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _15776_ (.A1(_11148_[0]),
    .A2(_09405_),
    .ZN(_09406_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15777_ (.A1(\cs_registers_i.mscratch_q[29] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[29] ),
    .ZN(_09407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15778_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(_09043_),
    .ZN(_09408_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15779_ (.A1(\cs_registers_i.dscratch1_q[29] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[29] ),
    .C1(net83),
    .C2(_08935_),
    .ZN(_09409_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15780_ (.A1(\cs_registers_i.mhpmcounter[1885] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .ZN(_09410_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15781_ (.A1(\cs_registers_i.mhpmcounter[1917] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .ZN(_09411_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15782_ (.A1(net3200),
    .A2(_09410_),
    .B1(_09411_),
    .B2(net3201),
    .ZN(_09412_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15783_ (.A1(\cs_registers_i.dscratch0_q[29] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09413_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15784_ (.A1(\cs_registers_i.mtval_q[29] ),
    .A2(_08938_),
    .B1(_09060_),
    .B2(net3674),
    .ZN(_09414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15785_ (.A1(_09413_),
    .A2(_09414_),
    .ZN(_09415_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15786_ (.A1(\cs_registers_i.csr_mtvec_o[29] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09412_),
    .C(_09415_),
    .ZN(_09416_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15787_ (.A1(_09407_),
    .A2(_09408_),
    .A3(_09409_),
    .A4(_09416_),
    .Z(_09417_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15788_ (.A1(_11626_[0]),
    .A2(_09417_),
    .Z(_09418_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15789_ (.A1(_09406_),
    .A2(_09418_),
    .Z(_09419_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15790_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .A2(_09003_),
    .ZN(_09420_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15791_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A4(_09350_),
    .Z(_09421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15792_ (.I0(_09420_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .S(_09421_),
    .Z(_09422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15793_ (.A1(_09003_),
    .A2(_09419_),
    .B(_09422_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _15794_ (.A1(_11409_[0]),
    .A2(_08982_),
    .B(_08956_),
    .ZN(_09423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15795_ (.A1(_08995_),
    .A2(_11165_[0]),
    .ZN(_09424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15796_ (.A1(_08997_),
    .A2(_09424_),
    .ZN(_09425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15797_ (.A1(_09178_),
    .A2(_09425_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .ZN(_09426_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15798_ (.A1(_09423_),
    .A2(_09003_),
    .B1(_09031_),
    .B2(_09030_),
    .C(_09426_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15799_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11638_[0]),
    .Z(_09427_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15800_ (.A1(_11148_[0]),
    .A2(_09427_),
    .Z(_09428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15801_ (.A1(\cs_registers_i.mscratch_q[30] ),
    .A2(_08899_),
    .B1(_08928_),
    .B2(\cs_registers_i.dscratch0_q[30] ),
    .ZN(_09429_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15802_ (.A1(net85),
    .A2(_08935_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[30] ),
    .ZN(_09430_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15803_ (.A1(\cs_registers_i.dscratch1_q[30] ),
    .A2(_08940_),
    .B(_08893_),
    .ZN(_09431_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15804_ (.A1(_09429_),
    .A2(_09430_),
    .A3(_09431_),
    .Z(_09432_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15805_ (.A1(\cs_registers_i.mie_q[14] ),
    .A2(_09043_),
    .ZN(_09433_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15806_ (.A1(\cs_registers_i.mhpmcounter[1886] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .ZN(_09434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15807_ (.A1(\cs_registers_i.mhpmcounter[1918] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .ZN(_09435_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15808_ (.A1(net3200),
    .A2(_09434_),
    .B1(_09435_),
    .B2(net3201),
    .ZN(_09436_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15809_ (.A1(\cs_registers_i.csr_mepc_o[30] ),
    .A2(_08932_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[30] ),
    .C1(net135),
    .C2(_09060_),
    .ZN(_09437_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15810_ (.I(_09437_),
    .ZN(_09438_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15811_ (.A1(\cs_registers_i.csr_mtvec_o[30] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09436_),
    .C(_09438_),
    .ZN(_09439_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15812_ (.A1(_09089_),
    .A2(_09432_),
    .A3(_09433_),
    .A4(_09439_),
    .ZN(_09440_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _15813_ (.A1(_11638_[0]),
    .A2(_09440_),
    .Z(_09441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15814_ (.A1(_09428_),
    .A2(_09441_),
    .ZN(_09442_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15815_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .Z(_09443_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15816_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .A2(_09370_),
    .A3(_09443_),
    .Z(_09444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15817_ (.A1(_09370_),
    .A2(_09443_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .C(_09003_),
    .ZN(_09445_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15818_ (.A1(_09003_),
    .A2(_09442_),
    .B(_09444_),
    .C(_09445_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15819_ (.A1(\cs_registers_i.mhpmcounter[1887] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .ZN(_09446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15820_ (.A1(\cs_registers_i.mhpmcounter[1919] ),
    .A2(net3211),
    .B1(net3209),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .ZN(_09447_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15821_ (.A1(net3200),
    .A2(_09446_),
    .B1(_09447_),
    .B2(net3201),
    .ZN(_09448_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15822_ (.A1(\cs_registers_i.mscratch_q[31] ),
    .A2(_08899_),
    .B1(_08928_),
    .B2(\cs_registers_i.dscratch0_q[31] ),
    .ZN(_09449_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15823_ (.A1(\cs_registers_i.mcause_q[5] ),
    .A2(_08898_),
    .B(_08924_),
    .ZN(_09450_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15824_ (.A1(\cs_registers_i.csr_mepc_o[31] ),
    .A2(_08932_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[31] ),
    .ZN(_09451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15825_ (.A1(\cs_registers_i.dscratch1_q[31] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[31] ),
    .C1(net86),
    .C2(_08935_),
    .ZN(_09452_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15826_ (.A1(_09449_),
    .A2(_09450_),
    .A3(_09451_),
    .A4(_09452_),
    .ZN(_09453_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _15827_ (.A1(\cs_registers_i.csr_mtvec_o[31] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09448_),
    .C(_09453_),
    .ZN(_09454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15828_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11143_[0]),
    .Z(_09455_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15829_ (.A1(_11148_[0]),
    .A2(_09455_),
    .ZN(_09456_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _15830_ (.A1(_11139_[0]),
    .A2(_09454_),
    .B(_09456_),
    .ZN(_09457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _15831_ (.I(_09457_),
    .ZN(_09458_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15832_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .A2(_09003_),
    .ZN(_09459_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15833_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .A2(_09350_),
    .A3(_09443_),
    .Z(_09460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15834_ (.I0(_09459_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .S(_09460_),
    .Z(_09461_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15835_ (.A1(_09003_),
    .A2(_09458_),
    .B(_09461_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3154 (.I(_03393_),
    .Z(net3154));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15837_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .A3(_09443_),
    .Z(_09463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15838_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .A2(_09463_),
    .Z(_09464_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15839_ (.A1(_09349_),
    .A2(_09464_),
    .Z(_09465_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15840_ (.A1(_09370_),
    .A2(_09463_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .C(_09000_),
    .ZN(_09466_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15841_ (.A1(_08985_),
    .A2(_09000_),
    .B1(_09180_),
    .B2(_09465_),
    .C(_09466_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3185 (.I(_03232_),
    .Z(net3185));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15843_ (.A1(_09234_),
    .A2(_09244_),
    .ZN(_09468_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15844_ (.A1(_09157_),
    .A2(_09349_),
    .Z(_09469_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15845_ (.A1(_08995_),
    .A2(_09464_),
    .A3(_09469_),
    .Z(_09470_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15846_ (.A1(_08990_),
    .A2(_09470_),
    .B(_08992_),
    .ZN(_09471_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15847_ (.A1(_08997_),
    .A2(_09470_),
    .Z(_09472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15848_ (.I0(_09471_),
    .I1(_09472_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .Z(_09473_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15849_ (.A1(_09000_),
    .A2(_09468_),
    .B(_09473_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15850_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(_09368_),
    .A3(_09464_),
    .Z(_09474_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15851_ (.A1(_08990_),
    .A2(_09474_),
    .Z(_09475_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15852_ (.A1(_08992_),
    .A2(_09475_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .ZN(_09476_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15853_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A2(_08997_),
    .A3(_09474_),
    .Z(_09477_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15854_ (.A1(_09423_),
    .A2(_09000_),
    .B(_09476_),
    .C(_09477_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15855_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11417_[0]),
    .Z(_09478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15856_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(_09041_),
    .ZN(_09479_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15857_ (.A1(\cs_registers_i.mie_q[17] ),
    .A2(_09043_),
    .ZN(_09480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15858_ (.A1(\cs_registers_i.dscratch1_q[3] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[3] ),
    .C1(net87),
    .C2(_08935_),
    .ZN(_09481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15859_ (.A1(\cs_registers_i.mhpmcounter[1859] ),
    .A2(_08897_),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .ZN(_09482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15860_ (.A1(\cs_registers_i.mhpmcounter[1891] ),
    .A2(_08897_),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .ZN(_09483_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15861_ (.A1(_08912_),
    .A2(_09482_),
    .B1(_09483_),
    .B2(_08910_),
    .ZN(_09484_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15862_ (.A1(_08906_),
    .A2(_09484_),
    .ZN(_09485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15863_ (.A1(\cs_registers_i.mscratch_q[3] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[3] ),
    .ZN(_09486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15864_ (.A1(\cs_registers_i.dscratch0_q[3] ),
    .A2(net3199),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[3] ),
    .C1(\cs_registers_i.mcause_q[3] ),
    .C2(_08898_),
    .ZN(_09487_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15865_ (.A1(net146),
    .A2(_09060_),
    .B(_08924_),
    .ZN(_09488_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15866_ (.A1(_09485_),
    .A2(_09486_),
    .A3(_09487_),
    .A4(_09488_),
    .Z(_09489_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _15867_ (.A1(_09479_),
    .A2(_09480_),
    .A3(_09481_),
    .A4(_09489_),
    .ZN(_09490_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15868_ (.A1(_11148_[0]),
    .A2(_09478_),
    .B1(_09490_),
    .B2(_11417_[0]),
    .ZN(_09491_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3153 (.I(_11255_[0]),
    .Z(net3153));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15870_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .A2(_09000_),
    .ZN(_09493_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15871_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A3(_09472_),
    .Z(_09494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15872_ (.I0(_09493_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .S(_09494_),
    .Z(_09495_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15873_ (.A1(_09000_),
    .A2(_09491_),
    .B(_09495_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3152 (.I(_11256_[0]),
    .Z(net3152));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15875_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(net3252),
    .Z(_09497_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15876_ (.A1(\cs_registers_i.mhpmcounter[1892] ),
    .A2(_08897_),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .ZN(_09498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15877_ (.A1(\cs_registers_i.mhpmcounter[1860] ),
    .A2(_08897_),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .ZN(_09499_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15878_ (.A1(_08910_),
    .A2(_09498_),
    .B1(_09499_),
    .B2(_08912_),
    .ZN(_09500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15879_ (.A1(\cs_registers_i.mcause_q[4] ),
    .A2(_08898_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[4] ),
    .ZN(_09501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15880_ (.A1(\cs_registers_i.dscratch0_q[4] ),
    .A2(net3199),
    .B(_08924_),
    .ZN(_09502_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15881_ (.A1(\cs_registers_i.mscratch_q[4] ),
    .A2(_08899_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[4] ),
    .ZN(_09503_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15882_ (.A1(\cs_registers_i.dscratch1_q[4] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[4] ),
    .C1(net88),
    .C2(_08935_),
    .ZN(_09504_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15883_ (.A1(_09501_),
    .A2(_09502_),
    .A3(_09503_),
    .A4(_09504_),
    .ZN(_09505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15884_ (.A1(_08906_),
    .A2(_09500_),
    .B(_09505_),
    .ZN(_09506_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _15885_ (.I(_09506_),
    .ZN(_09507_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15886_ (.A1(_11148_[0]),
    .A2(_09497_),
    .B1(_09507_),
    .B2(net3252),
    .ZN(_09508_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15887_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .Z(_09509_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15888_ (.A1(_09177_),
    .A2(_09465_),
    .A3(_09509_),
    .ZN(_09510_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15889_ (.A1(_08997_),
    .A2(_09510_),
    .Z(_09511_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15890_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(_09003_),
    .A3(_09511_),
    .Z(_09512_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15891_ (.A1(_08990_),
    .A2(_09510_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .ZN(_09513_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15892_ (.A1(_09000_),
    .A2(_09508_),
    .B1(_09512_),
    .B2(_09513_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15893_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11433_[0]),
    .Z(_09514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15894_ (.A1(\cs_registers_i.mhpmcounter[1893] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .ZN(_09515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15895_ (.A1(\cs_registers_i.mhpmcounter[1861] ),
    .A2(_08897_),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .ZN(_09516_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15896_ (.A1(_08910_),
    .A2(_09515_),
    .B1(_09516_),
    .B2(_08912_),
    .ZN(_09517_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15897_ (.A1(_08906_),
    .A2(_09517_),
    .ZN(_09518_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15898_ (.A1(\cs_registers_i.dscratch0_q[5] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15899_ (.A1(\cs_registers_i.mscratch_q[5] ),
    .A2(_08899_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[5] ),
    .C1(\cs_registers_i.mtval_q[5] ),
    .C2(_08938_),
    .ZN(_09520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15900_ (.A1(\cs_registers_i.dscratch1_q[5] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[5] ),
    .C1(net89),
    .C2(_08935_),
    .ZN(_09521_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15901_ (.A1(_09518_),
    .A2(_09519_),
    .A3(_09520_),
    .A4(_09521_),
    .Z(_09522_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15902_ (.A1(_11437_[0]),
    .A2(_09522_),
    .ZN(_09523_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _15903_ (.A1(_11148_[0]),
    .A2(_09514_),
    .B(_09523_),
    .ZN(_09524_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15904_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(_09509_),
    .Z(_09525_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15905_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(_09472_),
    .A3(_09525_),
    .Z(_09526_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15906_ (.A1(_09470_),
    .A2(_09525_),
    .Z(_09527_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15907_ (.A1(_08990_),
    .A2(_09527_),
    .Z(_09528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15908_ (.A1(_08992_),
    .A2(_09528_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .ZN(_09529_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15909_ (.A1(_09000_),
    .A2(_09524_),
    .B(_09526_),
    .C(_09529_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15910_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11441_[0]),
    .Z(_09530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15911_ (.A1(\cs_registers_i.mhpmcounter[1894] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .ZN(_09531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15912_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .ZN(_09532_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15913_ (.A1(_08910_),
    .A2(_09531_),
    .B1(_09532_),
    .B2(_08912_),
    .ZN(_09533_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15914_ (.A1(\cs_registers_i.dcsr_q[6] ),
    .A2(_08893_),
    .B1(_08899_),
    .B2(\cs_registers_i.mscratch_q[6] ),
    .ZN(_09534_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15915_ (.A1(\cs_registers_i.dscratch0_q[6] ),
    .A2(_08928_),
    .B(_08924_),
    .ZN(_09535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15916_ (.A1(\cs_registers_i.csr_mepc_o[6] ),
    .A2(_08932_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[6] ),
    .ZN(_09536_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15917_ (.A1(\cs_registers_i.dscratch1_q[6] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[6] ),
    .C1(net90),
    .C2(_08935_),
    .ZN(_09537_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15918_ (.A1(_09534_),
    .A2(_09535_),
    .A3(_09536_),
    .A4(_09537_),
    .ZN(_09538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15919_ (.A1(_08906_),
    .A2(_09533_),
    .B(_09538_),
    .ZN(_09539_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _15920_ (.I(_09539_),
    .ZN(_09540_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15921_ (.A1(_11148_[0]),
    .A2(_09530_),
    .B1(_09540_),
    .B2(_11441_[0]),
    .ZN(_09541_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15922_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(_09464_),
    .A3(_09525_),
    .Z(_09542_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15923_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(_08997_),
    .A3(_09368_),
    .A4(_09542_),
    .Z(_09543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15924_ (.A1(_09368_),
    .A2(_09542_),
    .ZN(_09544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15925_ (.A1(_08997_),
    .A2(_09544_),
    .ZN(_09545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15926_ (.A1(_08992_),
    .A2(_09545_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .ZN(_09546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15927_ (.A1(_09000_),
    .A2(_09541_),
    .B(_09543_),
    .C(_09546_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15928_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11449_[0]),
    .Z(_09547_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3211 (.I(_08897_),
    .Z(net3211));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15930_ (.A1(_06530_),
    .A2(_08310_),
    .A3(_08313_),
    .Z(_09549_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15931_ (.A1(net301),
    .A2(net263),
    .A3(_08313_),
    .A4(_08348_),
    .Z(_09550_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15932_ (.A1(_09549_),
    .A2(_08352_),
    .A3(_09550_),
    .Z(_09551_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15933_ (.A1(_11486_[0]),
    .A2(_08324_),
    .A3(_09549_),
    .Z(_09552_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _15934_ (.A1(_06388_),
    .A2(net485),
    .A3(_08327_),
    .B(_08313_),
    .ZN(_09553_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15935_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_09552_),
    .A3(_09553_),
    .Z(_09554_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15936_ (.A1(net91),
    .A2(_09551_),
    .B(_09554_),
    .ZN(_09555_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15937_ (.A1(_08314_),
    .A2(_08318_),
    .ZN(_09556_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15938_ (.A1(_09550_),
    .A2(_09556_),
    .Z(_09557_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15939_ (.A1(_06388_),
    .A2(net329),
    .A3(_08930_),
    .A4(_08313_),
    .Z(_09558_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15940_ (.A1(\cs_registers_i.csr_depc_o[7] ),
    .A2(_09552_),
    .A3(_09558_),
    .Z(_09559_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15941_ (.A1(net147),
    .A2(_09557_),
    .B(_09559_),
    .ZN(_09560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15942_ (.A1(net3287),
    .A2(_08280_),
    .ZN(_09561_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15943_ (.A1(_08314_),
    .A2(_09561_),
    .ZN(_09562_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15944_ (.A1(_11434_[0]),
    .A2(_09553_),
    .A3(_09562_),
    .Z(_09563_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15945_ (.A1(_06388_),
    .A2(net485),
    .A3(_08930_),
    .A4(_08313_),
    .Z(_09564_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15946_ (.A1(\cs_registers_i.mtval_q[7] ),
    .A2(_09556_),
    .A3(_09564_),
    .Z(_09565_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15947_ (.A1(_09563_),
    .A2(_09565_),
    .ZN(_09566_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15948_ (.A1(\cs_registers_i.mscratch_q[7] ),
    .A2(_09553_),
    .A3(_09556_),
    .Z(_09567_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15949_ (.A1(\cs_registers_i.dscratch1_q[7] ),
    .A2(_09552_),
    .A3(_09564_),
    .Z(_09568_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15950_ (.A1(_09567_),
    .A2(_09568_),
    .ZN(_09569_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15951_ (.A1(_09555_),
    .A2(_09560_),
    .A3(_09566_),
    .A4(_09569_),
    .Z(_09570_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _15952_ (.A1(_11434_[0]),
    .A2(_08314_),
    .A3(_09561_),
    .ZN(_09571_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15953_ (.A1(\cs_registers_i.mstatus_q[4] ),
    .A2(_09553_),
    .A3(_09571_),
    .Z(_09572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15954_ (.A1(_08327_),
    .A2(_08313_),
    .ZN(_09573_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15955_ (.A1(net301),
    .A2(net485),
    .A3(_08313_),
    .Z(_09574_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15956_ (.A1(\cs_registers_i.dscratch0_q[7] ),
    .A2(_09573_),
    .A3(_09552_),
    .A4(_09574_),
    .Z(_09575_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15957_ (.A1(_09572_),
    .A2(_09575_),
    .ZN(_09576_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15958_ (.A1(_09550_),
    .A2(_09571_),
    .Z(_09577_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15959_ (.A1(\cs_registers_i.csr_mepc_o[7] ),
    .A2(_09558_),
    .A3(_09556_),
    .Z(_09578_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15960_ (.A1(\cs_registers_i.mie_q[16] ),
    .A2(_09577_),
    .B(_09578_),
    .ZN(_09579_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _15961_ (.A1(_06530_),
    .A2(_08327_),
    .B(_08313_),
    .ZN(_09580_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15962_ (.A1(_06811_),
    .A2(_08313_),
    .A3(_08298_),
    .A4(_08339_),
    .Z(_09581_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15963_ (.A1(_09581_),
    .A2(_08909_),
    .Z(_09582_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15964_ (.A1(_08280_),
    .A2(_09582_),
    .ZN(_09583_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15965_ (.A1(\cs_registers_i.mhpmcounter[1863] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .ZN(_09584_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15966_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .ZN(_09585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15967_ (.I(_08313_),
    .ZN(_09586_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15968_ (.A1(_09586_),
    .A2(_08335_),
    .ZN(_09587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _15969_ (.A1(_09587_),
    .A2(_09582_),
    .ZN(_09588_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15970_ (.A1(_09583_),
    .A2(_09584_),
    .B1(_09585_),
    .B2(_09588_),
    .ZN(_09589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15971_ (.A1(_09580_),
    .A2(_09589_),
    .ZN(_09590_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15972_ (.A1(_09570_),
    .A2(_09576_),
    .A3(_09579_),
    .A4(_09590_),
    .Z(_09591_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15973_ (.I(_09591_),
    .ZN(_09592_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _15974_ (.A1(_11148_[0]),
    .A2(_09547_),
    .B1(_09592_),
    .B2(_11449_[0]),
    .ZN(_09593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15975_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(_09542_),
    .Z(_09594_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15976_ (.A1(_08995_),
    .A2(_09469_),
    .A3(_09594_),
    .Z(_09595_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15977_ (.A1(_08990_),
    .A2(_09595_),
    .B(_08992_),
    .ZN(_09596_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15978_ (.A1(_08997_),
    .A2(_09595_),
    .Z(_09597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15979_ (.I0(_09596_),
    .I1(_09597_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .Z(_09598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15980_ (.A1(_09000_),
    .A2(_09593_),
    .B(_09598_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15981_ (.A1(_08990_),
    .A2(_09069_),
    .B(_09178_),
    .ZN(_09599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15982_ (.I0(_09599_),
    .I1(_09070_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .Z(_09600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15983_ (.A1(_09003_),
    .A2(_09491_),
    .B(_09600_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15984_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11457_[0]),
    .Z(_09601_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15985_ (.A1(\cs_registers_i.mhpmcounter[1864] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .ZN(_09602_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15986_ (.A1(\cs_registers_i.mhpmcounter[1896] ),
    .A2(net3210),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .ZN(_09603_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15987_ (.A1(_08912_),
    .A2(_09602_),
    .B1(_09603_),
    .B2(_08910_),
    .ZN(_09604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15988_ (.A1(_08906_),
    .A2(_09604_),
    .ZN(_09605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15989_ (.A1(\cs_registers_i.csr_mtvec_o[8] ),
    .A2(_08926_),
    .ZN(_09606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15990_ (.A1(\cs_registers_i.dscratch1_q[8] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[8] ),
    .C1(net92),
    .C2(_08935_),
    .ZN(_09607_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15991_ (.A1(\cs_registers_i.dcsr_q[8] ),
    .A2(_08893_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[8] ),
    .ZN(_09608_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15992_ (.A1(_09089_),
    .A2(_09607_),
    .A3(_09608_),
    .Z(_09609_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15993_ (.A1(\cs_registers_i.dscratch0_q[8] ),
    .A2(_08928_),
    .B1(_08938_),
    .B2(\cs_registers_i.mtval_q[8] ),
    .C1(\cs_registers_i.mscratch_q[8] ),
    .C2(_08899_),
    .ZN(_09610_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _15994_ (.A1(_09605_),
    .A2(_09606_),
    .A3(_09609_),
    .A4(_09610_),
    .Z(_09611_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15995_ (.A1(_11461_[0]),
    .A2(_09611_),
    .ZN(_09612_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _15996_ (.A1(_11148_[0]),
    .A2(_09601_),
    .B(_09612_),
    .ZN(_09613_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _15997_ (.A1(_09370_),
    .A2(_09594_),
    .Z(_09614_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3150 (.I(net3149),
    .Z(net3150));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15999_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A3(_09614_),
    .Z(_09616_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16000_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(_09614_),
    .B(_09000_),
    .C(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .ZN(_09617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16001_ (.A1(_09000_),
    .A2(_09613_),
    .B(_09616_),
    .C(_09617_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16002_ (.I0(_11151_[0]),
    .I1(_06849_),
    .S(_11465_[0]),
    .Z(_09618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16003_ (.A1(\cs_registers_i.mhpmcounter[1865] ),
    .A2(_08897_),
    .B1(net3208),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .ZN(_09619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16004_ (.A1(\cs_registers_i.mhpmcounter[1897] ),
    .A2(net3210),
    .B1(_08959_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .ZN(_09620_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16005_ (.A1(_08912_),
    .A2(_09619_),
    .B1(_09620_),
    .B2(_08910_),
    .ZN(_09621_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16006_ (.A1(\cs_registers_i.csr_mtvec_o[9] ),
    .A2(_08926_),
    .B1(_08906_),
    .B2(_09621_),
    .ZN(_09622_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _16007_ (.A1(\cs_registers_i.dscratch0_q[9] ),
    .A2(_08928_),
    .B1(_08932_),
    .B2(\cs_registers_i.csr_mepc_o[9] ),
    .C1(\cs_registers_i.mscratch_q[9] ),
    .C2(_08899_),
    .ZN(_09623_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _16008_ (.A1(\cs_registers_i.dscratch1_q[9] ),
    .A2(_08940_),
    .B1(_09018_),
    .B2(\cs_registers_i.csr_depc_o[9] ),
    .C1(net93),
    .C2(_08935_),
    .ZN(_09624_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16009_ (.A1(\cs_registers_i.mtval_q[9] ),
    .A2(_08938_),
    .B(_08924_),
    .ZN(_09625_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16010_ (.A1(_09622_),
    .A2(_09623_),
    .A3(_09624_),
    .A4(_09625_),
    .Z(_09626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16011_ (.A1(_11469_[0]),
    .A2(_09626_),
    .ZN(_09627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _16012_ (.A1(_11148_[0]),
    .A2(_09618_),
    .B(_09627_),
    .ZN(_09628_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16013_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(_09000_),
    .ZN(_09629_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16014_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A3(_09597_),
    .Z(_09630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16015_ (.I0(_09629_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .S(_09630_),
    .Z(_09631_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16016_ (.A1(_09000_),
    .A2(_09628_),
    .B(_09631_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16017_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A4(_09614_),
    .Z(_09632_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16018_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A2(_09000_),
    .A3(_09632_),
    .Z(_09633_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16019_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .Z(_09634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16020_ (.A1(_09000_),
    .A2(_09029_),
    .B1(_09614_),
    .B2(_09634_),
    .ZN(_09635_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16021_ (.A1(_09633_),
    .A2(_09635_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16022_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(_09000_),
    .ZN(_09636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16023_ (.A1(_09597_),
    .A2(_09634_),
    .ZN(_09637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16024_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .I1(_09636_),
    .S(_09637_),
    .Z(_09638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16025_ (.A1(_09000_),
    .A2(_09066_),
    .B(_09638_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16026_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(_09000_),
    .ZN(_09639_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16027_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(_09614_),
    .A3(_09634_),
    .Z(_09640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16028_ (.I0(_09639_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .S(_09640_),
    .Z(_09641_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16029_ (.A1(_09000_),
    .A2(_09096_),
    .B(_09641_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16030_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A3(_09634_),
    .Z(_09642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16031_ (.A1(_09597_),
    .A2(_09642_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .C(_09000_),
    .ZN(_09643_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16032_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .A2(_09642_),
    .Z(_09644_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16033_ (.A1(_09597_),
    .A2(_09644_),
    .Z(_09645_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16034_ (.A1(_09000_),
    .A2(_09117_),
    .B(_09643_),
    .C(_09645_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16035_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(_09614_),
    .A3(_09644_),
    .Z(_09646_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16036_ (.A1(_09614_),
    .A2(_09644_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .C(_09000_),
    .ZN(_09647_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16037_ (.A1(_09000_),
    .A2(_09133_),
    .B(_09646_),
    .C(_09647_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16038_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(_09000_),
    .ZN(_09648_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16039_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(_09644_),
    .Z(_09649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16040_ (.A1(_09597_),
    .A2(_09649_),
    .ZN(_09650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16041_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .I1(_09648_),
    .S(_09650_),
    .Z(_09651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16042_ (.A1(_09000_),
    .A2(_09149_),
    .B(_09651_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16043_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(_09649_),
    .Z(_09652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16044_ (.A1(_09614_),
    .A2(_09652_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .C(_09000_),
    .ZN(_09653_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16045_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(_09652_),
    .Z(_09654_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16046_ (.A1(_09614_),
    .A2(_09654_),
    .Z(_09655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16047_ (.A1(_09000_),
    .A2(_09174_),
    .B(_09653_),
    .C(_09655_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16048_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .ZN(_09656_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16049_ (.A1(_09469_),
    .A2(_09594_),
    .A3(_09654_),
    .Z(_09657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16050_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .I1(_09656_),
    .S(_09657_),
    .Z(_09658_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16051_ (.A1(_08963_),
    .A2(_08989_),
    .B(_09030_),
    .ZN(_09659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16052_ (.A1(_08997_),
    .A2(_09658_),
    .B1(_09659_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .ZN(_09660_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16053_ (.A1(_09178_),
    .A2(_09194_),
    .B(_09660_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16054_ (.A1(_08995_),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A3(_09031_),
    .Z(_09661_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16055_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .A2(_09661_),
    .Z(_09662_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16056_ (.I(_09508_),
    .ZN(_09663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16057_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .I1(_09663_),
    .S(_08910_),
    .Z(_09664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16058_ (.I0(_09662_),
    .I1(_09664_),
    .S(_08990_),
    .Z(_00060_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16059_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .A2(_09654_),
    .Z(_09665_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16060_ (.A1(_09614_),
    .A2(_09665_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .C(_09000_),
    .ZN(_09666_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16061_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .A2(_09665_),
    .Z(_09667_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16062_ (.A1(_09614_),
    .A2(_09667_),
    .Z(_09668_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16063_ (.A1(_09000_),
    .A2(_09210_),
    .B(_09666_),
    .C(_09668_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16064_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .A2(_09667_),
    .Z(_09669_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16065_ (.A1(_09595_),
    .A2(_09667_),
    .ZN(_09670_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16066_ (.A1(_08997_),
    .A2(_09670_),
    .ZN(_09671_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16067_ (.A1(_08992_),
    .A2(_09671_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .ZN(_09672_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16068_ (.A1(_09000_),
    .A2(_09229_),
    .B1(_09597_),
    .B2(_09669_),
    .C(_09672_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16069_ (.A1(_09176_),
    .A2(_09349_),
    .A3(_09594_),
    .A4(_09669_),
    .ZN(_09673_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16070_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_09673_),
    .B(_08997_),
    .ZN(_09674_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16071_ (.A1(_08992_),
    .A2(_09674_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .ZN(_09675_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16072_ (.A1(_09176_),
    .A2(_09349_),
    .A3(_09594_),
    .A4(_09669_),
    .Z(_09676_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16073_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(_09030_),
    .A3(_09676_),
    .Z(_09677_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16074_ (.A1(_09000_),
    .A2(_09262_),
    .B(_09675_),
    .C(_09677_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16075_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .A2(_09000_),
    .ZN(_09678_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16076_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(_09469_),
    .A3(_09594_),
    .A4(_09669_),
    .Z(_09679_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16077_ (.A1(_09030_),
    .A2(_09679_),
    .ZN(_09680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16078_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .I1(_09678_),
    .S(_09680_),
    .Z(_09681_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16079_ (.A1(_09000_),
    .A2(_09277_),
    .B(_09681_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16080_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .Z(_09682_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16081_ (.A1(_09676_),
    .A2(_09682_),
    .Z(_09683_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16082_ (.A1(_08995_),
    .A2(_09683_),
    .B(_08990_),
    .ZN(_09684_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16083_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(_09003_),
    .A3(_09684_),
    .Z(_09685_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16084_ (.A1(_09030_),
    .A2(_09683_),
    .ZN(_09686_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16085_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(_09686_),
    .ZN(_09687_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16086_ (.A1(_09000_),
    .A2(_09293_),
    .B1(_09685_),
    .B2(_09687_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16087_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A2(_09000_),
    .ZN(_09688_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16088_ (.A1(_09469_),
    .A2(_09594_),
    .A3(_09669_),
    .A4(_09682_),
    .Z(_09689_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16089_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(_09030_),
    .A3(_09689_),
    .Z(_09690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16090_ (.I0(_09688_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .S(_09690_),
    .Z(_09691_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16091_ (.A1(_09000_),
    .A2(_09310_),
    .B(_09691_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16092_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(_09000_),
    .ZN(_09692_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16093_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A3(_09030_),
    .A4(_09683_),
    .Z(_09693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16094_ (.I0(_09692_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .S(_09693_),
    .Z(_09694_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16095_ (.A1(_09000_),
    .A2(_09330_),
    .B(_09694_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16096_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .Z(_09695_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16097_ (.A1(_09030_),
    .A2(_09689_),
    .A3(_09695_),
    .ZN(_09696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16098_ (.A1(net3201),
    .A2(_08999_),
    .B1(_09696_),
    .B2(_08997_),
    .ZN(_09697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16099_ (.I0(_09696_),
    .I1(_09697_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .Z(_09698_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16100_ (.A1(_09178_),
    .A2(_09348_),
    .B(_09698_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16101_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(_09695_),
    .Z(_09699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16102_ (.A1(_09683_),
    .A2(_09699_),
    .Z(_09700_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16103_ (.A1(_09030_),
    .A2(_09700_),
    .ZN(_09701_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16104_ (.I(_09700_),
    .ZN(_09702_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16105_ (.A1(_08997_),
    .A2(_09702_),
    .B(_09659_),
    .ZN(_09703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16106_ (.I0(_09701_),
    .I1(_09703_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .Z(_09704_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16107_ (.A1(_09178_),
    .A2(_09367_),
    .B(_09704_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16108_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(_09689_),
    .A3(_09699_),
    .Z(_09705_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16109_ (.A1(_09030_),
    .A2(_09705_),
    .ZN(_09706_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16110_ (.I(_09705_),
    .ZN(_09707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16111_ (.A1(_08997_),
    .A2(_09707_),
    .B(_09659_),
    .ZN(_09708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16112_ (.I0(_09706_),
    .I1(_09708_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .Z(_09709_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16113_ (.A1(_09178_),
    .A2(_09384_),
    .B(_09709_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16114_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .A3(_09069_),
    .Z(_09710_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16115_ (.A1(_08990_),
    .A2(_09710_),
    .Z(_09711_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16116_ (.A1(_09178_),
    .A2(_09711_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .ZN(_09712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16117_ (.A1(_09003_),
    .A2(_09524_),
    .B(_09712_),
    .C(_09071_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16118_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .ZN(_09713_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16119_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A3(_09700_),
    .Z(_09714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16120_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .I1(_09713_),
    .S(_09714_),
    .Z(_09715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16121_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A2(_09659_),
    .B1(_09715_),
    .B2(_08997_),
    .ZN(_09716_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16122_ (.A1(_09178_),
    .A2(_09401_),
    .B(_09716_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16123_ (.A1(_08995_),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A4(_09705_),
    .Z(_09717_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16124_ (.A1(_08990_),
    .A2(_09717_),
    .Z(_09718_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16125_ (.A1(_08992_),
    .A2(_09718_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .ZN(_09719_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16126_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .Z(_09720_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16127_ (.A1(_09030_),
    .A2(_09705_),
    .A3(_09720_),
    .Z(_09721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16128_ (.A1(_09000_),
    .A2(_09419_),
    .B(_09719_),
    .C(_09721_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16129_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(_09700_),
    .A3(_09720_),
    .ZN(_09722_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16130_ (.A1(_08997_),
    .A2(_09722_),
    .Z(_09723_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16131_ (.A1(_09659_),
    .A2(_09723_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .ZN(_09724_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16132_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .A2(_08999_),
    .A3(_09722_),
    .Z(_09725_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16133_ (.A1(_09178_),
    .A2(_09442_),
    .B(_09724_),
    .C(_09725_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16134_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .A2(_09705_),
    .A3(_09720_),
    .ZN(_09726_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16135_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .A2(_08999_),
    .A3(_09726_),
    .Z(_09727_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16136_ (.A1(_08997_),
    .A2(_09726_),
    .Z(_09728_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16137_ (.A1(_09659_),
    .A2(_09728_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .ZN(_09729_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16138_ (.A1(_09178_),
    .A2(_09458_),
    .B(_09727_),
    .C(_09729_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16139_ (.A1(_08995_),
    .A2(_09033_),
    .B(_08990_),
    .ZN(_09730_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16140_ (.A1(_09000_),
    .A2(_09730_),
    .Z(_09731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16141_ (.I0(_09731_),
    .I1(_09034_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .Z(_09732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16142_ (.A1(_09003_),
    .A2(_09541_),
    .B(_09732_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16143_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(_08992_),
    .ZN(_09733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16144_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .A2(_09071_),
    .ZN(_09734_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16145_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .I1(_09733_),
    .S(_09734_),
    .Z(_09735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16146_ (.A1(_08992_),
    .A2(_09593_),
    .B(_09735_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16147_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .A2(_08992_),
    .ZN(_09736_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16148_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A3(_09034_),
    .Z(_09737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16149_ (.I0(_09736_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .S(_09737_),
    .Z(_09738_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16150_ (.A1(_08992_),
    .A2(_09613_),
    .B(_09738_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16151_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .A2(_09003_),
    .ZN(_09739_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16152_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .A4(_09071_),
    .Z(_09740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16153_ (.I0(_09739_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .S(_09740_),
    .Z(_09741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16154_ (.A1(_09003_),
    .A2(_09628_),
    .B(_09741_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16155_ (.A1(_07000_),
    .A2(_06982_),
    .ZN(_09742_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16156_ (.I(_11004_[0]),
    .ZN(_09743_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16157_ (.A1(_09743_),
    .A2(_07004_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16158_ (.A1(net3215),
    .A2(_06993_),
    .B1(_09742_),
    .B2(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16159_ (.A1(_07295_),
    .A2(_01917_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16160_ (.A1(_06974_),
    .A2(_06982_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16161_ (.A1(_01919_),
    .A2(_01916_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16162_ (.I(_06993_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16163_ (.A1(net3215),
    .A2(_07000_),
    .A3(_06982_),
    .A4(_01921_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16164_ (.I(_11010_[0]),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16165_ (.A1(_07000_),
    .A2(_06982_),
    .B(_01923_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16166_ (.A1(_06993_),
    .A2(_01916_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16167_ (.A1(_01922_),
    .A2(_01924_),
    .A3(_01925_),
    .B(_07001_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16168_ (.A1(_01920_),
    .A2(_01926_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16169_ (.A1(_07005_),
    .A2(_06993_),
    .B(_07001_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16170_ (.A1(_06974_),
    .A2(_06982_),
    .A3(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16171_ (.A1(net3215),
    .A2(_07001_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16172_ (.A1(_07000_),
    .A2(_06982_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16173_ (.A1(_11012_[0]),
    .A2(_01929_),
    .B1(_01930_),
    .B2(_01931_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16174_ (.A1(_11139_[0]),
    .A2(_01932_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16175_ (.I0(_01918_),
    .I1(_01927_),
    .S(_01933_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16176_ (.A1(_11141_[0]),
    .A2(_01934_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16177_ (.A1(_08239_),
    .A2(_08241_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16178_ (.A1(_08234_),
    .A2(_08238_),
    .B(_01936_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16179_ (.A1(_08234_),
    .A2(_08238_),
    .A3(_01936_),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16180_ (.A1(net259),
    .A2(_08250_),
    .B(_01918_),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16181_ (.A1(_01920_),
    .A2(_01926_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16182_ (.A1(net259),
    .A2(_08250_),
    .A3(_01940_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16183_ (.A1(_01937_),
    .A2(_01938_),
    .B1(_01939_),
    .B2(_01941_),
    .C(_11141_[0]),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16184_ (.A1(_07295_),
    .A2(_01917_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16185_ (.A1(net259),
    .A2(_08250_),
    .A3(_01943_),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16186_ (.A1(net259),
    .A2(_08250_),
    .B(_01927_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16187_ (.A1(_08243_),
    .A2(_08244_),
    .B1(_01944_),
    .B2(_01945_),
    .C(_11141_[0]),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16188_ (.A1(_01935_),
    .A2(_01942_),
    .A3(_01946_),
    .Z(_01947_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16189_ (.A1(_11010_[0]),
    .A2(_06993_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16190_ (.A1(_07001_),
    .A2(_01948_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16191_ (.A1(_01947_),
    .A2(_01949_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16192_ (.A1(_08442_),
    .A2(_08444_),
    .B(_01950_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16193_ (.A1(_09743_),
    .A2(_07004_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16194_ (.A1(net3215),
    .A2(_11010_[0]),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16195_ (.A1(_01952_),
    .A2(_01953_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16196_ (.A1(_09742_),
    .A2(_01916_),
    .B1(_01954_),
    .B2(_06993_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16197_ (.A1(_01922_),
    .A2(_01924_),
    .B(_07001_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16198_ (.A1(_07295_),
    .A2(_01955_),
    .B(_01956_),
    .C(_01920_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16199_ (.A1(_08442_),
    .A2(_08444_),
    .A3(_01947_),
    .A4(_01957_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16200_ (.A1(_06246_),
    .A2(_08404_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16201_ (.A1(_06782_),
    .A2(_01959_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16202_ (.A1(net261),
    .A2(_01960_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _16203_ (.A1(\cs_registers_i.mcountinhibit_q[2] ),
    .A2(_08364_),
    .A3(_08392_),
    .A4(_08400_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16204_ (.A1(net59),
    .A2(_08395_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16205_ (.A1(\id_stage_i.id_fsm_q ),
    .A2(_01963_),
    .B(_06758_),
    .C(_06345_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16206_ (.A1(_06224_),
    .A2(_08620_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16207_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .A2(_06244_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _16208_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .A3(_08233_),
    .A4(_01966_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16209_ (.A1(_01965_),
    .A2(_01967_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16210_ (.A1(_01959_),
    .A2(_01968_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16211_ (.A1(_06994_),
    .A2(net3374),
    .A3(_01965_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16212_ (.A1(_06758_),
    .A2(_01963_),
    .B(_01967_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16213_ (.A1(\id_stage_i.id_fsm_q ),
    .A2(_08404_),
    .A3(_01970_),
    .A4(_01971_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16214_ (.A1(_01964_),
    .A2(_01969_),
    .A3(_01972_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16215_ (.A1(_06782_),
    .A2(_01973_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16216_ (.A1(_08948_),
    .A2(_08359_),
    .A3(_08404_),
    .A4(_08313_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16217_ (.A1(_08950_),
    .A2(_08337_),
    .A3(_09582_),
    .A4(_01975_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16218_ (.A1(_09574_),
    .A2(_09580_),
    .A3(_01976_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16219_ (.A1(_01974_),
    .A2(_01977_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _16220_ (.A1(\id_stage_i.controller_i.instr_fetch_err_i ),
    .A2(_08376_),
    .A3(_01962_),
    .A4(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _16221_ (.A1(net3091),
    .A2(_01958_),
    .A3(_01961_),
    .B(_01979_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16222_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(_01980_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16223_ (.A1(_09574_),
    .A2(_09580_),
    .A3(_01976_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16224_ (.A1(_09588_),
    .A2(_01982_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16225_ (.I0(_08945_),
    .I1(_01981_),
    .S(_01983_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _16226_ (.A1(_08988_),
    .A2(_08951_),
    .A3(_08897_),
    .A4(_08906_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16227_ (.A1(\id_stage_i.controller_i.instr_fetch_err_i ),
    .A2(_08376_),
    .A3(_01962_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16228_ (.I(_01985_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16229_ (.A1(_01951_),
    .A2(_01958_),
    .A3(_01961_),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16230_ (.A1(_01984_),
    .A2(_01986_),
    .A3(_01987_),
    .A4(_01974_),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3149 (.I(_11265_[0]),
    .Z(net3149));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3148 (.I(_11307_[0]),
    .Z(net3148));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16233_ (.A1(_11163_[0]),
    .A2(\cs_registers_i.mhpmcounter[1858] ),
    .A3(\cs_registers_i.mhpmcounter[1859] ),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16234_ (.A1(\cs_registers_i.mhpmcounter[1860] ),
    .A2(\cs_registers_i.mhpmcounter[1861] ),
    .A3(_01991_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16235_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(\cs_registers_i.mhpmcounter[1863] ),
    .A3(\cs_registers_i.mhpmcounter[1864] ),
    .A4(\cs_registers_i.mhpmcounter[1865] ),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16236_ (.A1(_01992_),
    .A2(_01993_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16237_ (.A1(_09588_),
    .A2(_01982_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16238_ (.A1(_01988_),
    .A2(_01994_),
    .B(_01995_),
    .C(\cs_registers_i.mhpmcounter[1866] ),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3155 (.I(_03391_),
    .Z(net3155));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16240_ (.A1(\cs_registers_i.mhpmcounter[1866] ),
    .A2(_01988_),
    .A3(_01994_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16241_ (.A1(_08988_),
    .A2(_08951_),
    .A3(_08897_),
    .A4(_08906_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16242_ (.A1(_08910_),
    .A2(_01999_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3143 (.I(_11319_[0]),
    .Z(net3143));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16244_ (.A1(_09029_),
    .A2(_02000_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16245_ (.A1(_01996_),
    .A2(_01998_),
    .A3(_02002_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16246_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(\cs_registers_i.mhpmcounter[1857] ),
    .A3(\cs_registers_i.mhpmcounter[1858] ),
    .A4(\cs_registers_i.mhpmcounter[1859] ),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16247_ (.A1(\cs_registers_i.mhpmcounter[1860] ),
    .A2(\cs_registers_i.mhpmcounter[1861] ),
    .A3(_02003_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16248_ (.A1(\cs_registers_i.mhpmcounter[1866] ),
    .A2(_01993_),
    .A3(_02004_),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16249_ (.A1(\cs_registers_i.mhpmcounter[1867] ),
    .A2(_02000_),
    .Z(_02006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16250_ (.A1(_01988_),
    .A2(_02005_),
    .B(_02006_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16251_ (.A1(\cs_registers_i.mhpmcounter[1867] ),
    .A2(_01988_),
    .A3(_02005_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16252_ (.A1(_09066_),
    .A2(_02000_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16253_ (.A1(_02007_),
    .A2(_02008_),
    .A3(_02009_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16254_ (.A1(_08910_),
    .A2(_01999_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3142 (.I(_11324_[0]),
    .Z(net3142));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16256_ (.A1(\cs_registers_i.mhpmcounter[1867] ),
    .A2(\cs_registers_i.mhpmcounter[1866] ),
    .A3(_01993_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16257_ (.A1(_01992_),
    .A2(_02012_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16258_ (.I(_02013_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3147 (.I(_11312_[0]),
    .Z(net3147));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16260_ (.I0(_02014_),
    .I1(_01983_),
    .S(net3085),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16261_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3157 (.I(_11245_[0]),
    .Z(net3157));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _16263_ (.A1(net3091),
    .A2(_01958_),
    .A3(_01961_),
    .B(_01974_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16264_ (.A1(_01999_),
    .A2(_01985_),
    .A3(net3083),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16265_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(_02020_),
    .A3(_02014_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16266_ (.A1(_09096_),
    .A2(_02010_),
    .B(_02017_),
    .C(_02021_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16267_ (.I(\cs_registers_i.mhpmcounter[1869] ),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16268_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(_02004_),
    .A3(_02012_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16269_ (.I0(_02000_),
    .I1(_02023_),
    .S(_01988_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16270_ (.A1(_11498_[0]),
    .A2(_09115_),
    .B(_09105_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16271_ (.A1(_02022_),
    .A2(_02023_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16272_ (.A1(_02025_),
    .A2(_02000_),
    .B1(_01988_),
    .B2(_02026_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16273_ (.A1(_02022_),
    .A2(_02024_),
    .B(_02027_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16274_ (.I(\cs_registers_i.mhpmcounter[1870] ),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16275_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(\cs_registers_i.mhpmcounter[1869] ),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16276_ (.A1(_02013_),
    .A2(_02029_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16277_ (.I0(_02000_),
    .I1(_02030_),
    .S(_01988_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16278_ (.A1(_09132_),
    .A2(_02000_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16279_ (.I(_02030_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16280_ (.A1(\cs_registers_i.mhpmcounter[1870] ),
    .A2(_02020_),
    .A3(_02033_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16281_ (.A1(_02028_),
    .A2(_02031_),
    .B(_02032_),
    .C(_02034_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16282_ (.I(\cs_registers_i.mhpmcounter[1871] ),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16283_ (.A1(\cs_registers_i.mhpmcounter[1870] ),
    .A2(_02004_),
    .A3(_02012_),
    .A4(_02029_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16284_ (.I0(_02000_),
    .I1(_02036_),
    .S(_01988_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16285_ (.I(_09149_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16286_ (.A1(_02035_),
    .A2(_02036_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16287_ (.A1(_02038_),
    .A2(_02000_),
    .B1(_01988_),
    .B2(_02039_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16288_ (.A1(_02035_),
    .A2(_02037_),
    .B(_02040_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_127_clk_i_regs (.I(clknet_6_58__leaf_clk_i_regs),
    .Z(clknet_leaf_127_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16290_ (.A1(_01985_),
    .A2(_02019_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16291_ (.A1(\cs_registers_i.mhpmcounter[1870] ),
    .A2(\cs_registers_i.mhpmcounter[1871] ),
    .A3(_02042_),
    .A4(_02030_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3141 (.I(_11325_[0]),
    .Z(net3141));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16293_ (.A1(\cs_registers_i.mhpmcounter[1872] ),
    .A2(_01977_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16294_ (.A1(_08963_),
    .A2(_01999_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 place3516 (.I(net3513),
    .Z(net3516));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16296_ (.A1(_02028_),
    .A2(_02035_),
    .A3(_02033_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3139 (.I(_11331_[0]),
    .Z(net3139));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16298_ (.A1(_01985_),
    .A2(net3083),
    .A3(_02048_),
    .B(net3194),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16299_ (.A1(_02046_),
    .A2(_02050_),
    .B(\cs_registers_i.mhpmcounter[1872] ),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16300_ (.A1(_09174_),
    .A2(_02000_),
    .B1(_02043_),
    .B2(_02045_),
    .C(_02051_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16301_ (.A1(\cs_registers_i.mhpmcounter[1871] ),
    .A2(\cs_registers_i.mhpmcounter[1872] ),
    .A3(_02042_),
    .A4(_02036_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16302_ (.A1(\cs_registers_i.mhpmcounter[1873] ),
    .A2(_01977_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16303_ (.A1(\cs_registers_i.mhpmcounter[1871] ),
    .A2(\cs_registers_i.mhpmcounter[1872] ),
    .A3(_02036_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16304_ (.A1(_01985_),
    .A2(net3083),
    .A3(_02054_),
    .B(net3194),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16305_ (.A1(_02046_),
    .A2(_02055_),
    .B(\cs_registers_i.mhpmcounter[1873] ),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16306_ (.A1(_09194_),
    .A2(_02000_),
    .B1(_02052_),
    .B2(_02053_),
    .C(_02056_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16307_ (.A1(\cs_registers_i.mhpmcounter[1870] ),
    .A2(\cs_registers_i.mhpmcounter[1871] ),
    .A3(\cs_registers_i.mhpmcounter[1872] ),
    .A4(\cs_registers_i.mhpmcounter[1873] ),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16308_ (.A1(_02029_),
    .A2(_02057_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16309_ (.A1(_02013_),
    .A2(_02058_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16310_ (.I(_02059_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16311_ (.I0(_02060_),
    .I1(_01983_),
    .S(net3085),
    .Z(_02061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16312_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(_02061_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16313_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(_02020_),
    .A3(_02060_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16314_ (.A1(_09210_),
    .A2(_02010_),
    .B(_02062_),
    .C(_02063_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16315_ (.A1(\cs_registers_i.mhpmcounter[1875] ),
    .A2(_02010_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3160 (.I(_11236_[0]),
    .Z(net3160));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3138 (.I(_11336_[0]),
    .Z(net3138));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16318_ (.A1(_02004_),
    .A2(_02012_),
    .A3(_02058_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16319_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(net3084),
    .A3(_01979_),
    .A4(_02067_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16320_ (.I0(\cs_registers_i.mhpmcounter[1875] ),
    .I1(_02064_),
    .S(_02068_),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16321_ (.A1(_09229_),
    .A2(_02010_),
    .B(_02069_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16322_ (.I0(_11164_[0]),
    .I1(\cs_registers_i.mhpmcounter[1857] ),
    .S(_01980_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16323_ (.I0(_09245_),
    .I1(_02070_),
    .S(_01983_),
    .Z(_00091_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16324_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(\cs_registers_i.mhpmcounter[1875] ),
    .A3(_02059_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16325_ (.A1(_01988_),
    .A2(_02071_),
    .B(_01995_),
    .C(\cs_registers_i.mhpmcounter[1876] ),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16326_ (.A1(net3084),
    .A2(_01979_),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16327_ (.A1(\cs_registers_i.mhpmcounter[1876] ),
    .A2(_02073_),
    .A3(_02071_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16328_ (.A1(_09262_),
    .A2(_02000_),
    .B(_02072_),
    .C(_02074_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16329_ (.A1(\cs_registers_i.mhpmcounter[1877] ),
    .A2(_02010_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16330_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(\cs_registers_i.mhpmcounter[1875] ),
    .A3(\cs_registers_i.mhpmcounter[1876] ),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16331_ (.A1(net3084),
    .A2(_01979_),
    .A3(_02067_),
    .A4(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16332_ (.I0(\cs_registers_i.mhpmcounter[1877] ),
    .I1(_02075_),
    .S(_02077_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16333_ (.A1(_09277_),
    .A2(_02010_),
    .B(_02078_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16334_ (.A1(\cs_registers_i.mhpmcounter[1877] ),
    .A2(_02042_),
    .A3(_02059_),
    .A4(_02076_),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16335_ (.A1(\cs_registers_i.mhpmcounter[1878] ),
    .A2(_01977_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16336_ (.A1(\cs_registers_i.mhpmcounter[1877] ),
    .A2(_02059_),
    .A3(_02076_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16337_ (.A1(_01985_),
    .A2(net3083),
    .A3(_02081_),
    .B(net3194),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16338_ (.A1(_02046_),
    .A2(_02082_),
    .B(\cs_registers_i.mhpmcounter[1878] ),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16339_ (.A1(_09293_),
    .A2(_02000_),
    .B1(_02079_),
    .B2(_02080_),
    .C(_02083_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16340_ (.A1(\cs_registers_i.mhpmcounter[1877] ),
    .A2(\cs_registers_i.mhpmcounter[1878] ),
    .A3(_02076_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16341_ (.A1(_02067_),
    .A2(_02084_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16342_ (.I0(_02085_),
    .I1(_01983_),
    .S(net3085),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16343_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(_02086_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16344_ (.I(\cs_registers_i.mhpmcounter[1879] ),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16345_ (.A1(_02088_),
    .A2(_01988_),
    .A3(_02067_),
    .A4(_02084_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16346_ (.A1(_09310_),
    .A2(_02010_),
    .B(_02087_),
    .C(_02089_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16347_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(_02012_),
    .A3(_02058_),
    .A4(_02084_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16348_ (.A1(_01992_),
    .A2(_02090_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16349_ (.I0(_02091_),
    .I1(_01983_),
    .S(net3085),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16350_ (.A1(\cs_registers_i.mhpmcounter[1880] ),
    .A2(_02092_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16351_ (.A1(\cs_registers_i.mhpmcounter[1880] ),
    .A2(net3085),
    .A3(_02091_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16352_ (.A1(_09330_),
    .A2(_01983_),
    .B(_02093_),
    .C(_02094_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16353_ (.I(\cs_registers_i.mhpmcounter[1881] ),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16354_ (.A1(\cs_registers_i.mhpmcounter[1880] ),
    .A2(_02004_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16355_ (.A1(_02090_),
    .A2(_02096_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16356_ (.I0(_02097_),
    .I1(_01995_),
    .S(net3085),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16357_ (.A1(_11594_[0]),
    .A2(_09346_),
    .B(_09335_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16358_ (.A1(_02095_),
    .A2(_02097_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16359_ (.A1(_02099_),
    .A2(_01995_),
    .B1(_02100_),
    .B2(_02073_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16360_ (.A1(_02095_),
    .A2(_02098_),
    .B(_02101_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16361_ (.A1(\cs_registers_i.mhpmcounter[1882] ),
    .A2(_02000_),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16362_ (.I(\cs_registers_i.mhpmcounter[1880] ),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16363_ (.A1(_02103_),
    .A2(_02095_),
    .A3(_01980_),
    .A4(_02091_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16364_ (.I0(\cs_registers_i.mhpmcounter[1882] ),
    .I1(_02102_),
    .S(_02104_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16365_ (.A1(_09367_),
    .A2(_02000_),
    .B(_02105_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16366_ (.A1(\cs_registers_i.mhpmcounter[1881] ),
    .A2(\cs_registers_i.mhpmcounter[1882] ),
    .A3(_02097_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16367_ (.I(_02106_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16368_ (.I0(_02107_),
    .I1(_01983_),
    .S(net3085),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16369_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(_02108_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16370_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(net3085),
    .A3(_02107_),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16371_ (.A1(_09384_),
    .A2(_01983_),
    .B(_02109_),
    .C(_02110_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16372_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(_02012_),
    .A3(_02058_),
    .A4(_02084_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16373_ (.A1(\cs_registers_i.mhpmcounter[1880] ),
    .A2(\cs_registers_i.mhpmcounter[1881] ),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16374_ (.A1(\cs_registers_i.mhpmcounter[1882] ),
    .A2(_01992_),
    .A3(_02111_),
    .A4(_02112_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16375_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(_02042_),
    .A3(_02113_),
    .Z(_02114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16376_ (.A1(\cs_registers_i.mhpmcounter[1884] ),
    .A2(_01977_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16377_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(_02113_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16378_ (.A1(_01985_),
    .A2(net3083),
    .A3(_02116_),
    .B(net3194),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16379_ (.A1(_02046_),
    .A2(_02117_),
    .B(\cs_registers_i.mhpmcounter[1884] ),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16380_ (.A1(_09401_),
    .A2(_02000_),
    .B1(_02114_),
    .B2(_02115_),
    .C(_02118_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16381_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(_02012_),
    .A3(_02058_),
    .A4(_02084_),
    .Z(_02119_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16382_ (.A1(\cs_registers_i.mhpmcounter[1881] ),
    .A2(\cs_registers_i.mhpmcounter[1882] ),
    .A3(_02119_),
    .A4(_02096_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16383_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(\cs_registers_i.mhpmcounter[1884] ),
    .A3(_02120_),
    .Z(_02121_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16384_ (.A1(\cs_registers_i.mhpmcounter[1885] ),
    .A2(_02000_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16385_ (.A1(_01988_),
    .A2(_02121_),
    .B(_02122_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16386_ (.A1(\cs_registers_i.mhpmcounter[1885] ),
    .A2(_01988_),
    .A3(_02121_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16387_ (.A1(_09419_),
    .A2(_02000_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16388_ (.A1(_02123_),
    .A2(_02124_),
    .A3(_02125_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16389_ (.I(_11163_[0]),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16390_ (.A1(_02126_),
    .A2(_01980_),
    .B(_02010_),
    .C(\cs_registers_i.mhpmcounter[1858] ),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16391_ (.A1(_02126_),
    .A2(\cs_registers_i.mhpmcounter[1858] ),
    .A3(_02020_),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16392_ (.A1(_09423_),
    .A2(_01983_),
    .B(_02127_),
    .C(_02128_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16393_ (.I(\cs_registers_i.mhpmcounter[1886] ),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16394_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(\cs_registers_i.mhpmcounter[1884] ),
    .A3(\cs_registers_i.mhpmcounter[1885] ),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16395_ (.A1(_02113_),
    .A2(_02130_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16396_ (.I0(_02000_),
    .I1(_02131_),
    .S(_01988_),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16397_ (.A1(_02129_),
    .A2(_01988_),
    .A3(_02131_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16398_ (.A1(_09428_),
    .A2(_09441_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16399_ (.A1(_02134_),
    .A2(_02000_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16400_ (.A1(_02129_),
    .A2(_02132_),
    .B(_02133_),
    .C(_02135_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16401_ (.I(\cs_registers_i.mhpmcounter[1887] ),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16402_ (.A1(\cs_registers_i.mhpmcounter[1886] ),
    .A2(_02120_),
    .A3(_02130_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16403_ (.I0(_02000_),
    .I1(_02137_),
    .S(_01988_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16404_ (.A1(_02136_),
    .A2(_02137_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16405_ (.A1(_09457_),
    .A2(_02000_),
    .B1(_01988_),
    .B2(_02139_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16406_ (.A1(_02136_),
    .A2(_02138_),
    .B(_02140_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16407_ (.A1(\cs_registers_i.mhpmcounter[1886] ),
    .A2(\cs_registers_i.mhpmcounter[1887] ),
    .A3(_02131_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16408_ (.A1(_01999_),
    .A2(_02141_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16409_ (.A1(_08946_),
    .A2(_08951_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16410_ (.A1(_08897_),
    .A2(_08906_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16411_ (.A1(_02143_),
    .A2(_02144_),
    .A3(_08910_),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _16412_ (.A1(_01999_),
    .A2(_01985_),
    .A3(_02019_),
    .B(_02145_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16413_ (.A1(_02142_),
    .A2(_02146_),
    .B(_08908_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16414_ (.A1(_08985_),
    .A2(_02145_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16415_ (.A1(_08908_),
    .A2(_01988_),
    .A3(_02141_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16416_ (.A1(_02147_),
    .A2(_02148_),
    .A3(_02149_),
    .Z(_00105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16417_ (.I(\cs_registers_i.mhpmcounter[1889] ),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16418_ (.A1(\cs_registers_i.mhpmcounter[1886] ),
    .A2(\cs_registers_i.mhpmcounter[1887] ),
    .A3(_02106_),
    .A4(_02130_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16419_ (.A1(\cs_registers_i.mhpmcounter[1888] ),
    .A2(_02151_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16420_ (.A1(_02150_),
    .A2(_02042_),
    .A3(_01977_),
    .A4(_02152_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16421_ (.A1(_09588_),
    .A2(_01977_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_128_clk_i_regs (.I(clknet_6_58__leaf_clk_i_regs),
    .Z(clknet_leaf_128_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16423_ (.A1(_01980_),
    .A2(_02154_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16424_ (.A1(\cs_registers_i.mhpmcounter[1889] ),
    .A2(_02156_),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_129_clk_i_regs (.I(clknet_6_58__leaf_clk_i_regs),
    .Z(clknet_leaf_129_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _16426_ (.A1(_02150_),
    .A2(_01982_),
    .A3(_02152_),
    .B1(_02154_),
    .B2(_09468_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16427_ (.A1(_02153_),
    .A2(_02157_),
    .A3(_02159_),
    .Z(_00106_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16428_ (.A1(\cs_registers_i.mhpmcounter[1888] ),
    .A2(\cs_registers_i.mhpmcounter[1889] ),
    .A3(_02141_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16429_ (.A1(_01999_),
    .A2(_01985_),
    .A3(_02019_),
    .A4(_02160_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16430_ (.A1(\cs_registers_i.mhpmcounter[1890] ),
    .A2(_02161_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16431_ (.I0(_08984_),
    .I1(_02162_),
    .S(_02145_),
    .Z(_00107_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16432_ (.A1(\cs_registers_i.mhpmcounter[1888] ),
    .A2(\cs_registers_i.mhpmcounter[1889] ),
    .A3(\cs_registers_i.mhpmcounter[1890] ),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16433_ (.A1(_02151_),
    .A2(_02163_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16434_ (.A1(\cs_registers_i.mhpmcounter[1891] ),
    .A2(_01977_),
    .A3(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16435_ (.A1(\cs_registers_i.mhpmcounter[1891] ),
    .A2(_01982_),
    .A3(_02164_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16436_ (.A1(\cs_registers_i.mhpmcounter[1891] ),
    .A2(_02156_),
    .B1(_02166_),
    .B2(_02042_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16437_ (.A1(_09491_),
    .A2(_02154_),
    .B(_02165_),
    .C(_02167_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16438_ (.A1(\cs_registers_i.mhpmcounter[1891] ),
    .A2(_02163_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16439_ (.A1(_02141_),
    .A2(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16440_ (.A1(_01999_),
    .A2(_01985_),
    .A3(_02019_),
    .A4(_02169_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16441_ (.A1(\cs_registers_i.mhpmcounter[1892] ),
    .A2(_02170_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16442_ (.I0(_09663_),
    .I1(_02171_),
    .S(_02145_),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16443_ (.I(\cs_registers_i.mhpmcounter[1893] ),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16444_ (.A1(\cs_registers_i.mhpmcounter[1892] ),
    .A2(_02168_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16445_ (.A1(_02151_),
    .A2(_02173_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16446_ (.A1(_02172_),
    .A2(_01988_),
    .A3(_02174_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16447_ (.A1(\cs_registers_i.mhpmcounter[1893] ),
    .A2(_02156_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _16448_ (.A1(_02172_),
    .A2(_01982_),
    .A3(_02174_),
    .B1(_02154_),
    .B2(_09524_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16449_ (.A1(_02175_),
    .A2(_02176_),
    .A3(_02177_),
    .Z(_00110_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_134_clk_i_regs (.I(clknet_6_58__leaf_clk_i_regs),
    .Z(clknet_leaf_134_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_136_clk_i_regs (.I(clknet_6_58__leaf_clk_i_regs),
    .Z(clknet_leaf_136_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16452_ (.A1(\cs_registers_i.mhpmcounter[1893] ),
    .A2(_02141_),
    .A3(_02173_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16453_ (.A1(_01984_),
    .A2(_02180_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16454_ (.I(\cs_registers_i.mhpmcounter[1894] ),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16455_ (.A1(_02146_),
    .A2(_02181_),
    .B(_02182_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16456_ (.A1(\cs_registers_i.mhpmcounter[1894] ),
    .A2(_02020_),
    .A3(_02180_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16457_ (.A1(_09541_),
    .A2(_02145_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16458_ (.A1(_02183_),
    .A2(_02184_),
    .A3(_02185_),
    .Z(_00111_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_137_clk_i_regs (.I(clknet_6_47__leaf_clk_i_regs),
    .Z(clknet_leaf_137_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16460_ (.A1(\cs_registers_i.mhpmcounter[1893] ),
    .A2(\cs_registers_i.mhpmcounter[1894] ),
    .A3(_02174_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16461_ (.A1(_01982_),
    .A2(_02187_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16462_ (.A1(_02156_),
    .A2(_02188_),
    .B(\cs_registers_i.mhpmcounter[1895] ),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16463_ (.I(\cs_registers_i.mhpmcounter[1895] ),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16464_ (.A1(_02190_),
    .A2(_02073_),
    .A3(_02187_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16465_ (.A1(_09593_),
    .A2(_02154_),
    .B(_02189_),
    .C(_02191_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16466_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(\cs_registers_i.mhpmcounter[1857] ),
    .A3(\cs_registers_i.mhpmcounter[1858] ),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16467_ (.A1(_01985_),
    .A2(net3083),
    .A3(_02192_),
    .B(_01984_),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16468_ (.A1(_02046_),
    .A2(_02193_),
    .B(\cs_registers_i.mhpmcounter[1859] ),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16469_ (.A1(_09491_),
    .A2(_02000_),
    .B1(_01988_),
    .B2(_02003_),
    .C(_02194_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16470_ (.I(\cs_registers_i.mhpmcounter[1896] ),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16471_ (.A1(_02182_),
    .A2(_02190_),
    .A3(_02180_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16472_ (.A1(_02195_),
    .A2(_01988_),
    .A3(_02196_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16473_ (.A1(\cs_registers_i.mhpmcounter[1896] ),
    .A2(_02156_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _16474_ (.A1(_02195_),
    .A2(_01982_),
    .A3(_02196_),
    .B1(_02154_),
    .B2(_09613_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16475_ (.A1(_02197_),
    .A2(_02198_),
    .A3(_02199_),
    .Z(_00114_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16476_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(\cs_registers_i.mhpmcounter[1896] ),
    .A3(_02187_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16477_ (.A1(\cs_registers_i.mhpmcounter[1897] ),
    .A2(_02020_),
    .A3(_02200_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16478_ (.A1(\cs_registers_i.mhpmcounter[1897] ),
    .A2(_02156_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16479_ (.A1(\cs_registers_i.mhpmcounter[1897] ),
    .A2(_01977_),
    .A3(_02200_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16480_ (.A1(_09628_),
    .A2(_02154_),
    .B(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16481_ (.A1(_02201_),
    .A2(_02202_),
    .A3(_02204_),
    .Z(_00115_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16482_ (.A1(\cs_registers_i.mhpmcounter[1896] ),
    .A2(\cs_registers_i.mhpmcounter[1897] ),
    .A3(_02196_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16483_ (.A1(\cs_registers_i.mhpmcounter[1898] ),
    .A2(_01982_),
    .A3(_02205_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16484_ (.A1(\cs_registers_i.mhpmcounter[1898] ),
    .A2(_02156_),
    .B1(_02206_),
    .B2(_02042_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16485_ (.A1(_09588_),
    .A2(_01977_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16486_ (.A1(\cs_registers_i.mhpmcounter[1898] ),
    .A2(_01977_),
    .A3(_02205_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16487_ (.A1(_09028_),
    .A2(_02208_),
    .B(_02209_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16488_ (.A1(_02207_),
    .A2(_02210_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_138_clk_i_regs (.I(clknet_6_47__leaf_clk_i_regs),
    .Z(clknet_leaf_138_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_139_clk_i_regs (.I(clknet_6_58__leaf_clk_i_regs),
    .Z(clknet_leaf_139_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16491_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(\cs_registers_i.mhpmcounter[1896] ),
    .A3(_02187_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16492_ (.A1(\cs_registers_i.mhpmcounter[1897] ),
    .A2(\cs_registers_i.mhpmcounter[1898] ),
    .A3(_02213_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16493_ (.A1(_01999_),
    .A2(_02214_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16494_ (.A1(net3077),
    .A2(_02215_),
    .B(\cs_registers_i.mhpmcounter[1899] ),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16495_ (.A1(_09040_),
    .A2(_09065_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16496_ (.A1(\cs_registers_i.mhpmcounter[1899] ),
    .A2(_02214_),
    .B(_01982_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16497_ (.A1(_02217_),
    .A2(_02208_),
    .B(_02156_),
    .C(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16498_ (.A1(_02216_),
    .A2(_02219_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_141_clk_i_regs (.I(clknet_6_47__leaf_clk_i_regs),
    .Z(clknet_leaf_141_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16500_ (.A1(_09075_),
    .A2(_09095_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16501_ (.A1(_08963_),
    .A2(_02221_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16502_ (.A1(\cs_registers_i.mhpmcounter[1899] ),
    .A2(\cs_registers_i.mhpmcounter[1898] ),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16503_ (.A1(_02205_),
    .A2(_02223_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16504_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(_02224_),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16505_ (.I0(_02222_),
    .I1(_02225_),
    .S(_01984_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16506_ (.A1(_01999_),
    .A2(_02224_),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16507_ (.A1(net3077),
    .A2(_02227_),
    .B(\cs_registers_i.mhpmcounter[1900] ),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16508_ (.A1(net3077),
    .A2(_02226_),
    .B(_02228_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_142_clk_i_regs (.I(clknet_6_47__leaf_clk_i_regs),
    .Z(clknet_leaf_142_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16510_ (.A1(\cs_registers_i.mhpmcounter[1899] ),
    .A2(\cs_registers_i.mhpmcounter[1897] ),
    .A3(\cs_registers_i.mhpmcounter[1898] ),
    .A4(_02213_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16511_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(_02230_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16512_ (.A1(_01984_),
    .A2(_02231_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16513_ (.A1(net3077),
    .A2(_02232_),
    .B(\cs_registers_i.mhpmcounter[1901] ),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16514_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(\cs_registers_i.mhpmcounter[1899] ),
    .A3(\cs_registers_i.mhpmcounter[1901] ),
    .A4(_02214_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16515_ (.A1(_01982_),
    .A2(_02234_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16516_ (.A1(_02025_),
    .A2(_02208_),
    .B(_02156_),
    .C(_02235_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16517_ (.A1(_02233_),
    .A2(_02236_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16518_ (.I(\cs_registers_i.mhpmcounter[1902] ),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16519_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(\cs_registers_i.mhpmcounter[1901] ),
    .A3(_02224_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16520_ (.A1(_02237_),
    .A2(_01977_),
    .A3(_02238_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16521_ (.A1(_09132_),
    .A2(_02208_),
    .B(_02239_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16522_ (.A1(_01982_),
    .A2(_02238_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16523_ (.A1(_02156_),
    .A2(_02241_),
    .B(\cs_registers_i.mhpmcounter[1902] ),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16524_ (.A1(_02156_),
    .A2(_02240_),
    .B(_02242_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16525_ (.A1(\cs_registers_i.mhpmcounter[1902] ),
    .A2(_02234_),
    .B(_01982_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16526_ (.I(\cs_registers_i.mhpmcounter[1903] ),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16527_ (.A1(_02156_),
    .A2(_02243_),
    .B(_02244_),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16528_ (.A1(\cs_registers_i.mhpmcounter[1902] ),
    .A2(\cs_registers_i.mhpmcounter[1903] ),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16529_ (.A1(_02234_),
    .A2(_02246_),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16530_ (.A1(_09149_),
    .A2(_02154_),
    .B1(_02247_),
    .B2(_01982_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16531_ (.A1(_02156_),
    .A2(_02248_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16532_ (.A1(_02245_),
    .A2(_02249_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16533_ (.I(_09174_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16534_ (.A1(_02238_),
    .A2(_02246_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16535_ (.A1(\cs_registers_i.mhpmcounter[1904] ),
    .A2(net3194),
    .A3(_02251_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16536_ (.A1(_02250_),
    .A2(net3194),
    .B(_02252_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16537_ (.A1(_01999_),
    .A2(_02251_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16538_ (.A1(net3077),
    .A2(_02254_),
    .B(\cs_registers_i.mhpmcounter[1904] ),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16539_ (.A1(net3077),
    .A2(_02253_),
    .B(_02255_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16540_ (.A1(\cs_registers_i.mhpmcounter[1904] ),
    .A2(_02247_),
    .B(_01982_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16541_ (.I(\cs_registers_i.mhpmcounter[1905] ),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16542_ (.A1(_02156_),
    .A2(_02256_),
    .B(_02257_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16543_ (.A1(\cs_registers_i.mhpmcounter[1904] ),
    .A2(\cs_registers_i.mhpmcounter[1905] ),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16544_ (.A1(_02247_),
    .A2(_02259_),
    .B(_01982_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16545_ (.A1(_09194_),
    .A2(_02154_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16546_ (.A1(_02156_),
    .A2(_02260_),
    .A3(_02261_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16547_ (.A1(_02258_),
    .A2(_02262_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16548_ (.A1(\cs_registers_i.mhpmcounter[1860] ),
    .A2(_01991_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16549_ (.I(_01991_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16550_ (.A1(_01985_),
    .A2(net3083),
    .A3(_02264_),
    .B(_01984_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16551_ (.A1(_02046_),
    .A2(_02265_),
    .B(\cs_registers_i.mhpmcounter[1860] ),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16552_ (.A1(_09508_),
    .A2(_02000_),
    .B1(_01988_),
    .B2(_02263_),
    .C(_02266_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16553_ (.I(\cs_registers_i.mhpmcounter[1906] ),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16554_ (.A1(_02267_),
    .A2(_01977_),
    .A3(_02251_),
    .A4(_02259_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16555_ (.A1(_02251_),
    .A2(_02259_),
    .B(_02267_),
    .C(_01982_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16556_ (.A1(_02042_),
    .A2(_02268_),
    .B(_02269_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16557_ (.I(_09210_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16558_ (.A1(_02271_),
    .A2(_02208_),
    .B1(_02156_),
    .B2(\cs_registers_i.mhpmcounter[1906] ),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16559_ (.A1(_02270_),
    .A2(_02272_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16560_ (.A1(\cs_registers_i.mhpmcounter[1906] ),
    .A2(\cs_registers_i.mhpmcounter[1907] ),
    .A3(_02259_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16561_ (.A1(_02247_),
    .A2(_02273_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16562_ (.A1(_01982_),
    .A2(_02274_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16563_ (.A1(_01986_),
    .A2(net3084),
    .A3(_01974_),
    .A4(_02275_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16564_ (.A1(_11546_[0]),
    .A2(_09227_),
    .B(_09216_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16565_ (.A1(_02277_),
    .A2(_02208_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16566_ (.A1(_02156_),
    .A2(_02276_),
    .A3(_02278_),
    .B(\cs_registers_i.mhpmcounter[1907] ),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16567_ (.A1(\cs_registers_i.mhpmcounter[1906] ),
    .A2(_02247_),
    .A3(_02259_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16568_ (.A1(_02276_),
    .A2(_02278_),
    .B1(_02280_),
    .B2(_01982_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16569_ (.A1(_02279_),
    .A2(_02281_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16570_ (.I(_09262_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16571_ (.A1(\cs_registers_i.mhpmcounter[1908] ),
    .A2(_02273_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16572_ (.A1(net3194),
    .A2(_02251_),
    .A3(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16573_ (.A1(_02282_),
    .A2(net3194),
    .B(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16574_ (.A1(_02251_),
    .A2(_02273_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16575_ (.A1(net3194),
    .A2(_02286_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16576_ (.A1(net3077),
    .A2(_02287_),
    .B(\cs_registers_i.mhpmcounter[1908] ),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16577_ (.A1(net3077),
    .A2(_02285_),
    .B(_02288_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16578_ (.A1(\cs_registers_i.mhpmcounter[1908] ),
    .A2(_02274_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16579_ (.A1(net3085),
    .A2(_02289_),
    .B(_02154_),
    .C(\cs_registers_i.mhpmcounter[1909] ),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16580_ (.A1(\cs_registers_i.mhpmcounter[1909] ),
    .A2(net3085),
    .A3(_02208_),
    .A4(_02289_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16581_ (.A1(_02290_),
    .A2(_02291_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16582_ (.A1(_09588_),
    .A2(_09277_),
    .A3(_01977_),
    .B(_02292_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16583_ (.A1(\cs_registers_i.mhpmcounter[1909] ),
    .A2(_02251_),
    .A3(_02283_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16584_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(_02293_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16585_ (.I0(_09293_),
    .I1(_02294_),
    .S(net3194),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16586_ (.A1(_01999_),
    .A2(_02293_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16587_ (.A1(net3077),
    .A2(_02296_),
    .B(\cs_registers_i.mhpmcounter[1910] ),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16588_ (.A1(net3077),
    .A2(_02295_),
    .B(_02297_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16589_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(\cs_registers_i.mhpmcounter[1901] ),
    .A3(_02230_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16590_ (.A1(\cs_registers_i.mhpmcounter[1909] ),
    .A2(_02298_),
    .A3(_02246_),
    .A4(_02283_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16591_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(\cs_registers_i.mhpmcounter[1911] ),
    .A3(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16592_ (.A1(_09310_),
    .A2(_02046_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16593_ (.A1(net3194),
    .A2(_02300_),
    .B(_02301_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16594_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(_02299_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16595_ (.A1(net3194),
    .A2(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16596_ (.A1(net3077),
    .A2(_02304_),
    .B(\cs_registers_i.mhpmcounter[1911] ),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16597_ (.A1(net3077),
    .A2(_02302_),
    .B(_02305_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16598_ (.I(_09330_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16599_ (.A1(_08963_),
    .A2(_02306_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16600_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(\cs_registers_i.mhpmcounter[1911] ),
    .A3(\cs_registers_i.mhpmcounter[1912] ),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16601_ (.A1(_02293_),
    .A2(_02308_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16602_ (.I0(_02307_),
    .I1(_02309_),
    .S(net3194),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16603_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(\cs_registers_i.mhpmcounter[1911] ),
    .A3(_02293_),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16604_ (.A1(_01999_),
    .A2(_02311_),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16605_ (.A1(net3077),
    .A2(_02312_),
    .B(\cs_registers_i.mhpmcounter[1912] ),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16606_ (.A1(net3077),
    .A2(_02310_),
    .B(_02313_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16607_ (.A1(\cs_registers_i.mhpmcounter[1913] ),
    .A2(_02299_),
    .A3(_02308_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16608_ (.I0(_09348_),
    .I1(_02314_),
    .S(net3194),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16609_ (.A1(_02299_),
    .A2(_02308_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16610_ (.A1(net3194),
    .A2(_02316_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16611_ (.A1(net3077),
    .A2(_02317_),
    .B(\cs_registers_i.mhpmcounter[1913] ),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16612_ (.A1(net3077),
    .A2(_02315_),
    .B(_02318_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16613_ (.A1(\cs_registers_i.mhpmcounter[1913] ),
    .A2(\cs_registers_i.mhpmcounter[1914] ),
    .A3(_02308_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16614_ (.A1(_02293_),
    .A2(_02319_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _16615_ (.I(_09367_),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16616_ (.A1(_08963_),
    .A2(_02321_),
    .A3(_01999_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16617_ (.A1(net3194),
    .A2(_02320_),
    .B(_02322_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16618_ (.A1(\cs_registers_i.mhpmcounter[1913] ),
    .A2(_02293_),
    .A3(_02308_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16619_ (.A1(_01999_),
    .A2(_02324_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16620_ (.A1(net3077),
    .A2(_02325_),
    .B(\cs_registers_i.mhpmcounter[1914] ),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16621_ (.A1(net3077),
    .A2(_02323_),
    .B(_02326_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16622_ (.I(\cs_registers_i.mhpmcounter[1915] ),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16623_ (.A1(_02299_),
    .A2(_02319_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16624_ (.A1(_01999_),
    .A2(_02328_),
    .B(net3077),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _16625_ (.I(_09384_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16626_ (.A1(net3194),
    .A2(_02328_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16627_ (.A1(_02330_),
    .A2(net3194),
    .B1(_02331_),
    .B2(_02327_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16628_ (.A1(_02327_),
    .A2(_02329_),
    .B1(_02332_),
    .B2(net3077),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16629_ (.I(\cs_registers_i.mhpmcounter[1861] ),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16630_ (.I0(_02333_),
    .I1(_02004_),
    .S(_02042_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16631_ (.A1(\cs_registers_i.mhpmcounter[1860] ),
    .A2(_02003_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16632_ (.A1(_01984_),
    .A2(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16633_ (.A1(_02046_),
    .A2(_02336_),
    .B(\cs_registers_i.mhpmcounter[1861] ),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16634_ (.A1(_09524_),
    .A2(_01995_),
    .B1(_02334_),
    .B2(_01984_),
    .C(_02337_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16635_ (.A1(_11618_[0]),
    .A2(_09399_),
    .B(_09388_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16636_ (.A1(_01999_),
    .A2(_02320_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16637_ (.A1(\cs_registers_i.mhpmcounter[1915] ),
    .A2(\cs_registers_i.mhpmcounter[1916] ),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16638_ (.A1(_02338_),
    .A2(net3194),
    .B1(_02339_),
    .B2(_02340_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16639_ (.A1(_02327_),
    .A2(_02320_),
    .B(net3194),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16640_ (.A1(net3077),
    .A2(_02342_),
    .B(\cs_registers_i.mhpmcounter[1916] ),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16641_ (.A1(net3077),
    .A2(_02341_),
    .B(_02343_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16642_ (.A1(_11626_[0]),
    .A2(_09417_),
    .B(_09406_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16643_ (.A1(\cs_registers_i.mhpmcounter[1915] ),
    .A2(\cs_registers_i.mhpmcounter[1916] ),
    .A3(\cs_registers_i.mhpmcounter[1917] ),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16644_ (.A1(_02344_),
    .A2(net3194),
    .B1(_02331_),
    .B2(_02345_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16645_ (.A1(\cs_registers_i.mhpmcounter[1915] ),
    .A2(\cs_registers_i.mhpmcounter[1916] ),
    .A3(_02328_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16646_ (.A1(_01999_),
    .A2(_02347_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16647_ (.A1(net3077),
    .A2(_02348_),
    .B(\cs_registers_i.mhpmcounter[1917] ),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16648_ (.A1(net3077),
    .A2(_02346_),
    .B(_02349_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16649_ (.A1(\cs_registers_i.mhpmcounter[1915] ),
    .A2(\cs_registers_i.mhpmcounter[1916] ),
    .A3(\cs_registers_i.mhpmcounter[1917] ),
    .A4(\cs_registers_i.mhpmcounter[1918] ),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16650_ (.I(_02350_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16651_ (.A1(_02134_),
    .A2(net3194),
    .B1(_02339_),
    .B2(_02351_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16652_ (.A1(_02320_),
    .A2(_02345_),
    .B(net3194),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16653_ (.A1(net3077),
    .A2(_02353_),
    .B(\cs_registers_i.mhpmcounter[1918] ),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16654_ (.A1(net3077),
    .A2(_02352_),
    .B(_02354_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16655_ (.A1(_08963_),
    .A2(_09457_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16656_ (.A1(\cs_registers_i.mhpmcounter[1919] ),
    .A2(_02328_),
    .A3(_02350_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16657_ (.I0(_02355_),
    .I1(_02356_),
    .S(net3194),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16658_ (.A1(_02328_),
    .A2(_02350_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16659_ (.A1(net3194),
    .A2(_02358_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16660_ (.A1(net3077),
    .A2(_02359_),
    .B(\cs_registers_i.mhpmcounter[1919] ),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16661_ (.A1(net3077),
    .A2(_02357_),
    .B(_02360_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16662_ (.I(_01992_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16663_ (.A1(_01985_),
    .A2(net3083),
    .A3(_02361_),
    .B(_01984_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16664_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(_02046_),
    .A3(_02362_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16665_ (.A1(_01988_),
    .A2(_01992_),
    .B(\cs_registers_i.mhpmcounter[1862] ),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16666_ (.A1(_09541_),
    .A2(_02010_),
    .B1(_02363_),
    .B2(_02364_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16667_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(_02004_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16668_ (.A1(\cs_registers_i.mhpmcounter[1863] ),
    .A2(_02010_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16669_ (.A1(_01988_),
    .A2(_02365_),
    .B(_02366_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16670_ (.A1(_09593_),
    .A2(_02010_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16671_ (.I(\cs_registers_i.mhpmcounter[1863] ),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16672_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(_02369_),
    .A3(_01988_),
    .A4(_02004_),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16673_ (.A1(_02367_),
    .A2(_02368_),
    .A3(_02370_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16674_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(\cs_registers_i.mhpmcounter[1863] ),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16675_ (.A1(_01992_),
    .A2(_02371_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16676_ (.A1(\cs_registers_i.mhpmcounter[1864] ),
    .A2(_02000_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16677_ (.A1(_01988_),
    .A2(_02372_),
    .B(_02373_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16678_ (.A1(\cs_registers_i.mhpmcounter[1864] ),
    .A2(_01988_),
    .A3(_01992_),
    .A4(_02371_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16679_ (.A1(_09613_),
    .A2(_02000_),
    .B(_02374_),
    .C(_02375_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16680_ (.A1(_01993_),
    .A2(_02004_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16681_ (.A1(\cs_registers_i.mhpmcounter[1864] ),
    .A2(_02371_),
    .A3(_02004_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16682_ (.A1(_01985_),
    .A2(net3083),
    .A3(_02377_),
    .B(_01984_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16683_ (.A1(_02046_),
    .A2(_02378_),
    .B(\cs_registers_i.mhpmcounter[1865] ),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16684_ (.A1(_09628_),
    .A2(_02000_),
    .B1(_01988_),
    .B2(_02376_),
    .C(_02379_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _16685_ (.A1(_08391_),
    .A2(_08664_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16686_ (.A1(\cs_registers_i.dcsr_q[0] ),
    .A2(_08380_),
    .B1(_08385_),
    .B2(\cs_registers_i.mstatus_q[2] ),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16687_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_08660_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16688_ (.I0(_08724_),
    .I1(_02382_),
    .S(_08632_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16689_ (.A1(_08370_),
    .A2(_02383_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _16690_ (.A1(_08629_),
    .A2(_08636_),
    .B(_02384_),
    .C(_08662_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16691_ (.A1(_08380_),
    .A2(_08385_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16692_ (.A1(_08665_),
    .A2(_02386_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16693_ (.A1(\cs_registers_i.priv_mode_id_o[0] ),
    .A2(_02385_),
    .B(_02387_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16694_ (.A1(_02380_),
    .A2(_02381_),
    .B(_02388_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16695_ (.A1(\cs_registers_i.dcsr_q[1] ),
    .A2(_08380_),
    .B1(_08385_),
    .B2(\cs_registers_i.mstatus_q[3] ),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16696_ (.A1(\cs_registers_i.priv_mode_id_o[1] ),
    .A2(_02385_),
    .B(_02387_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16697_ (.A1(_02380_),
    .A2(_02389_),
    .B(_02390_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16698_ (.I(\cs_registers_i.dcsr_q[0] ),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16699_ (.A1(_08946_),
    .A2(_08951_),
    .A3(_08893_),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16700_ (.A1(_02391_),
    .A2(_02392_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16701_ (.A1(_08945_),
    .A2(_09245_),
    .A3(_02392_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16702_ (.A1(_02393_),
    .A2(_02394_),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16703_ (.A1(_08389_),
    .A2(_08657_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16704_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_08370_),
    .A3(_08632_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _16705_ (.A1(_02396_),
    .A2(_02397_),
    .B(_08681_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _16706_ (.I(_02398_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16707_ (.I0(\cs_registers_i.priv_mode_id_o[0] ),
    .I1(_02395_),
    .S(_02399_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16708_ (.I0(_02217_),
    .I1(\cs_registers_i.dcsr_q[11] ),
    .S(_02392_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16709_ (.I0(_02221_),
    .I1(\cs_registers_i.dcsr_q[12] ),
    .S(_02392_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16710_ (.I0(_02025_),
    .I1(\cs_registers_i.dcsr_q[13] ),
    .S(_02392_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16711_ (.I0(_02038_),
    .I1(\cs_registers_i.dcsr_q[15] ),
    .S(_02392_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16712_ (.I(\cs_registers_i.dcsr_q[1] ),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16713_ (.A1(_02400_),
    .A2(_02392_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16714_ (.A1(_02394_),
    .A2(_02401_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16715_ (.I0(\cs_registers_i.priv_mode_id_o[1] ),
    .I1(_02402_),
    .S(_02399_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16716_ (.I0(_08984_),
    .I1(\cs_registers_i.dcsr_q[2] ),
    .S(_02392_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16717_ (.I(\cs_registers_i.dcsr_q[6] ),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16718_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_08661_),
    .B1(_02399_),
    .B2(_02403_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16719_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_02399_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16720_ (.I(\cs_registers_i.dcsr_q[2] ),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16721_ (.A1(_02405_),
    .A2(net60),
    .A3(_08661_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16722_ (.A1(_02404_),
    .A2(_02406_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16723_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_08661_),
    .B1(_02399_),
    .B2(\cs_registers_i.dcsr_q[8] ),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16724_ (.I(_02407_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16725_ (.A1(_08946_),
    .A2(_08951_),
    .A3(_09018_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_143_clk_i_regs (.I(clknet_6_47__leaf_clk_i_regs),
    .Z(clknet_leaf_143_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16727_ (.A1(_02399_),
    .A2(_02408_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_145_clk_i_regs (.I(clknet_6_46__leaf_clk_i_regs),
    .Z(clknet_leaf_145_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16729_ (.A1(\cs_registers_i.csr_depc_o[10] ),
    .A2(_02410_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3554 (.I(net3553),
    .Z(net3554));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place3515 (.I(net314),
    .Z(net3515));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16732_ (.I0(\cs_registers_i.pc_if_i[10] ),
    .I1(\cs_registers_i.pc_id_i[10] ),
    .S(_08662_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16733_ (.A1(net3290),
    .A2(_02415_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16734_ (.A1(_09029_),
    .A2(_02408_),
    .B(_02412_),
    .C(_02416_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_147_clk_i_regs (.I(clknet_6_46__leaf_clk_i_regs),
    .Z(clknet_leaf_147_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16736_ (.I0(\cs_registers_i.pc_if_i[11] ),
    .I1(\cs_registers_i.pc_id_i[11] ),
    .S(_08662_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16737_ (.A1(_02398_),
    .A2(_02418_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16738_ (.A1(\cs_registers_i.csr_depc_o[11] ),
    .A2(_02410_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16739_ (.A1(_09066_),
    .A2(_02408_),
    .B(_02419_),
    .C(_02420_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16740_ (.I0(\cs_registers_i.pc_if_i[12] ),
    .I1(\cs_registers_i.pc_id_i[12] ),
    .S(_08662_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16741_ (.A1(net3290),
    .A2(_02421_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16742_ (.A1(\cs_registers_i.csr_depc_o[12] ),
    .A2(_02410_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16743_ (.A1(_09096_),
    .A2(_02408_),
    .B(_02422_),
    .C(_02423_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16744_ (.I0(\cs_registers_i.pc_if_i[13] ),
    .I1(\cs_registers_i.pc_id_i[13] ),
    .S(_08662_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16745_ (.A1(net3290),
    .A2(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16746_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(_02410_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16747_ (.A1(_09117_),
    .A2(_02408_),
    .B(_02425_),
    .C(_02426_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16748_ (.I0(\cs_registers_i.pc_if_i[14] ),
    .I1(\cs_registers_i.pc_id_i[14] ),
    .S(net3291),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16749_ (.A1(net3290),
    .A2(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16750_ (.A1(\cs_registers_i.csr_depc_o[14] ),
    .A2(_02410_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16751_ (.A1(_09133_),
    .A2(_02408_),
    .B(_02428_),
    .C(_02429_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16752_ (.I0(\cs_registers_i.pc_if_i[15] ),
    .I1(\cs_registers_i.pc_id_i[15] ),
    .S(_08662_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16753_ (.A1(net3290),
    .A2(_02430_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16754_ (.A1(\cs_registers_i.csr_depc_o[15] ),
    .A2(_02410_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16755_ (.A1(_09149_),
    .A2(_02408_),
    .B(_02431_),
    .C(_02432_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3128 (.I(_03700_),
    .Z(net3128));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16757_ (.I0(\cs_registers_i.pc_if_i[16] ),
    .I1(\cs_registers_i.pc_id_i[16] ),
    .S(net3291),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16758_ (.A1(net3290),
    .A2(_02434_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16759_ (.A1(\cs_registers_i.csr_depc_o[16] ),
    .A2(_02410_),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16760_ (.A1(_09174_),
    .A2(_02408_),
    .B(_02435_),
    .C(_02436_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16761_ (.I0(\cs_registers_i.pc_if_i[17] ),
    .I1(\cs_registers_i.pc_id_i[17] ),
    .S(net3291),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16762_ (.A1(net3290),
    .A2(_02437_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16763_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(_02410_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16764_ (.A1(_09194_),
    .A2(_02408_),
    .B(_02438_),
    .C(_02439_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16765_ (.I0(\cs_registers_i.pc_if_i[18] ),
    .I1(\cs_registers_i.pc_id_i[18] ),
    .S(net3291),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16766_ (.A1(net3290),
    .A2(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16767_ (.A1(\cs_registers_i.csr_depc_o[18] ),
    .A2(_02410_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16768_ (.A1(_09210_),
    .A2(_02408_),
    .B(_02441_),
    .C(_02442_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16769_ (.I0(\cs_registers_i.pc_if_i[19] ),
    .I1(\cs_registers_i.pc_id_i[19] ),
    .S(net3291),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16770_ (.A1(net3290),
    .A2(_02443_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3553 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(net3553));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16772_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(_02410_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16773_ (.A1(_09229_),
    .A2(_02408_),
    .B(_02444_),
    .C(_02446_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_149_clk_i_regs (.I(clknet_6_47__leaf_clk_i_regs),
    .Z(clknet_leaf_149_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16775_ (.I0(net3653),
    .I1(\cs_registers_i.pc_id_i[1] ),
    .S(_08662_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16776_ (.A1(_02398_),
    .A2(_02448_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16777_ (.A1(\cs_registers_i.csr_depc_o[1] ),
    .A2(_02410_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16778_ (.A1(_09468_),
    .A2(_02408_),
    .B(_02449_),
    .C(_02450_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3129 (.I(_03454_),
    .Z(net3129));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16780_ (.I0(\cs_registers_i.pc_if_i[20] ),
    .I1(\cs_registers_i.pc_id_i[20] ),
    .S(net3291),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16781_ (.A1(net3290),
    .A2(_02452_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16782_ (.A1(\cs_registers_i.csr_depc_o[20] ),
    .A2(_02410_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16783_ (.A1(_09262_),
    .A2(_02408_),
    .B(_02453_),
    .C(_02454_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16784_ (.I0(\cs_registers_i.pc_if_i[21] ),
    .I1(\cs_registers_i.pc_id_i[21] ),
    .S(net3291),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16785_ (.A1(net3290),
    .A2(_02455_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16786_ (.A1(\cs_registers_i.csr_depc_o[21] ),
    .A2(_02410_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16787_ (.A1(_09277_),
    .A2(_02408_),
    .B(_02456_),
    .C(_02457_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16788_ (.I0(\cs_registers_i.pc_if_i[22] ),
    .I1(\cs_registers_i.pc_id_i[22] ),
    .S(net3291),
    .Z(_02458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16789_ (.A1(net3290),
    .A2(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16790_ (.A1(\cs_registers_i.csr_depc_o[22] ),
    .A2(_02410_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16791_ (.A1(_09293_),
    .A2(_02408_),
    .B(_02459_),
    .C(_02460_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16792_ (.I0(\cs_registers_i.pc_if_i[23] ),
    .I1(\cs_registers_i.pc_id_i[23] ),
    .S(net3291),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16793_ (.A1(net3290),
    .A2(_02461_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16794_ (.A1(\cs_registers_i.csr_depc_o[23] ),
    .A2(_02410_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16795_ (.A1(_09310_),
    .A2(_02408_),
    .B(_02462_),
    .C(_02463_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16796_ (.I0(\cs_registers_i.pc_if_i[24] ),
    .I1(\cs_registers_i.pc_id_i[24] ),
    .S(net3291),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16797_ (.A1(net3290),
    .A2(_02464_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16798_ (.A1(\cs_registers_i.csr_depc_o[24] ),
    .A2(_02410_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16799_ (.A1(_09330_),
    .A2(_02408_),
    .B(_02465_),
    .C(_02466_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3127 (.I(_03746_),
    .Z(net3127));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16801_ (.I0(\cs_registers_i.pc_if_i[25] ),
    .I1(\cs_registers_i.pc_id_i[25] ),
    .S(net3291),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16802_ (.A1(net3290),
    .A2(_02468_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16803_ (.A1(\cs_registers_i.csr_depc_o[25] ),
    .A2(_02410_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16804_ (.A1(_09348_),
    .A2(_02408_),
    .B(_02469_),
    .C(_02470_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16805_ (.I0(\cs_registers_i.pc_if_i[26] ),
    .I1(\cs_registers_i.pc_id_i[26] ),
    .S(net3291),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16806_ (.A1(net3290),
    .A2(_02471_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16807_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(_02410_),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16808_ (.A1(_09367_),
    .A2(_02408_),
    .B(_02472_),
    .C(_02473_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16809_ (.I0(\cs_registers_i.pc_if_i[27] ),
    .I1(\cs_registers_i.pc_id_i[27] ),
    .S(net3291),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16810_ (.A1(net3290),
    .A2(_02474_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16811_ (.A1(\cs_registers_i.csr_depc_o[27] ),
    .A2(_02410_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16812_ (.A1(_09384_),
    .A2(_02408_),
    .B(_02475_),
    .C(_02476_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16813_ (.I0(\cs_registers_i.pc_if_i[28] ),
    .I1(\cs_registers_i.pc_id_i[28] ),
    .S(net3291),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16814_ (.A1(net3290),
    .A2(_02477_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3642 (.I(net333),
    .Z(net3642));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16816_ (.A1(\cs_registers_i.csr_depc_o[28] ),
    .A2(_02410_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16817_ (.A1(_09401_),
    .A2(_02408_),
    .B(_02478_),
    .C(_02480_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3126 (.I(_09859_[0]),
    .Z(net3126));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16819_ (.I0(\cs_registers_i.pc_if_i[29] ),
    .I1(\cs_registers_i.pc_id_i[29] ),
    .S(net3291),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16820_ (.A1(net3290),
    .A2(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16821_ (.A1(\cs_registers_i.csr_depc_o[29] ),
    .A2(_02410_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16822_ (.A1(_09419_),
    .A2(_02408_),
    .B(_02483_),
    .C(_02484_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16823_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(_02410_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16824_ (.I0(\cs_registers_i.pc_if_i[2] ),
    .I1(\cs_registers_i.pc_id_i[2] ),
    .S(_08662_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16825_ (.A1(_02398_),
    .A2(_02486_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16826_ (.A1(_09423_),
    .A2(_02408_),
    .B(_02485_),
    .C(_02487_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16827_ (.I0(\cs_registers_i.pc_if_i[30] ),
    .I1(\cs_registers_i.pc_id_i[30] ),
    .S(net3291),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16828_ (.A1(net3290),
    .A2(_02488_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16829_ (.A1(\cs_registers_i.csr_depc_o[30] ),
    .A2(_02410_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16830_ (.A1(_09442_),
    .A2(_02408_),
    .B(_02489_),
    .C(_02490_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16831_ (.I0(\cs_registers_i.pc_if_i[31] ),
    .I1(\cs_registers_i.pc_id_i[31] ),
    .S(net3291),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16832_ (.A1(_02398_),
    .A2(_02491_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16833_ (.A1(\cs_registers_i.csr_depc_o[31] ),
    .A2(_02410_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16834_ (.A1(_09458_),
    .A2(_02408_),
    .B(_02492_),
    .C(_02493_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16835_ (.I0(\cs_registers_i.pc_if_i[3] ),
    .I1(\cs_registers_i.pc_id_i[3] ),
    .S(_08662_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16836_ (.A1(_02398_),
    .A2(_02494_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16837_ (.A1(\cs_registers_i.csr_depc_o[3] ),
    .A2(_02410_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16838_ (.A1(_09491_),
    .A2(_02408_),
    .B(_02495_),
    .C(_02496_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16839_ (.I0(\cs_registers_i.pc_if_i[4] ),
    .I1(\cs_registers_i.pc_id_i[4] ),
    .S(_08662_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16840_ (.A1(_02398_),
    .A2(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16841_ (.A1(\cs_registers_i.csr_depc_o[4] ),
    .A2(_02410_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16842_ (.A1(_09508_),
    .A2(_02408_),
    .B(_02498_),
    .C(_02499_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16843_ (.I0(\cs_registers_i.pc_if_i[5] ),
    .I1(\cs_registers_i.pc_id_i[5] ),
    .S(_08662_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16844_ (.A1(_02398_),
    .A2(_02500_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16845_ (.A1(\cs_registers_i.csr_depc_o[5] ),
    .A2(_02410_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16846_ (.A1(_09524_),
    .A2(_02408_),
    .B(_02501_),
    .C(_02502_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16847_ (.I0(\cs_registers_i.pc_if_i[6] ),
    .I1(\cs_registers_i.pc_id_i[6] ),
    .S(_08662_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16848_ (.A1(_02398_),
    .A2(_02503_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16849_ (.A1(\cs_registers_i.csr_depc_o[6] ),
    .A2(_02410_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16850_ (.A1(_09541_),
    .A2(_02408_),
    .B(_02504_),
    .C(_02505_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16851_ (.I0(\cs_registers_i.pc_if_i[7] ),
    .I1(\cs_registers_i.pc_id_i[7] ),
    .S(_08662_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16852_ (.A1(_02398_),
    .A2(_02506_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16853_ (.A1(\cs_registers_i.csr_depc_o[7] ),
    .A2(_02410_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16854_ (.A1(_09593_),
    .A2(_02408_),
    .B(_02507_),
    .C(_02508_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16855_ (.I0(\cs_registers_i.pc_if_i[8] ),
    .I1(\cs_registers_i.pc_id_i[8] ),
    .S(net3291),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16856_ (.A1(_02398_),
    .A2(_02509_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16857_ (.A1(\cs_registers_i.csr_depc_o[8] ),
    .A2(_02410_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16858_ (.A1(_09613_),
    .A2(_02408_),
    .B(_02510_),
    .C(_02511_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16859_ (.I0(\cs_registers_i.pc_if_i[9] ),
    .I1(\cs_registers_i.pc_id_i[9] ),
    .S(net3291),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16860_ (.A1(net3290),
    .A2(_02512_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16861_ (.A1(\cs_registers_i.csr_depc_o[9] ),
    .A2(_02410_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16862_ (.A1(_09628_),
    .A2(_02408_),
    .B(_02513_),
    .C(_02514_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16863_ (.A1(_08946_),
    .A2(_08951_),
    .A3(net3199),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3131 (.I(_11355_[0]),
    .Z(net3131));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16865_ (.I0(_08945_),
    .I1(\cs_registers_i.dscratch0_q[0] ),
    .S(_02515_),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16866_ (.I0(_09028_),
    .I1(\cs_registers_i.dscratch0_q[10] ),
    .S(_02515_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16867_ (.I0(_02217_),
    .I1(\cs_registers_i.dscratch0_q[11] ),
    .S(_02515_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16868_ (.I0(_02221_),
    .I1(\cs_registers_i.dscratch0_q[12] ),
    .S(net3193),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16869_ (.I0(_02025_),
    .I1(\cs_registers_i.dscratch0_q[13] ),
    .S(net3193),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16870_ (.I0(_09132_),
    .I1(\cs_registers_i.dscratch0_q[14] ),
    .S(net3193),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16871_ (.I0(_02038_),
    .I1(\cs_registers_i.dscratch0_q[15] ),
    .S(_02515_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16872_ (.I0(_02250_),
    .I1(\cs_registers_i.dscratch0_q[16] ),
    .S(net3193),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16873_ (.I(_09194_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3123 (.I(_11273_[0]),
    .Z(net3123));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16875_ (.I0(_02517_),
    .I1(\cs_registers_i.dscratch0_q[17] ),
    .S(net3193),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16876_ (.I0(_02271_),
    .I1(\cs_registers_i.dscratch0_q[18] ),
    .S(_02515_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16877_ (.I0(_02277_),
    .I1(\cs_registers_i.dscratch0_q[19] ),
    .S(net3193),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16878_ (.I0(_09245_),
    .I1(\cs_registers_i.dscratch0_q[1] ),
    .S(_02515_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16879_ (.I0(_02282_),
    .I1(\cs_registers_i.dscratch0_q[20] ),
    .S(_02515_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16880_ (.I(_09277_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16881_ (.I0(_02519_),
    .I1(\cs_registers_i.dscratch0_q[21] ),
    .S(net3193),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16882_ (.I(_09293_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16883_ (.I0(_02520_),
    .I1(\cs_registers_i.dscratch0_q[22] ),
    .S(net3193),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16884_ (.I(_09310_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16885_ (.I0(_02521_),
    .I1(\cs_registers_i.dscratch0_q[23] ),
    .S(net3193),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16886_ (.I0(_02306_),
    .I1(\cs_registers_i.dscratch0_q[24] ),
    .S(_02515_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16887_ (.I0(_02099_),
    .I1(\cs_registers_i.dscratch0_q[25] ),
    .S(_02515_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3561 (.I(net3558),
    .Z(net3561));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16889_ (.I0(_02321_),
    .I1(\cs_registers_i.dscratch0_q[26] ),
    .S(_02515_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16890_ (.I0(_02330_),
    .I1(\cs_registers_i.dscratch0_q[27] ),
    .S(_02515_),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16891_ (.I0(_02338_),
    .I1(\cs_registers_i.dscratch0_q[28] ),
    .S(_02515_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16892_ (.I0(_02344_),
    .I1(\cs_registers_i.dscratch0_q[29] ),
    .S(_02515_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16893_ (.I0(_08984_),
    .I1(\cs_registers_i.dscratch0_q[2] ),
    .S(_02515_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16894_ (.I0(_02134_),
    .I1(\cs_registers_i.dscratch0_q[30] ),
    .S(net3193),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16895_ (.I0(_09457_),
    .I1(\cs_registers_i.dscratch0_q[31] ),
    .S(_02515_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16896_ (.A1(\cs_registers_i.dscratch0_q[3] ),
    .A2(_02515_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16897_ (.A1(_09491_),
    .A2(_02515_),
    .B(_02523_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16898_ (.I0(_09663_),
    .I1(\cs_registers_i.dscratch0_q[4] ),
    .S(_02515_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16899_ (.I(_09524_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16900_ (.I0(_02524_),
    .I1(\cs_registers_i.dscratch0_q[5] ),
    .S(_02515_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16901_ (.I(_09541_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16902_ (.I0(_02525_),
    .I1(\cs_registers_i.dscratch0_q[6] ),
    .S(_02515_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16903_ (.I(_09593_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16904_ (.I0(_02526_),
    .I1(\cs_registers_i.dscratch0_q[7] ),
    .S(_02515_),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16905_ (.I(_09613_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16906_ (.I0(_02527_),
    .I1(\cs_registers_i.dscratch0_q[8] ),
    .S(_02515_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16907_ (.I(_09628_),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16908_ (.I0(_02528_),
    .I1(\cs_registers_i.dscratch0_q[9] ),
    .S(net3193),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16909_ (.A1(_08946_),
    .A2(_08951_),
    .A3(_08940_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3125 (.I(_11272_[0]),
    .Z(net3125));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16911_ (.I0(_08945_),
    .I1(\cs_registers_i.dscratch1_q[0] ),
    .S(_02529_),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16912_ (.I0(_09028_),
    .I1(\cs_registers_i.dscratch1_q[10] ),
    .S(_02529_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16913_ (.I0(_02217_),
    .I1(\cs_registers_i.dscratch1_q[11] ),
    .S(_02529_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16914_ (.I0(_02221_),
    .I1(\cs_registers_i.dscratch1_q[12] ),
    .S(_02529_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16915_ (.I0(_02025_),
    .I1(\cs_registers_i.dscratch1_q[13] ),
    .S(_02529_),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16916_ (.I0(_09132_),
    .I1(\cs_registers_i.dscratch1_q[14] ),
    .S(net3192),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16917_ (.I0(_02038_),
    .I1(\cs_registers_i.dscratch1_q[15] ),
    .S(net3192),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16918_ (.I0(_02250_),
    .I1(\cs_registers_i.dscratch1_q[16] ),
    .S(net3192),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16919_ (.I0(_02517_),
    .I1(\cs_registers_i.dscratch1_q[17] ),
    .S(net3192),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16920_ (.I0(_02271_),
    .I1(\cs_registers_i.dscratch1_q[18] ),
    .S(net3192),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3121 (.I(net3120),
    .Z(net3121));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16922_ (.I0(_02277_),
    .I1(\cs_registers_i.dscratch1_q[19] ),
    .S(net3192),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16923_ (.I0(_09245_),
    .I1(\cs_registers_i.dscratch1_q[1] ),
    .S(_02529_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16924_ (.I0(_02282_),
    .I1(\cs_registers_i.dscratch1_q[20] ),
    .S(net3192),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16925_ (.I0(_02519_),
    .I1(\cs_registers_i.dscratch1_q[21] ),
    .S(net3192),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16926_ (.I0(_02520_),
    .I1(\cs_registers_i.dscratch1_q[22] ),
    .S(net3192),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16927_ (.I0(_02521_),
    .I1(\cs_registers_i.dscratch1_q[23] ),
    .S(net3192),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16928_ (.I0(_02306_),
    .I1(\cs_registers_i.dscratch1_q[24] ),
    .S(net3192),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16929_ (.I0(_02099_),
    .I1(\cs_registers_i.dscratch1_q[25] ),
    .S(net3192),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16930_ (.I0(_02321_),
    .I1(\cs_registers_i.dscratch1_q[26] ),
    .S(net3192),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16931_ (.I0(_02330_),
    .I1(\cs_registers_i.dscratch1_q[27] ),
    .S(net3192),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 place3117 (.I(_11288_[0]),
    .Z(net3117));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16933_ (.I0(_02338_),
    .I1(\cs_registers_i.dscratch1_q[28] ),
    .S(net3192),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16934_ (.I0(_02344_),
    .I1(\cs_registers_i.dscratch1_q[29] ),
    .S(net3192),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16935_ (.I0(_08984_),
    .I1(\cs_registers_i.dscratch1_q[2] ),
    .S(_02529_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16936_ (.I0(_02134_),
    .I1(\cs_registers_i.dscratch1_q[30] ),
    .S(net3192),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16937_ (.I0(_09457_),
    .I1(\cs_registers_i.dscratch1_q[31] ),
    .S(_02529_),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16938_ (.I(\cs_registers_i.dscratch1_q[3] ),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16939_ (.I0(_09491_),
    .I1(_02533_),
    .S(_02529_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16940_ (.I(_02534_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16941_ (.I0(_09663_),
    .I1(\cs_registers_i.dscratch1_q[4] ),
    .S(_02529_),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16942_ (.I0(_02524_),
    .I1(\cs_registers_i.dscratch1_q[5] ),
    .S(_02529_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16943_ (.I0(_02525_),
    .I1(\cs_registers_i.dscratch1_q[6] ),
    .S(_02529_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16944_ (.I0(_02526_),
    .I1(\cs_registers_i.dscratch1_q[7] ),
    .S(_02529_),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16945_ (.I0(_02527_),
    .I1(\cs_registers_i.dscratch1_q[8] ),
    .S(_02529_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16946_ (.I0(_02528_),
    .I1(\cs_registers_i.dscratch1_q[9] ),
    .S(net3192),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _16947_ (.A1(_08370_),
    .A2(_02385_),
    .A3(_02399_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3118 (.I(_11288_[0]),
    .Z(net3118));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _16949_ (.A1(\cs_registers_i.nmi_mode_i ),
    .A2(_08709_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16950_ (.A1(_02535_),
    .A2(_02537_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3116 (.I(_11289_[0]),
    .Z(net3116));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3119 (.I(_11287_[0]),
    .Z(net3119));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16953_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.load_err_q ),
    .A3(_08393_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16954_ (.A1(net3560),
    .A2(_08381_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16955_ (.A1(net3560),
    .A2(_08633_),
    .B(_02542_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16956_ (.I(_02543_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16957_ (.A1(_08393_),
    .A2(_02544_),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16958_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_02541_),
    .A3(_02545_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16959_ (.A1(_08626_),
    .A2(_02546_),
    .B(_08629_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16960_ (.A1(_08707_),
    .A2(_02547_),
    .Z(_02548_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3114 (.I(_11294_[0]),
    .Z(net3114));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16962_ (.A1(\cs_registers_i.mstack_cause_q[0] ),
    .A2(_02537_),
    .B1(_02548_),
    .B2(_02535_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16963_ (.A1(_08985_),
    .A2(_02538_),
    .B(_02550_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16964_ (.I(_08898_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16965_ (.A1(_02535_),
    .A2(_02537_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _16966_ (.A1(_02143_),
    .A2(_02552_),
    .B(_02553_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16967_ (.I0(\cs_registers_i.mcause_q[0] ),
    .I1(_02551_),
    .S(_02554_),
    .Z(_00251_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place3115 (.I(_11290_[0]),
    .Z(net3115));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16969_ (.I0(\id_stage_i.controller_i.store_err_q ),
    .I1(_02543_),
    .S(_08393_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16970_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_02556_),
    .B(_08724_),
    .C(_08626_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _16971_ (.A1(_08370_),
    .A2(_02385_),
    .A3(_02399_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16972_ (.A1(_08723_),
    .A2(_02557_),
    .B(_02558_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16973_ (.A1(\cs_registers_i.mstack_cause_q[1] ),
    .A2(_02537_),
    .B1(_02553_),
    .B2(_09245_),
    .C(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16974_ (.I(_02560_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16975_ (.I0(\cs_registers_i.mcause_q[1] ),
    .I1(_02561_),
    .S(_02554_),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_151_clk_i_regs (.I(clknet_6_45__leaf_clk_i_regs),
    .Z(clknet_leaf_151_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16977_ (.A1(_09423_),
    .A2(_02538_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16978_ (.A1(net3382),
    .A2(_08655_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16979_ (.A1(net3406),
    .A2(net3405),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16980_ (.A1(_02565_),
    .A2(net3402),
    .A3(net3401),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16981_ (.A1(net3403),
    .A2(_02564_),
    .A3(_08720_),
    .A4(_02566_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16982_ (.A1(_08706_),
    .A2(_02567_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16983_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.load_err_q ),
    .B(_08635_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16984_ (.A1(_08393_),
    .A2(_02569_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16985_ (.A1(_08391_),
    .A2(_02570_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16986_ (.A1(_02568_),
    .A2(_02571_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_154_clk_i_regs (.I(clknet_6_45__leaf_clk_i_regs),
    .Z(clknet_leaf_154_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16988_ (.A1(\cs_registers_i.mstack_cause_q[2] ),
    .A2(_02537_),
    .B1(_02572_),
    .B2(_02535_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16989_ (.A1(_02563_),
    .A2(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16990_ (.I0(\cs_registers_i.mcause_q[2] ),
    .I1(_02575_),
    .S(_02554_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _16991_ (.A1(_09491_),
    .A2(_02538_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16992_ (.A1(net129),
    .A2(\cs_registers_i.mie_q[15] ),
    .A3(_08648_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16993_ (.A1(_08652_),
    .A2(_08720_),
    .A3(_02577_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _16994_ (.A1(_08706_),
    .A2(_02578_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16995_ (.A1(net3449),
    .A2(_08393_),
    .A3(_08724_),
    .A4(_08635_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16996_ (.A1(_02579_),
    .A2(_02580_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3113 (.I(_11295_[0]),
    .Z(net3113));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16998_ (.A1(\cs_registers_i.mstack_cause_q[3] ),
    .A2(_02537_),
    .B1(_02581_),
    .B2(_02535_),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16999_ (.A1(_02576_),
    .A2(_02583_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17000_ (.I0(\cs_registers_i.mcause_q[3] ),
    .I1(_02584_),
    .S(_02554_),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17001_ (.A1(_09508_),
    .A2(_02538_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17002_ (.A1(net3382),
    .A2(_08719_),
    .B(_08641_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17003_ (.A1(\cs_registers_i.mstack_cause_q[4] ),
    .A2(_02537_),
    .B(_02586_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17004_ (.A1(_02585_),
    .A2(_02587_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17005_ (.I0(\cs_registers_i.mcause_q[4] ),
    .I1(_02588_),
    .S(_02554_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17006_ (.A1(_09457_),
    .A2(_02553_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17007_ (.A1(\cs_registers_i.mstack_cause_q[5] ),
    .A2(_02537_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17008_ (.A1(_08706_),
    .A2(_02589_),
    .A3(_02590_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17009_ (.I0(\cs_registers_i.mcause_q[5] ),
    .I1(_02591_),
    .S(_02554_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17010_ (.I(_08932_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17011_ (.A1(_02143_),
    .A2(_02592_),
    .B(_02553_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3566 (.I(net3558),
    .Z(net3566));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17013_ (.I(_02593_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17014_ (.A1(\cs_registers_i.mstack_epc_q[0] ),
    .A2(_02537_),
    .B1(_02595_),
    .B2(\cs_registers_i.csr_mepc_o[0] ),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17015_ (.I(_02596_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17016_ (.A1(_02415_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[10] ),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17017_ (.A1(_09029_),
    .A2(_02538_),
    .B(_02597_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17018_ (.I0(\cs_registers_i.csr_mepc_o[10] ),
    .I1(_02598_),
    .S(net3189),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17019_ (.A1(_02418_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[11] ),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17020_ (.A1(_09066_),
    .A2(_02538_),
    .B(_02599_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17021_ (.I0(\cs_registers_i.csr_mepc_o[11] ),
    .I1(_02600_),
    .S(net3189),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17022_ (.A1(_02421_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[12] ),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17023_ (.A1(_09096_),
    .A2(_02538_),
    .B(_02601_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17024_ (.I0(\cs_registers_i.csr_mepc_o[12] ),
    .I1(_02602_),
    .S(net3189),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17025_ (.A1(_02424_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[13] ),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17026_ (.A1(_09117_),
    .A2(_02538_),
    .B(_02603_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17027_ (.I0(\cs_registers_i.csr_mepc_o[13] ),
    .I1(_02604_),
    .S(net3189),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17028_ (.A1(_02427_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[14] ),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17029_ (.A1(_09133_),
    .A2(_02538_),
    .B(_02605_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17030_ (.I0(\cs_registers_i.csr_mepc_o[14] ),
    .I1(_02606_),
    .S(net3189),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17031_ (.A1(_02430_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[15] ),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17032_ (.A1(_09149_),
    .A2(_02538_),
    .B(_02607_),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17033_ (.I0(\cs_registers_i.csr_mepc_o[15] ),
    .I1(_02608_),
    .S(net3189),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17034_ (.A1(_02434_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[16] ),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17035_ (.A1(_09174_),
    .A2(_02538_),
    .B(_02609_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17036_ (.I0(\cs_registers_i.csr_mepc_o[16] ),
    .I1(_02610_),
    .S(net3189),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3641 (.I(net3634),
    .Z(net3641));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17038_ (.A1(_02437_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[17] ),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17039_ (.A1(_09194_),
    .A2(_02538_),
    .B(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17040_ (.I0(\cs_registers_i.csr_mepc_o[17] ),
    .I1(_02613_),
    .S(net3189),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17041_ (.A1(_02440_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[18] ),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17042_ (.A1(_09210_),
    .A2(_02538_),
    .B(_02614_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17043_ (.I0(\cs_registers_i.csr_mepc_o[18] ),
    .I1(_02615_),
    .S(net3189),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3109 (.I(_03513_),
    .Z(net3109));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3640 (.I(net3634),
    .Z(net3640));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17046_ (.A1(_02443_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[19] ),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17047_ (.A1(_09229_),
    .A2(_02538_),
    .B(_02618_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3108 (.I(_03515_),
    .Z(net3108));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17049_ (.I0(\cs_registers_i.csr_mepc_o[19] ),
    .I1(_02619_),
    .S(net3189),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17050_ (.A1(_02448_),
    .A2(_02535_),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[1] ),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17051_ (.A1(_09468_),
    .A2(_02538_),
    .B(_02621_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17052_ (.I0(\cs_registers_i.csr_mepc_o[1] ),
    .I1(_02622_),
    .S(_02593_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17053_ (.A1(_02452_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[20] ),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17054_ (.A1(_09262_),
    .A2(_02538_),
    .B(_02623_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17055_ (.I0(\cs_registers_i.csr_mepc_o[20] ),
    .I1(_02624_),
    .S(net3189),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17056_ (.A1(_02455_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[21] ),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17057_ (.A1(_09277_),
    .A2(_02538_),
    .B(_02625_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17058_ (.I0(\cs_registers_i.csr_mepc_o[21] ),
    .I1(_02626_),
    .S(net3189),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17059_ (.A1(_02458_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[22] ),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17060_ (.A1(_09293_),
    .A2(_02538_),
    .B(_02627_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17061_ (.I0(\cs_registers_i.csr_mepc_o[22] ),
    .I1(_02628_),
    .S(net3189),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17062_ (.A1(_02461_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[23] ),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17063_ (.A1(_09310_),
    .A2(_02538_),
    .B(_02629_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17064_ (.I0(\cs_registers_i.csr_mepc_o[23] ),
    .I1(_02630_),
    .S(net3189),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17065_ (.A1(_02464_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[24] ),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17066_ (.A1(_09330_),
    .A2(_02538_),
    .B(_02631_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17067_ (.I0(\cs_registers_i.csr_mepc_o[24] ),
    .I1(_02632_),
    .S(net3189),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17068_ (.A1(_02468_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[25] ),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17069_ (.A1(_09348_),
    .A2(_02538_),
    .B(_02633_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17070_ (.I0(\cs_registers_i.csr_mepc_o[25] ),
    .I1(_02634_),
    .S(net3189),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3565 (.I(net3558),
    .Z(net3565));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17072_ (.A1(_02471_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[26] ),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17073_ (.A1(_09367_),
    .A2(_02538_),
    .B(_02636_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17074_ (.I0(\cs_registers_i.csr_mepc_o[26] ),
    .I1(_02637_),
    .S(net3189),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17075_ (.A1(_02474_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[27] ),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17076_ (.A1(_09384_),
    .A2(_02538_),
    .B(_02638_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17077_ (.I0(\cs_registers_i.csr_mepc_o[27] ),
    .I1(_02639_),
    .S(net3189),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17078_ (.A1(_02477_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[28] ),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17079_ (.A1(_09401_),
    .A2(_02538_),
    .B(_02640_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_156_clk_i_regs (.I(clknet_6_44__leaf_clk_i_regs),
    .Z(clknet_leaf_156_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17081_ (.I0(\cs_registers_i.csr_mepc_o[28] ),
    .I1(_02641_),
    .S(net3189),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17082_ (.A1(_02482_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[29] ),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17083_ (.A1(_09419_),
    .A2(_02538_),
    .B(_02643_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17084_ (.I0(\cs_registers_i.csr_mepc_o[29] ),
    .I1(_02644_),
    .S(net3189),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17085_ (.A1(_02486_),
    .A2(_02535_),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[2] ),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17086_ (.A1(_02563_),
    .A2(_02645_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17087_ (.I0(\cs_registers_i.csr_mepc_o[2] ),
    .I1(_02646_),
    .S(_02593_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17088_ (.A1(_02488_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[30] ),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17089_ (.A1(_09442_),
    .A2(_02538_),
    .B(_02647_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17090_ (.I0(\cs_registers_i.csr_mepc_o[30] ),
    .I1(_02648_),
    .S(net3189),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17091_ (.A1(_02491_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[31] ),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17092_ (.A1(_02589_),
    .A2(_02649_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17093_ (.I0(\cs_registers_i.csr_mepc_o[31] ),
    .I1(_02650_),
    .S(net3189),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17094_ (.A1(_02494_),
    .A2(_02535_),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[3] ),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17095_ (.A1(_02576_),
    .A2(_02651_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17096_ (.I0(\cs_registers_i.csr_mepc_o[3] ),
    .I1(_02652_),
    .S(_02593_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17097_ (.A1(_02497_),
    .A2(_02535_),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[4] ),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17098_ (.A1(_02585_),
    .A2(_02653_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17099_ (.I0(\cs_registers_i.csr_mepc_o[4] ),
    .I1(_02654_),
    .S(_02593_),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17100_ (.A1(_02500_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[5] ),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17101_ (.A1(_09524_),
    .A2(_02538_),
    .B(_02655_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17102_ (.I0(\cs_registers_i.csr_mepc_o[5] ),
    .I1(_02656_),
    .S(net3189),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17103_ (.A1(_02503_),
    .A2(_02535_),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[6] ),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17104_ (.A1(_09541_),
    .A2(_02538_),
    .B(_02657_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17105_ (.I0(\cs_registers_i.csr_mepc_o[6] ),
    .I1(_02658_),
    .S(net3189),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17106_ (.A1(_02506_),
    .A2(_02535_),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[7] ),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17107_ (.A1(_09593_),
    .A2(_02538_),
    .B(_02659_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17108_ (.I0(\cs_registers_i.csr_mepc_o[7] ),
    .I1(_02660_),
    .S(net3189),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17109_ (.A1(_02509_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[8] ),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17110_ (.A1(_09613_),
    .A2(_02538_),
    .B(_02661_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17111_ (.I0(\cs_registers_i.csr_mepc_o[8] ),
    .I1(_02662_),
    .S(net3189),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17112_ (.A1(_02512_),
    .A2(net3220),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_epc_q[9] ),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17113_ (.A1(_09628_),
    .A2(_02538_),
    .B(_02663_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17114_ (.I0(\cs_registers_i.csr_mepc_o[9] ),
    .I1(_02664_),
    .S(net3189),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17115_ (.A1(_08946_),
    .A2(_08951_),
    .A3(_09043_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_158_clk_i_regs (.I(clknet_6_44__leaf_clk_i_regs),
    .Z(clknet_leaf_158_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17117_ (.I0(_02250_),
    .I1(\cs_registers_i.mie_q[0] ),
    .S(_02665_),
    .Z(_00289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17118_ (.I0(_02321_),
    .I1(\cs_registers_i.mie_q[10] ),
    .S(_02665_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17119_ (.I0(_02330_),
    .I1(\cs_registers_i.mie_q[11] ),
    .S(_02665_),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17120_ (.I0(_02338_),
    .I1(\cs_registers_i.mie_q[12] ),
    .S(_02665_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17121_ (.I0(_02344_),
    .I1(\cs_registers_i.mie_q[13] ),
    .S(_02665_),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17122_ (.I0(_02134_),
    .I1(\cs_registers_i.mie_q[14] ),
    .S(_02665_),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17123_ (.I0(_02217_),
    .I1(\cs_registers_i.mie_q[15] ),
    .S(_02665_),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17124_ (.I0(_02526_),
    .I1(\cs_registers_i.mie_q[16] ),
    .S(_02665_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17125_ (.I(\cs_registers_i.mie_q[17] ),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17126_ (.I0(_09491_),
    .I1(_02667_),
    .S(_02665_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17127_ (.I(_02668_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17128_ (.I0(_02517_),
    .I1(\cs_registers_i.mie_q[1] ),
    .S(_02665_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17129_ (.I0(_02271_),
    .I1(\cs_registers_i.mie_q[2] ),
    .S(_02665_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17130_ (.I0(_02277_),
    .I1(\cs_registers_i.mie_q[3] ),
    .S(_02665_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17131_ (.I0(_02282_),
    .I1(\cs_registers_i.mie_q[4] ),
    .S(_02665_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17132_ (.I0(_02519_),
    .I1(\cs_registers_i.mie_q[5] ),
    .S(_02665_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17133_ (.I0(_02520_),
    .I1(\cs_registers_i.mie_q[6] ),
    .S(_02665_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17134_ (.I0(_02521_),
    .I1(\cs_registers_i.mie_q[7] ),
    .S(_02665_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17135_ (.I0(_02306_),
    .I1(\cs_registers_i.mie_q[8] ),
    .S(_02665_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17136_ (.I0(_02099_),
    .I1(\cs_registers_i.mie_q[9] ),
    .S(_02665_),
    .Z(_00306_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17137_ (.A1(_08946_),
    .A2(_08951_),
    .A3(_08899_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3107 (.I(_03658_),
    .Z(net3107));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17139_ (.I0(_08945_),
    .I1(\cs_registers_i.mscratch_q[0] ),
    .S(_02669_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17140_ (.I0(_09028_),
    .I1(\cs_registers_i.mscratch_q[10] ),
    .S(_02669_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17141_ (.I0(_02217_),
    .I1(\cs_registers_i.mscratch_q[11] ),
    .S(_02669_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17142_ (.I0(_02221_),
    .I1(\cs_registers_i.mscratch_q[12] ),
    .S(_02669_),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17143_ (.I0(_02025_),
    .I1(\cs_registers_i.mscratch_q[13] ),
    .S(_02669_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17144_ (.I0(_09132_),
    .I1(\cs_registers_i.mscratch_q[14] ),
    .S(net3191),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17145_ (.I0(_02038_),
    .I1(\cs_registers_i.mscratch_q[15] ),
    .S(_02669_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17146_ (.I0(_02250_),
    .I1(\cs_registers_i.mscratch_q[16] ),
    .S(net3191),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_162_clk_i_regs (.I(clknet_6_35__leaf_clk_i_regs),
    .Z(clknet_leaf_162_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17148_ (.I0(_02517_),
    .I1(\cs_registers_i.mscratch_q[17] ),
    .S(net3191),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17149_ (.I0(_02271_),
    .I1(\cs_registers_i.mscratch_q[18] ),
    .S(net3191),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17150_ (.I0(_02277_),
    .I1(\cs_registers_i.mscratch_q[19] ),
    .S(net3191),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17151_ (.I0(_09245_),
    .I1(\cs_registers_i.mscratch_q[1] ),
    .S(_02669_),
    .Z(_00318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17152_ (.I0(_02282_),
    .I1(\cs_registers_i.mscratch_q[20] ),
    .S(net3191),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17153_ (.I0(_02519_),
    .I1(\cs_registers_i.mscratch_q[21] ),
    .S(net3191),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17154_ (.I0(_02520_),
    .I1(\cs_registers_i.mscratch_q[22] ),
    .S(net3191),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17155_ (.I0(_02521_),
    .I1(\cs_registers_i.mscratch_q[23] ),
    .S(net3191),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17156_ (.I0(_02306_),
    .I1(\cs_registers_i.mscratch_q[24] ),
    .S(net3191),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17157_ (.I0(_02099_),
    .I1(\cs_registers_i.mscratch_q[25] ),
    .S(net3191),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_160_clk_i_regs (.I(clknet_6_35__leaf_clk_i_regs),
    .Z(clknet_leaf_160_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17159_ (.I0(_02321_),
    .I1(\cs_registers_i.mscratch_q[26] ),
    .S(net3191),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17160_ (.I0(_02330_),
    .I1(\cs_registers_i.mscratch_q[27] ),
    .S(net3191),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17161_ (.I0(_02338_),
    .I1(\cs_registers_i.mscratch_q[28] ),
    .S(net3191),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17162_ (.I0(_02344_),
    .I1(\cs_registers_i.mscratch_q[29] ),
    .S(net3191),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17163_ (.I0(_08984_),
    .I1(\cs_registers_i.mscratch_q[2] ),
    .S(_02669_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17164_ (.I0(_02134_),
    .I1(\cs_registers_i.mscratch_q[30] ),
    .S(net3191),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17165_ (.I0(_09457_),
    .I1(\cs_registers_i.mscratch_q[31] ),
    .S(_02669_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17166_ (.A1(\cs_registers_i.mscratch_q[3] ),
    .A2(_02669_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17167_ (.A1(_09491_),
    .A2(_02669_),
    .B(_02673_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17168_ (.I0(_09663_),
    .I1(\cs_registers_i.mscratch_q[4] ),
    .S(_02669_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17169_ (.I0(_02524_),
    .I1(\cs_registers_i.mscratch_q[5] ),
    .S(_02669_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17170_ (.I0(_02525_),
    .I1(\cs_registers_i.mscratch_q[6] ),
    .S(_02669_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17171_ (.I0(_02526_),
    .I1(\cs_registers_i.mscratch_q[7] ),
    .S(_02669_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17172_ (.I0(_02527_),
    .I1(\cs_registers_i.mscratch_q[8] ),
    .S(_02669_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17173_ (.I0(_02528_),
    .I1(\cs_registers_i.mscratch_q[9] ),
    .S(net3191),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_165_clk_i_regs (.I(clknet_6_35__leaf_clk_i_regs),
    .Z(clknet_leaf_165_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17175_ (.I0(\cs_registers_i.mcause_q[0] ),
    .I1(\cs_registers_i.mstack_cause_q[0] ),
    .S(_02558_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17176_ (.I0(\cs_registers_i.mcause_q[1] ),
    .I1(\cs_registers_i.mstack_cause_q[1] ),
    .S(_02558_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17177_ (.I0(\cs_registers_i.mcause_q[2] ),
    .I1(\cs_registers_i.mstack_cause_q[2] ),
    .S(_02558_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17178_ (.I0(\cs_registers_i.mcause_q[3] ),
    .I1(\cs_registers_i.mstack_cause_q[3] ),
    .S(_02558_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17179_ (.I0(\cs_registers_i.mcause_q[4] ),
    .I1(\cs_registers_i.mstack_cause_q[4] ),
    .S(_02558_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17180_ (.I0(\cs_registers_i.mcause_q[5] ),
    .I1(\cs_registers_i.mstack_cause_q[5] ),
    .S(_02558_),
    .Z(_00344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17181_ (.I0(\cs_registers_i.mstatus_q[2] ),
    .I1(\cs_registers_i.mstack_q[0] ),
    .S(_02558_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17182_ (.I0(\cs_registers_i.mstatus_q[3] ),
    .I1(\cs_registers_i.mstack_q[1] ),
    .S(_02558_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17183_ (.I0(\cs_registers_i.mstatus_q[4] ),
    .I1(\cs_registers_i.mstack_q[2] ),
    .S(_02558_),
    .Z(_00347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17184_ (.I0(\cs_registers_i.csr_mepc_o[0] ),
    .I1(\cs_registers_i.mstack_epc_q[0] ),
    .S(_02558_),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_166_clk_i_regs (.I(clknet_6_50__leaf_clk_i_regs),
    .Z(clknet_leaf_166_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17186_ (.I0(\cs_registers_i.csr_mepc_o[10] ),
    .I1(\cs_registers_i.mstack_epc_q[10] ),
    .S(net3219),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17187_ (.I0(\cs_registers_i.csr_mepc_o[11] ),
    .I1(\cs_registers_i.mstack_epc_q[11] ),
    .S(_02558_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17188_ (.I0(\cs_registers_i.csr_mepc_o[12] ),
    .I1(\cs_registers_i.mstack_epc_q[12] ),
    .S(_02558_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17189_ (.I0(\cs_registers_i.csr_mepc_o[13] ),
    .I1(\cs_registers_i.mstack_epc_q[13] ),
    .S(net3219),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17190_ (.I0(\cs_registers_i.csr_mepc_o[14] ),
    .I1(\cs_registers_i.mstack_epc_q[14] ),
    .S(net3219),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17191_ (.I0(\cs_registers_i.csr_mepc_o[15] ),
    .I1(\cs_registers_i.mstack_epc_q[15] ),
    .S(_02558_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17192_ (.I0(\cs_registers_i.csr_mepc_o[16] ),
    .I1(\cs_registers_i.mstack_epc_q[16] ),
    .S(net3219),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17193_ (.I0(\cs_registers_i.csr_mepc_o[17] ),
    .I1(\cs_registers_i.mstack_epc_q[17] ),
    .S(net3219),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17194_ (.I0(\cs_registers_i.csr_mepc_o[18] ),
    .I1(\cs_registers_i.mstack_epc_q[18] ),
    .S(net3219),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17195_ (.I0(\cs_registers_i.csr_mepc_o[19] ),
    .I1(\cs_registers_i.mstack_epc_q[19] ),
    .S(net3219),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3106 (.I(_03701_),
    .Z(net3106));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17197_ (.I0(\cs_registers_i.csr_mepc_o[1] ),
    .I1(\cs_registers_i.mstack_epc_q[1] ),
    .S(_02558_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17198_ (.I0(\cs_registers_i.csr_mepc_o[20] ),
    .I1(\cs_registers_i.mstack_epc_q[20] ),
    .S(_02558_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17199_ (.I0(\cs_registers_i.csr_mepc_o[21] ),
    .I1(\cs_registers_i.mstack_epc_q[21] ),
    .S(net3219),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17200_ (.I0(\cs_registers_i.csr_mepc_o[22] ),
    .I1(\cs_registers_i.mstack_epc_q[22] ),
    .S(net3219),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17201_ (.I0(\cs_registers_i.csr_mepc_o[23] ),
    .I1(\cs_registers_i.mstack_epc_q[23] ),
    .S(net3219),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17202_ (.I0(\cs_registers_i.csr_mepc_o[24] ),
    .I1(\cs_registers_i.mstack_epc_q[24] ),
    .S(net3219),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17203_ (.I0(\cs_registers_i.csr_mepc_o[25] ),
    .I1(\cs_registers_i.mstack_epc_q[25] ),
    .S(net3219),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17204_ (.I0(\cs_registers_i.csr_mepc_o[26] ),
    .I1(\cs_registers_i.mstack_epc_q[26] ),
    .S(net3219),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17205_ (.I0(\cs_registers_i.csr_mepc_o[27] ),
    .I1(\cs_registers_i.mstack_epc_q[27] ),
    .S(net3219),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17206_ (.I0(\cs_registers_i.csr_mepc_o[28] ),
    .I1(\cs_registers_i.mstack_epc_q[28] ),
    .S(net3219),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3105 (.I(_03747_),
    .Z(net3105));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17208_ (.I0(\cs_registers_i.csr_mepc_o[29] ),
    .I1(\cs_registers_i.mstack_epc_q[29] ),
    .S(net3219),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17209_ (.I0(\cs_registers_i.csr_mepc_o[2] ),
    .I1(\cs_registers_i.mstack_epc_q[2] ),
    .S(_02558_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17210_ (.I0(\cs_registers_i.csr_mepc_o[30] ),
    .I1(\cs_registers_i.mstack_epc_q[30] ),
    .S(net3219),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17211_ (.I0(\cs_registers_i.csr_mepc_o[31] ),
    .I1(\cs_registers_i.mstack_epc_q[31] ),
    .S(_02558_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17212_ (.I0(\cs_registers_i.csr_mepc_o[3] ),
    .I1(\cs_registers_i.mstack_epc_q[3] ),
    .S(_02558_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17213_ (.I0(\cs_registers_i.csr_mepc_o[4] ),
    .I1(\cs_registers_i.mstack_epc_q[4] ),
    .S(_02558_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17214_ (.I0(\cs_registers_i.csr_mepc_o[5] ),
    .I1(\cs_registers_i.mstack_epc_q[5] ),
    .S(_02558_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17215_ (.I0(\cs_registers_i.csr_mepc_o[6] ),
    .I1(\cs_registers_i.mstack_epc_q[6] ),
    .S(_02558_),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17216_ (.I0(\cs_registers_i.csr_mepc_o[7] ),
    .I1(\cs_registers_i.mstack_epc_q[7] ),
    .S(_02558_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17217_ (.I0(\cs_registers_i.csr_mepc_o[8] ),
    .I1(\cs_registers_i.mstack_epc_q[8] ),
    .S(_02558_),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17218_ (.I0(\cs_registers_i.csr_mepc_o[9] ),
    .I1(\cs_registers_i.mstack_epc_q[9] ),
    .S(net3219),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17219_ (.A1(_08946_),
    .A2(_08951_),
    .A3(_09041_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17220_ (.I0(_02519_),
    .I1(\cs_registers_i.csr_mstatus_tw_o ),
    .S(_02678_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17221_ (.I0(_02517_),
    .I1(\cs_registers_i.mstatus_q[1] ),
    .S(_02678_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3564 (.I(net3558),
    .Z(net3564));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_167_clk_i_regs (.I(clknet_6_45__leaf_clk_i_regs),
    .Z(clknet_leaf_167_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17224_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_08626_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_169_clk_i_regs (.I(clknet_6_56__leaf_clk_i_regs),
    .Z(clknet_leaf_169_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_171_clk_i_regs (.I(clknet_6_56__leaf_clk_i_regs),
    .Z(clknet_leaf_171_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17227_ (.I0(\id_stage_i.controller_i.instr_i[0] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17228_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .A2(_02570_),
    .B1(_02681_),
    .B2(_02684_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _17229_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_08634_),
    .A3(_02570_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17230_ (.A1(_08724_),
    .A2(_02535_),
    .A3(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17231_ (.A1(_08985_),
    .A2(_02535_),
    .B1(_02685_),
    .B2(_02687_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17232_ (.I(_08938_),
    .ZN(_02689_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17233_ (.A1(_02143_),
    .A2(_02689_),
    .B(_02558_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_174_clk_i_regs (.I(clknet_6_56__leaf_clk_i_regs),
    .Z(clknet_leaf_174_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17235_ (.I0(\cs_registers_i.mtval_q[0] ),
    .I1(_02688_),
    .S(_02690_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_177_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_177_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17237_ (.A1(\cs_registers_i.pc_id_i[3] ),
    .A2(\cs_registers_i.pc_id_i[4] ),
    .A3(\cs_registers_i.pc_id_i[5] ),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17238_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .A4(_02693_),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17239_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(\cs_registers_i.pc_id_i[7] ),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17240_ (.A1(\cs_registers_i.pc_id_i[8] ),
    .A2(\cs_registers_i.pc_id_i[9] ),
    .A3(_02694_),
    .A4(_02695_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17241_ (.A1(\cs_registers_i.pc_id_i[10] ),
    .A2(_02696_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_178_clk_i_regs (.I(clknet_6_54__leaf_clk_i_regs),
    .Z(clknet_leaf_178_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17243_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17244_ (.A1(_02681_),
    .A2(_02699_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17245_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(net3289),
    .B1(_02697_),
    .B2(_08634_),
    .C(_02700_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17246_ (.A1(_09029_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02701_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17247_ (.I0(\cs_registers_i.mtval_q[10] ),
    .I1(_02702_),
    .S(_02690_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_179_clk_i_regs (.I(clknet_6_51__leaf_clk_i_regs),
    .Z(clknet_leaf_179_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17249_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17250_ (.A1(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .A2(_11167_[0]),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17251_ (.A1(_02693_),
    .A2(_02705_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17252_ (.A1(\cs_registers_i.pc_id_i[8] ),
    .A2(\cs_registers_i.pc_id_i[9] ),
    .A3(\cs_registers_i.pc_id_i[10] ),
    .A4(_02695_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17253_ (.A1(_02706_),
    .A2(_02707_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17254_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_02708_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_180_clk_i_regs (.I(clknet_6_51__leaf_clk_i_regs),
    .Z(clknet_leaf_180_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17256_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(net3289),
    .B1(_02681_),
    .B2(_02704_),
    .C1(_02709_),
    .C2(_08634_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17257_ (.A1(_09066_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02711_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17258_ (.I0(\cs_registers_i.mtval_q[11] ),
    .I1(_02712_),
    .S(_02690_),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17259_ (.I0(\id_stage_i.controller_i.instr_i[12] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17260_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_02694_),
    .A3(_02707_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17261_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_02714_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17262_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(net3289),
    .B1(_02681_),
    .B2(_02713_),
    .C1(_02715_),
    .C2(_08634_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17263_ (.A1(_09096_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02716_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17264_ (.I0(\cs_registers_i.mtval_q[12] ),
    .I1(_02717_),
    .S(_02690_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17265_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_02708_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17266_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_02718_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17267_ (.A1(\cs_registers_i.pc_id_i[13] ),
    .A2(_02719_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17268_ (.I0(\id_stage_i.controller_i.instr_i[13] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02721_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17269_ (.A1(_02681_),
    .A2(_02721_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17270_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(net3289),
    .B1(_02720_),
    .B2(_08634_),
    .C(_02722_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17271_ (.A1(_09117_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02723_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17272_ (.I0(\cs_registers_i.mtval_q[13] ),
    .I1(_02724_),
    .S(_02690_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17273_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(\cs_registers_i.pc_id_i[13] ),
    .A3(_02714_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17274_ (.A1(\cs_registers_i.pc_id_i[14] ),
    .A2(_02725_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17275_ (.I0(\id_stage_i.controller_i.instr_i[14] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17276_ (.A1(_02681_),
    .A2(_02727_),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17277_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(net3289),
    .B1(_02726_),
    .B2(_08634_),
    .C(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17278_ (.A1(_09133_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17279_ (.I0(\cs_registers_i.mtval_q[14] ),
    .I1(_02730_),
    .S(_02690_),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17280_ (.I0(net3607),
    .I1(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02731_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17281_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(\cs_registers_i.pc_id_i[13] ),
    .A3(\cs_registers_i.pc_id_i[14] ),
    .A4(_02718_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17282_ (.A1(\cs_registers_i.pc_id_i[15] ),
    .A2(_02732_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17283_ (.A1(_08634_),
    .A2(_02733_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17284_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(net3289),
    .B1(_02681_),
    .B2(_02731_),
    .C(_02734_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17285_ (.A1(_09149_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17286_ (.I0(\cs_registers_i.mtval_q[15] ),
    .I1(_02736_),
    .S(_02690_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3103 (.I(_03518_),
    .Z(net3103));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17288_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(\cs_registers_i.pc_id_i[13] ),
    .A3(\cs_registers_i.pc_id_i[14] ),
    .A4(\cs_registers_i.pc_id_i[15] ),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17289_ (.A1(_02714_),
    .A2(_02738_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17290_ (.A1(_07512_),
    .A2(_02739_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17291_ (.I(\id_stage_i.controller_i.instr_is_compressed_i ),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17292_ (.A1(_02741_),
    .A2(_02681_),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_182_clk_i_regs (.I(clknet_6_50__leaf_clk_i_regs),
    .Z(clknet_leaf_182_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17294_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(net3289),
    .B1(_02740_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3605),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17295_ (.A1(_09174_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02744_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17296_ (.I0(\cs_registers_i.mtval_q[16] ),
    .I1(_02745_),
    .S(_02690_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17297_ (.A1(_02718_),
    .A2(_02738_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17298_ (.A1(\cs_registers_i.pc_id_i[16] ),
    .A2(_02746_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17299_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(_02747_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_185_clk_i_regs (.I(clknet_6_49__leaf_clk_i_regs),
    .Z(clknet_leaf_185_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17301_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(net3289),
    .B1(_02748_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3582),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17302_ (.A1(_09194_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02750_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17303_ (.I0(\cs_registers_i.mtval_q[17] ),
    .I1(_02751_),
    .S(_02690_),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17304_ (.I(\cs_registers_i.pc_id_i[18] ),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17305_ (.A1(\cs_registers_i.pc_id_i[16] ),
    .A2(\cs_registers_i.pc_id_i[17] ),
    .A3(_02739_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17306_ (.A1(_02752_),
    .A2(_02753_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17307_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(net3289),
    .B1(_02754_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3580),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17308_ (.A1(_09210_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02755_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17309_ (.I0(\cs_registers_i.mtval_q[18] ),
    .I1(_02756_),
    .S(net3188),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17310_ (.A1(\cs_registers_i.pc_id_i[16] ),
    .A2(\cs_registers_i.pc_id_i[17] ),
    .A3(\cs_registers_i.pc_id_i[18] ),
    .A4(_02746_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17311_ (.A1(\cs_registers_i.pc_id_i[19] ),
    .A2(_02757_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17312_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(net3289),
    .B1(_02758_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3576),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17313_ (.A1(_09229_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_183_clk_i_regs (.I(clknet_6_50__leaf_clk_i_regs),
    .Z(clknet_leaf_183_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17315_ (.I0(\cs_registers_i.mtval_q[19] ),
    .I1(_02760_),
    .S(_02690_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_186_clk_i_regs (.I(clknet_6_48__leaf_clk_i_regs),
    .Z(clknet_leaf_186_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17317_ (.I0(net398),
    .I1(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17318_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17319_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A2(_02570_),
    .B1(_02681_),
    .B2(_02763_),
    .C1(_02764_),
    .C2(_08634_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17320_ (.A1(_09468_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02765_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17321_ (.I0(\cs_registers_i.mtval_q[1] ),
    .I1(_02766_),
    .S(_02690_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17322_ (.A1(\cs_registers_i.pc_id_i[16] ),
    .A2(\cs_registers_i.pc_id_i[17] ),
    .A3(\cs_registers_i.pc_id_i[18] ),
    .A4(\cs_registers_i.pc_id_i[19] ),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17323_ (.A1(_02739_),
    .A2(_02767_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17324_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(_02768_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17325_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(net3289),
    .B1(_02769_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3560),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17326_ (.A1(_09262_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02770_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17327_ (.I0(\cs_registers_i.mtval_q[20] ),
    .I1(_02771_),
    .S(_02690_),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17328_ (.A1(_02746_),
    .A2(_02767_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17329_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17330_ (.A1(\cs_registers_i.pc_id_i[21] ),
    .A2(_02773_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17331_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(net3289),
    .B1(_02774_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3552),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17332_ (.A1(_09277_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02775_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17333_ (.I0(\cs_registers_i.mtval_q[21] ),
    .I1(_02776_),
    .S(_02690_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_187_clk_i_regs (.I(clknet_6_49__leaf_clk_i_regs),
    .Z(clknet_leaf_187_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17335_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(\cs_registers_i.pc_id_i[21] ),
    .A3(_02768_),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17336_ (.A1(\cs_registers_i.pc_id_i[22] ),
    .A2(_02778_),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17337_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(net3289),
    .B1(_02779_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3499),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17338_ (.A1(_09293_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02780_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17339_ (.I0(\cs_registers_i.mtval_q[22] ),
    .I1(_02781_),
    .S(net3188),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17340_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(\cs_registers_i.pc_id_i[21] ),
    .A3(\cs_registers_i.pc_id_i[22] ),
    .A4(_02772_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17341_ (.A1(\cs_registers_i.pc_id_i[23] ),
    .A2(_02782_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17342_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(net3289),
    .B1(_02783_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3498),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17343_ (.A1(_09310_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17344_ (.I0(\cs_registers_i.mtval_q[23] ),
    .I1(_02785_),
    .S(net3188),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17345_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(\cs_registers_i.pc_id_i[21] ),
    .A3(\cs_registers_i.pc_id_i[22] ),
    .A4(\cs_registers_i.pc_id_i[23] ),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17346_ (.A1(_02768_),
    .A2(_02786_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17347_ (.A1(\cs_registers_i.pc_id_i[24] ),
    .A2(_02787_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17348_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(net3289),
    .B1(_02788_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3487),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17349_ (.A1(_09330_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17350_ (.I0(\cs_registers_i.mtval_q[24] ),
    .I1(_02790_),
    .S(net3188),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_188_clk_i_regs (.I(clknet_6_49__leaf_clk_i_regs),
    .Z(clknet_leaf_188_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17352_ (.A1(\cs_registers_i.pc_id_i[24] ),
    .A2(_02786_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17353_ (.A1(_02772_),
    .A2(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17354_ (.A1(\cs_registers_i.pc_id_i[25] ),
    .A2(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17355_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(net3289),
    .B1(_02794_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3486),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17356_ (.A1(_09348_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02795_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17357_ (.I0(\cs_registers_i.mtval_q[25] ),
    .I1(_02796_),
    .S(net3188),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17358_ (.A1(\cs_registers_i.pc_id_i[25] ),
    .A2(_02792_),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17359_ (.A1(_02768_),
    .A2(_02797_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17360_ (.A1(\cs_registers_i.pc_id_i[26] ),
    .A2(_02798_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17361_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(net3289),
    .B1(_02799_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3485),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17362_ (.A1(_09367_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02800_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17363_ (.I0(\cs_registers_i.mtval_q[26] ),
    .I1(_02801_),
    .S(net3188),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17364_ (.A1(\cs_registers_i.pc_id_i[26] ),
    .A2(_02797_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17365_ (.A1(_02772_),
    .A2(_02802_),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17366_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(_02803_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17367_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(net3289),
    .B1(_02804_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3484),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17368_ (.A1(_09384_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02805_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17369_ (.I0(\cs_registers_i.mtval_q[27] ),
    .I1(_02806_),
    .S(net3188),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17370_ (.A1(_02768_),
    .A2(_02802_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17371_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(_02807_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17372_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(_02808_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17373_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(net3289),
    .B1(_02809_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3483),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17374_ (.A1(_09401_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_191_clk_i_regs (.I(clknet_6_50__leaf_clk_i_regs),
    .Z(clknet_leaf_191_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17376_ (.I0(\cs_registers_i.mtval_q[28] ),
    .I1(_02811_),
    .S(net3188),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3563 (.I(net3558),
    .Z(net3563));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17378_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(\cs_registers_i.pc_id_i[28] ),
    .A3(_02803_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17379_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(_02814_),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17380_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(net3289),
    .B1(_02815_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3482),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17381_ (.A1(_09419_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02816_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17382_ (.I0(\cs_registers_i.mtval_q[29] ),
    .I1(_02817_),
    .S(net3188),
    .Z(_00407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17383_ (.I0(net3481),
    .I1(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17384_ (.I0(\cs_registers_i.pc_id_i[2] ),
    .I1(_11168_[0]),
    .S(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17385_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .A2(_02570_),
    .B1(_02681_),
    .B2(_02818_),
    .C1(_02819_),
    .C2(_08634_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17386_ (.A1(_09423_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02820_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17387_ (.I0(\cs_registers_i.mtval_q[2] ),
    .I1(_02821_),
    .S(_02690_),
    .Z(_00408_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17388_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(\cs_registers_i.pc_id_i[28] ),
    .A3(\cs_registers_i.pc_id_i[29] ),
    .A4(_02807_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17389_ (.A1(\cs_registers_i.pc_id_i[30] ),
    .A2(_02822_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17390_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(net3289),
    .B1(_02823_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3480),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17391_ (.A1(_09442_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02824_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17392_ (.I0(\cs_registers_i.mtval_q[30] ),
    .I1(_02825_),
    .S(_02690_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17393_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(\cs_registers_i.pc_id_i[28] ),
    .A3(\cs_registers_i.pc_id_i[29] ),
    .A4(\cs_registers_i.pc_id_i[30] ),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17394_ (.A1(_02803_),
    .A2(_02826_),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17395_ (.A1(\cs_registers_i.pc_id_i[31] ),
    .A2(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17396_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(net3289),
    .B1(_02828_),
    .B2(_08634_),
    .C1(_02742_),
    .C2(net3479),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17397_ (.A1(_09458_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17398_ (.I0(\cs_registers_i.mtval_q[31] ),
    .I1(_02830_),
    .S(_02690_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17399_ (.A1(\cs_registers_i.pc_id_i[3] ),
    .A2(_02705_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17400_ (.I0(net3478),
    .I1(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02832_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17401_ (.A1(_02681_),
    .A2(_02832_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17402_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A2(_02570_),
    .B1(_02831_),
    .B2(_08634_),
    .C(_02833_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17403_ (.A1(_09491_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02834_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17404_ (.I0(\cs_registers_i.mtval_q[3] ),
    .I1(_02835_),
    .S(_02690_),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17405_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(\cs_registers_i.pc_id_i[3] ),
    .A4(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Z(_02836_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17406_ (.A1(\cs_registers_i.pc_id_i[4] ),
    .A2(_02836_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17407_ (.I0(\id_stage_i.controller_i.instr_i[4] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17408_ (.A1(_02681_),
    .A2(_02838_),
    .Z(_02839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17409_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .A2(_02570_),
    .B1(_02837_),
    .B2(_08634_),
    .C(_02839_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17410_ (.A1(_09508_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02840_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17411_ (.I0(\cs_registers_i.mtval_q[4] ),
    .I1(_02841_),
    .S(_02690_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17412_ (.A1(\cs_registers_i.pc_id_i[3] ),
    .A2(\cs_registers_i.pc_id_i[4] ),
    .A3(_02705_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17413_ (.A1(\cs_registers_i.pc_id_i[5] ),
    .A2(_02842_),
    .Z(_02843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17414_ (.I0(\id_stage_i.controller_i.instr_i[5] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17415_ (.A1(_02681_),
    .A2(_02844_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17416_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(_02570_),
    .B1(_02843_),
    .B2(_08634_),
    .C(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17417_ (.A1(_09524_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02846_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17418_ (.I0(\cs_registers_i.mtval_q[5] ),
    .I1(_02847_),
    .S(_02690_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17419_ (.I0(net354),
    .I1(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17420_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(_02694_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17421_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(net3289),
    .B1(_02681_),
    .B2(_02848_),
    .C1(_02849_),
    .C2(_08634_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17422_ (.A1(_09541_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02850_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17423_ (.I0(\cs_registers_i.mtval_q[6] ),
    .I1(_02851_),
    .S(_02690_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17424_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(_02706_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17425_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17426_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17427_ (.A1(_02681_),
    .A2(_02854_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17428_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(net3289),
    .B1(_02853_),
    .B2(_08634_),
    .C(_02855_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17429_ (.A1(_09593_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02856_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17430_ (.I0(\cs_registers_i.mtval_q[7] ),
    .I1(_02857_),
    .S(_02690_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17431_ (.A1(_02694_),
    .A2(_02695_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17432_ (.A1(\cs_registers_i.pc_id_i[8] ),
    .A2(_02858_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17433_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17434_ (.A1(_02681_),
    .A2(_02860_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17435_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(net3289),
    .B1(_02859_),
    .B2(_08634_),
    .C(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17436_ (.A1(_09613_),
    .A2(_02535_),
    .B1(_02687_),
    .B2(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17437_ (.I0(\cs_registers_i.mtval_q[8] ),
    .I1(_02863_),
    .S(_02690_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17438_ (.A1(\cs_registers_i.pc_id_i[8] ),
    .A2(_02695_),
    .A3(_02706_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17439_ (.A1(\cs_registers_i.pc_id_i[9] ),
    .A2(_02864_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17440_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17441_ (.A1(_02681_),
    .A2(_02866_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17442_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(net3289),
    .B1(_02865_),
    .B2(_08634_),
    .C(_02867_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17443_ (.A1(_09628_),
    .A2(net3220),
    .B1(_02687_),
    .B2(_02868_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17444_ (.I0(\cs_registers_i.mtval_q[9] ),
    .I1(_02869_),
    .S(_02690_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17445_ (.A1(_08951_),
    .A2(_08926_),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_193_clk_i_regs (.I(clknet_6_39__leaf_clk_i_regs),
    .Z(clknet_leaf_193_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17447_ (.A1(_08361_),
    .A2(_08659_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_196_clk_i_regs (.I(clknet_6_39__leaf_clk_i_regs),
    .Z(clknet_leaf_196_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17449_ (.I(_02872_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17450_ (.A1(_02874_),
    .A2(_02870_),
    .Z(_02875_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_197_clk_i_regs (.I(clknet_6_39__leaf_clk_i_regs),
    .Z(clknet_leaf_197_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17452_ (.A1(net1),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[10] ),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17453_ (.A1(_09029_),
    .A2(_02870_),
    .B(_02877_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17454_ (.A1(net2),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[11] ),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17455_ (.A1(_09066_),
    .A2(_02870_),
    .B(_02878_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17456_ (.A1(net3),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[12] ),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17457_ (.A1(_09096_),
    .A2(_02870_),
    .B(_02879_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17458_ (.A1(net4),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[13] ),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17459_ (.A1(_09117_),
    .A2(_02870_),
    .B(_02880_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17460_ (.A1(net5),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[14] ),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17461_ (.A1(_09133_),
    .A2(_02870_),
    .B(_02881_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17462_ (.A1(net6),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[15] ),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17463_ (.A1(_09149_),
    .A2(_02870_),
    .B(_02882_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17464_ (.A1(net7),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[16] ),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17465_ (.A1(_09174_),
    .A2(_02870_),
    .B(_02883_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17466_ (.A1(net8),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[17] ),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17467_ (.A1(_09194_),
    .A2(_02870_),
    .B(_02884_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17468_ (.A1(net9),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[18] ),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17469_ (.A1(_09210_),
    .A2(_02870_),
    .B(_02885_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17470_ (.A1(net10),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[19] ),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17471_ (.A1(_09229_),
    .A2(_02870_),
    .B(_02886_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_198_clk_i_regs (.I(clknet_6_38__leaf_clk_i_regs),
    .Z(clknet_leaf_198_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_200_clk_i_regs (.I(clknet_6_39__leaf_clk_i_regs),
    .Z(clknet_leaf_200_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_201_clk_i_regs (.I(clknet_6_39__leaf_clk_i_regs),
    .Z(clknet_leaf_201_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17475_ (.A1(net11),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[20] ),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17476_ (.A1(_09262_),
    .A2(_02870_),
    .B(_02890_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17477_ (.A1(net12),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[21] ),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17478_ (.A1(_09277_),
    .A2(_02870_),
    .B(_02891_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17479_ (.A1(net13),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[22] ),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17480_ (.A1(_09293_),
    .A2(_02870_),
    .B(_02892_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17481_ (.A1(net14),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[23] ),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17482_ (.A1(_09310_),
    .A2(_02870_),
    .B(_02893_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17483_ (.A1(net15),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[24] ),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17484_ (.A1(_09330_),
    .A2(_02870_),
    .B(_02894_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17485_ (.A1(net16),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[25] ),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17486_ (.A1(_09348_),
    .A2(_02870_),
    .B(_02895_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17487_ (.A1(net17),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[26] ),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17488_ (.A1(_09367_),
    .A2(_02870_),
    .B(_02896_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17489_ (.A1(net18),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[27] ),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17490_ (.A1(_09384_),
    .A2(_02870_),
    .B(_02897_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17491_ (.A1(net19),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[28] ),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17492_ (.A1(_09401_),
    .A2(_02870_),
    .B(_02898_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17493_ (.A1(net20),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[29] ),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17494_ (.A1(_09419_),
    .A2(_02870_),
    .B(_02899_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17495_ (.A1(net21),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[30] ),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17496_ (.A1(_09442_),
    .A2(_02870_),
    .B(_02900_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17497_ (.A1(net22),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[31] ),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17498_ (.A1(_09458_),
    .A2(_02870_),
    .B(_02901_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17499_ (.A1(net23),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[8] ),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17500_ (.A1(_09613_),
    .A2(_02870_),
    .B(_02902_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17501_ (.A1(net24),
    .A2(_02872_),
    .B1(_02875_),
    .B2(\cs_registers_i.csr_mtvec_o[9] ),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17502_ (.A1(_09628_),
    .A2(_02870_),
    .B(_02903_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_202_clk_i_regs (.I(clknet_6_39__leaf_clk_i_regs),
    .Z(clknet_leaf_202_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17504_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_08407_),
    .A3(_08456_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17505_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .I1(_08445_),
    .S(_02905_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17506_ (.A1(net3647),
    .A2(net3371),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_205_clk_i_regs (.I(clknet_6_36__leaf_clk_i_regs),
    .Z(clknet_leaf_205_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17508_ (.A1(_08405_),
    .A2(_02906_),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _17509_ (.A1(net3655),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17510_ (.A1(_02908_),
    .A2(_02909_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17511_ (.I0(_08407_),
    .I1(_02910_),
    .S(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17512_ (.A1(_11172_[0]),
    .A2(_02909_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17513_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .I1(_02911_),
    .S(_08407_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17514_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(_11173_[0]),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17515_ (.A1(_02909_),
    .A2(_02912_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17516_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .I1(_02913_),
    .S(_08407_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17517_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17518_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_02914_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17519_ (.A1(_02909_),
    .A2(_02915_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17520_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .I1(_02916_),
    .S(_08407_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17521_ (.A1(_11173_[0]),
    .A2(_08402_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17522_ (.A1(_02909_),
    .A2(_02917_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17523_ (.A1(_02908_),
    .A2(_02918_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _17524_ (.A1(_11173_[0]),
    .A2(_08402_),
    .A3(_02908_),
    .A4(_02909_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17525_ (.I0(_02919_),
    .I1(_02920_),
    .S(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17526_ (.I0(\alu_adder_result_ex[0] ),
    .I1(net3376),
    .S(_08455_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17527_ (.A1(net3655),
    .A2(_08407_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_207_clk_i_regs (.I(clknet_6_36__leaf_clk_i_regs),
    .Z(clknet_leaf_207_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_208_clk_i_regs (.I(clknet_6_37__leaf_clk_i_regs),
    .Z(clknet_leaf_208_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17530_ (.I0(_02921_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .S(_02922_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_211_clk_i_regs (.I(clknet_6_31__leaf_clk_i_regs),
    .Z(clknet_leaf_211_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17532_ (.I0(net3312),
    .I1(net151),
    .S(_08458_),
    .Z(_02926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17533_ (.I0(_02926_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .S(_02922_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _17534_ (.I(net152),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_214_clk_i_regs (.I(clknet_6_36__leaf_clk_i_regs),
    .Z(clknet_leaf_214_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17536_ (.I0(net3377),
    .I1(_02927_),
    .S(_08458_),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17537_ (.I(_02929_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17538_ (.I0(_02930_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .S(_02922_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17539_ (.I(net153),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17540_ (.I0(net3381),
    .I1(_02931_),
    .S(_08458_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17541_ (.I(_02932_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17542_ (.I0(_02933_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .S(_02922_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17543_ (.I0(net3361),
    .I1(net154),
    .S(_08458_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17544_ (.I0(_02934_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .S(_02922_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17545_ (.I0(net3262),
    .I1(net365),
    .S(_08458_),
    .Z(_02935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17546_ (.I0(_02935_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .S(_02922_),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17547_ (.I0(net3350),
    .I1(net156),
    .S(_08458_),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_215_clk_i_regs (.I(clknet_6_36__leaf_clk_i_regs),
    .Z(clknet_leaf_215_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17549_ (.I0(_02936_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .S(_02922_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17550_ (.I0(net3360),
    .I1(net404),
    .S(_08458_),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17551_ (.I0(_02938_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .S(_02922_),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17552_ (.I0(net3349),
    .I1(_08436_),
    .S(_08458_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17553_ (.I(_02939_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17554_ (.I0(_02940_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .S(_02922_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_217_clk_i_regs (.I(clknet_6_5__leaf_clk_i_regs),
    .Z(clknet_leaf_217_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17556_ (.I0(net3359),
    .I1(net159),
    .S(_08458_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17557_ (.I0(_02942_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .S(_02922_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17558_ (.I0(net3283),
    .I1(net160),
    .S(_08458_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17559_ (.I0(_02943_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .S(_02922_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17560_ (.I0(net3355),
    .I1(\alu_adder_result_ex[1] ),
    .S(_08458_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17561_ (.I0(_02944_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .S(_02922_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17562_ (.I0(net3358),
    .I1(net161),
    .S(_08458_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17563_ (.I0(_02945_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .S(_02922_),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3562 (.I(net3558),
    .Z(net3562));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17565_ (.I0(net3347),
    .I1(_07787_),
    .S(_08458_),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17566_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .A2(_02922_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17567_ (.A1(_02922_),
    .A2(_02947_),
    .B(_02948_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17568_ (.I(net3346),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17569_ (.I0(_02949_),
    .I1(net163),
    .S(_08458_),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17570_ (.I0(_02950_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .S(_02922_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17571_ (.I0(net3277),
    .I1(net164),
    .S(_08458_),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17572_ (.I0(_02951_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .S(_02922_),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17573_ (.I(net3344),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17574_ (.I0(_02952_),
    .I1(net165),
    .S(_08458_),
    .Z(_02953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17575_ (.I0(_02953_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .S(_02922_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17576_ (.I(net3343),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17577_ (.I0(_02954_),
    .I1(net166),
    .S(_08458_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_219_clk_i_regs (.I(clknet_6_5__leaf_clk_i_regs),
    .Z(clknet_leaf_219_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17579_ (.I0(_02955_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .S(_02922_),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17580_ (.I0(net3342),
    .I1(_08078_),
    .S(_08458_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17581_ (.I(_02957_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17582_ (.I0(_02958_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .S(_02922_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17583_ (.A1(net168),
    .A2(_08455_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17584_ (.A1(net3357),
    .A2(_08455_),
    .B(_02959_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17585_ (.I0(_02960_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .S(_02922_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17586_ (.I(net169),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17587_ (.I0(net3341),
    .I1(_02961_),
    .S(_08458_),
    .Z(_02962_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17588_ (.I(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17589_ (.I0(_02963_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .S(_02922_),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17590_ (.I0(net3267),
    .I1(net170),
    .S(_08458_),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17591_ (.I0(_02964_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .S(_02922_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17592_ (.I0(net3372),
    .I1(net171),
    .S(_08458_),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17593_ (.I0(_02965_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .S(_02922_),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17594_ (.I0(net3261),
    .I1(net257),
    .S(_08458_),
    .Z(_02966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17595_ (.I0(_02966_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .S(_02922_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17596_ (.A1(net280),
    .A2(_08569_),
    .B(_08235_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17597_ (.I0(_02967_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .S(_02922_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17598_ (.I0(net3369),
    .I1(net174),
    .S(_08458_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17599_ (.I0(_02968_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .S(_02922_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17600_ (.I0(net3368),
    .I1(net175),
    .S(_08458_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17601_ (.I0(_02969_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .S(_02922_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17602_ (.I0(net3320),
    .I1(net176),
    .S(_08458_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17603_ (.I0(_02970_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .S(_02922_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17604_ (.A1(net177),
    .A2(_08458_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17605_ (.A1(net3366),
    .A2(_08458_),
    .B(_02971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17606_ (.I0(_02972_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .S(_02922_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17607_ (.I0(net3316),
    .I1(net178),
    .S(_08458_),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17608_ (.I0(_02973_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .S(_02922_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17609_ (.I(net179),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17610_ (.I0(net3364),
    .I1(_02974_),
    .S(_08458_),
    .Z(_02975_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17611_ (.I(_02975_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17612_ (.I0(_02976_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .S(_02922_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17613_ (.A1(net180),
    .A2(_08458_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17614_ (.A1(net3363),
    .A2(_08458_),
    .B(_02977_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17615_ (.I0(_02978_),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .S(_02922_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _17616_ (.A1(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .A2(_08252_),
    .A3(_08253_),
    .B(_08240_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17617_ (.A1(_08252_),
    .A2(net273),
    .B(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17618_ (.A1(_02979_),
    .A2(_02980_),
    .Z(_02981_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3104 (.I(_07258_),
    .Z(net3104));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3639 (.I(net3634),
    .Z(net3639));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17621_ (.A1(_08401_),
    .A2(_08402_),
    .A3(_02981_),
    .Z(_02984_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17622_ (.A1(_11171_[0]),
    .A2(_08407_),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17623_ (.A1(_02984_),
    .A2(_02985_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_222_clk_i_regs (.I(clknet_6_38__leaf_clk_i_regs),
    .Z(clknet_leaf_222_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17625_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17626_ (.A1(_02986_),
    .A2(_02988_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17627_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17628_ (.A1(_08401_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A3(_02989_),
    .A4(_02981_),
    .Z(_02990_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_226_clk_i_regs (.I(clknet_6_38__leaf_clk_i_regs),
    .Z(clknet_leaf_226_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17630_ (.A1(_11175_[0]),
    .A2(_08407_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17631_ (.A1(_02990_),
    .A2(_02992_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17632_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17633_ (.A1(_02993_),
    .A2(_02994_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17634_ (.A1(_11179_[0]),
    .A2(_08407_),
    .Z(_02995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17635_ (.A1(_02990_),
    .A2(_02995_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17636_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17637_ (.A1(_02996_),
    .A2(_02997_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17638_ (.A1(_08401_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A4(_02981_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_229_clk_i_regs (.I(clknet_6_33__leaf_clk_i_regs),
    .Z(clknet_leaf_229_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17640_ (.A1(_02985_),
    .A2(_02998_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17641_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17642_ (.A1(_03000_),
    .A2(_03001_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17643_ (.A1(_11177_[0]),
    .A2(_08407_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17644_ (.A1(_02998_),
    .A2(_03002_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17645_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17646_ (.A1(_03003_),
    .A2(_03004_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17647_ (.A1(_02992_),
    .A2(_02998_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17648_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17649_ (.A1(_03005_),
    .A2(_03006_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17650_ (.A1(_02995_),
    .A2(_02998_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17651_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17652_ (.A1(_03007_),
    .A2(_03008_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_230_clk_i_regs (.I(clknet_6_34__leaf_clk_i_regs),
    .Z(clknet_leaf_230_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17654_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(_08402_),
    .A3(_02981_),
    .Z(_03010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17655_ (.A1(_02985_),
    .A2(_03010_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17656_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17657_ (.A1(_03011_),
    .A2(_03012_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17658_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(_08409_),
    .A3(_02981_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17659_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .A2(_03013_),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17660_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .A2(_02922_),
    .B1(_03014_),
    .B2(net3654),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17661_ (.I(_03015_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17662_ (.A1(_02992_),
    .A2(_03010_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_231_clk_i_regs (.I(clknet_6_34__leaf_clk_i_regs),
    .Z(clknet_leaf_231_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17664_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17665_ (.A1(_03016_),
    .A2(_03018_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17666_ (.A1(_02995_),
    .A2(_03010_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_233_clk_i_regs (.I(clknet_6_32__leaf_clk_i_regs),
    .Z(clknet_leaf_233_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17668_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17669_ (.A1(_03019_),
    .A2(_03021_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17670_ (.A1(_08401_),
    .A2(_02981_),
    .Z(_03022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17671_ (.A1(_08409_),
    .A2(_03022_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17672_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .A2(_02922_),
    .B(net3654),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17673_ (.A1(_03023_),
    .A2(_03024_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17674_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_02989_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17675_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(_02979_),
    .A3(_02980_),
    .A4(_03025_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17676_ (.A1(_02985_),
    .A2(_03026_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17677_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17678_ (.A1(_03027_),
    .A2(_03028_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17679_ (.A1(_03002_),
    .A2(_03026_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17680_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17681_ (.A1(_03029_),
    .A2(_03030_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17682_ (.A1(_02992_),
    .A2(_03026_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17683_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17684_ (.A1(_03031_),
    .A2(_03032_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17685_ (.A1(_02995_),
    .A2(_03026_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17686_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17687_ (.A1(_03033_),
    .A2(_03034_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17688_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(_02989_),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17689_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_02979_),
    .A3(_02980_),
    .A4(_03035_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17690_ (.A1(_02985_),
    .A2(_03036_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17691_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17692_ (.A1(_03037_),
    .A2(_03038_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17693_ (.A1(_03002_),
    .A2(_03036_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17694_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17695_ (.A1(_03039_),
    .A2(_03040_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17696_ (.A1(_02992_),
    .A2(_03036_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17697_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17698_ (.A1(_03041_),
    .A2(_03042_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17699_ (.A1(_02995_),
    .A2(_03036_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_234_clk_i_regs (.I(clknet_6_33__leaf_clk_i_regs),
    .Z(clknet_leaf_234_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17701_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17702_ (.A1(_03043_),
    .A2(_03045_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17703_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A4(_02981_),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17704_ (.A1(_02985_),
    .A2(_03046_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3638 (.I(net3634),
    .Z(net3638));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17706_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17707_ (.A1(_03047_),
    .A2(_03049_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17708_ (.A1(_03002_),
    .A2(_03046_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17709_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17710_ (.A1(_03050_),
    .A2(_03051_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17711_ (.A1(_02984_),
    .A2(_02992_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17712_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17713_ (.A1(_03052_),
    .A2(_03053_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17714_ (.A1(_02992_),
    .A2(_03046_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17715_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17716_ (.A1(_03054_),
    .A2(_03055_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17717_ (.A1(_02995_),
    .A2(_03046_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17718_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17719_ (.A1(_03056_),
    .A2(_03057_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17720_ (.A1(_02984_),
    .A2(_02995_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17721_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17722_ (.A1(_03058_),
    .A2(_03059_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17723_ (.A1(_08401_),
    .A2(_02981_),
    .A3(_03025_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17724_ (.A1(_02985_),
    .A2(_03060_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17725_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .A2(_02922_),
    .B(net3654),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17726_ (.A1(_03061_),
    .A2(_03062_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17727_ (.A1(_03002_),
    .A2(_03060_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17728_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17729_ (.A1(_03063_),
    .A2(_03064_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17730_ (.A1(_02992_),
    .A2(_03060_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17731_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17732_ (.A1(_03065_),
    .A2(_03066_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17733_ (.A1(_02995_),
    .A2(_03060_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17734_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .A2(net3218),
    .B(net3654),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17735_ (.A1(_03067_),
    .A2(_03068_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17736_ (.A1(_02985_),
    .A2(_02990_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17737_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .A2(_02922_),
    .B(net3654),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17738_ (.A1(_03069_),
    .A2(_03070_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17739_ (.A1(_02990_),
    .A2(_03002_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17740_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .A2(_02922_),
    .B(net3654),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17741_ (.A1(_03071_),
    .A2(_03072_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17742_ (.A1(fetch_enable_q),
    .A2(net61),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_235_clk_i_regs (.I(clknet_6_32__leaf_clk_i_regs),
    .Z(clknet_leaf_235_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17744_ (.I0(net43),
    .I1(net27),
    .S(net3471),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17745_ (.I0(net57),
    .I1(net34),
    .S(net3471),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 _17746_ (.I(\load_store_unit_i.rdata_offset_q[1] ),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_237_clk_i_regs (.I(clknet_6_33__leaf_clk_i_regs),
    .Z(clknet_leaf_237_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17748_ (.I0(_03074_),
    .I1(_03075_),
    .S(_03076_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _17749_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(\load_store_unit_i.data_type_q[1] ),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_238_clk_i_regs (.I(clknet_6_33__leaf_clk_i_regs),
    .Z(clknet_leaf_238_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_241_clk_i_regs (.I(clknet_6_32__leaf_clk_i_regs),
    .Z(clknet_leaf_241_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_242_clk_i_regs (.I(clknet_6_32__leaf_clk_i_regs),
    .Z(clknet_leaf_242_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_244_clk_i_regs (.I(clknet_6_32__leaf_clk_i_regs),
    .Z(clknet_leaf_244_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17754_ (.I0(net57),
    .I1(\load_store_unit_i.rdata_q[8] ),
    .I2(\load_store_unit_i.rdata_q[16] ),
    .I3(net27),
    .S0(net3471),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17755_ (.I0(net56),
    .I1(net42),
    .I2(net33),
    .I3(net51),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17756_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(\load_store_unit_i.data_sign_ext_q ),
    .A3(_03085_),
    .Z(_03086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17757_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_03078_),
    .B1(_03079_),
    .B2(_03084_),
    .C(_03086_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17758_ (.I(_03087_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17759_ (.A1(_06993_),
    .A2(_07003_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17760_ (.A1(_07004_),
    .A2(_01953_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _17761_ (.A1(_11004_[0]),
    .A2(_03089_),
    .A3(_03090_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17762_ (.A1(_06388_),
    .A2(net484),
    .A3(_11410_[0]),
    .B(_06253_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17763_ (.A1(net3288),
    .A2(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_247_clk_i_regs (.I(clknet_6_13__leaf_clk_i_regs),
    .Z(clknet_leaf_247_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_248_clk_i_regs (.I(clknet_6_12__leaf_clk_i_regs),
    .Z(clknet_leaf_248_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17766_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A2(_06398_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _17767_ (.A1(_06404_),
    .A2(_06414_),
    .A3(_06438_),
    .Z(_03097_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17768_ (.A1(_11394_[0]),
    .A2(net299),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _17769_ (.A1(_06253_),
    .A2(_03096_),
    .A3(_03097_),
    .B(_03098_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _17770_ (.A1(_11004_[0]),
    .A2(_06993_),
    .A3(_07003_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_250_clk_i_regs (.I(clknet_6_13__leaf_clk_i_regs),
    .Z(clknet_leaf_250_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17772_ (.I0(_11437_[0]),
    .I1(_11453_[0]),
    .I2(_11602_[0]),
    .I3(_11586_[0]),
    .S0(net3207),
    .S1(_03100_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17773_ (.I0(_11429_[0]),
    .I1(_11445_[0]),
    .I2(_11610_[0]),
    .I3(_11594_[0]),
    .S0(net3207),
    .S1(_03100_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17774_ (.I0(_03102_),
    .I1(_03103_),
    .S(_06388_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_251_clk_i_regs (.I(clknet_6_13__leaf_clk_i_regs),
    .Z(clknet_leaf_251_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _17776_ (.I0(_11399_[0]),
    .I1(_11406_[0]),
    .I2(_11139_[0]),
    .I3(_11634_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17777_ (.I0(_11413_[0]),
    .I1(_11421_[0]),
    .I2(_11626_[0]),
    .I3(_11618_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3098 (.I(_03699_),
    .Z(net3098));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17779_ (.I0(_03106_),
    .I1(_03107_),
    .S(net3207),
    .Z(_03109_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17780_ (.A1(_11393_[0]),
    .A2(net299),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17781_ (.A1(_11414_[0]),
    .A2(_03110_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3097 (.I(net155),
    .Z(net3097));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17783_ (.I0(_03104_),
    .I1(_03109_),
    .S(_03111_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17784_ (.A1(_11004_[0]),
    .A2(_06993_),
    .A3(_07003_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_252_clk_i_regs (.I(clknet_6_32__leaf_clk_i_regs),
    .Z(clknet_leaf_252_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17786_ (.I0(_11485_[0]),
    .I1(_11477_[0]),
    .I2(_11554_[0]),
    .I3(_11562_[0]),
    .S0(net3253),
    .S1(_03114_),
    .Z(_03116_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_254_clk_i_regs (.I(clknet_6_40__leaf_clk_i_regs),
    .Z(clknet_leaf_254_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17788_ (.I0(_11461_[0]),
    .I1(_11469_[0]),
    .I2(_11578_[0]),
    .I3(_11570_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17789_ (.I0(_03116_),
    .I1(_03118_),
    .S(net3207),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17790_ (.I0(_11514_[0]),
    .I1(_11522_[0]),
    .S(_03114_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17791_ (.I0(_11498_[0]),
    .I1(_11538_[0]),
    .S(_03114_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17792_ (.I0(_11506_[0]),
    .I1(_11530_[0]),
    .S(_03114_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17793_ (.I0(_11490_[0]),
    .I1(_11546_[0]),
    .S(_03114_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17794_ (.I0(_03120_),
    .I1(_03121_),
    .I2(_03122_),
    .I3(_03123_),
    .S0(net3207),
    .S1(net3253),
    .Z(_03124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17795_ (.I0(_03119_),
    .I1(_03124_),
    .S(_03111_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17796_ (.A1(_11393_[0]),
    .A2(_08930_),
    .B(net299),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17797_ (.A1(_06530_),
    .A2(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_255_clk_i_regs (.I(clknet_6_40__leaf_clk_i_regs),
    .Z(clknet_leaf_255_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17799_ (.I0(_03113_),
    .I1(_03125_),
    .S(_03127_),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17800_ (.A1(_03093_),
    .A2(_03129_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17801_ (.A1(net3287),
    .A2(_03126_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _17802_ (.A1(_09743_),
    .A2(_06895_),
    .A3(_06918_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _17803_ (.A1(_11004_[0]),
    .A2(_08201_),
    .A3(_08216_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17804_ (.A1(_01923_),
    .A2(_03089_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17805_ (.A1(_03132_),
    .A2(_03133_),
    .B(_03134_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_256_clk_i_regs (.I(clknet_6_40__leaf_clk_i_regs),
    .Z(clknet_leaf_256_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17807_ (.A1(_03131_),
    .A2(_03135_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17808_ (.I0(_11490_[0]),
    .I1(_11498_[0]),
    .I2(_11546_[0]),
    .I3(_11538_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17809_ (.I0(_11461_[0]),
    .I1(_11469_[0]),
    .I2(_11578_[0]),
    .I3(_11570_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17810_ (.I0(_11510_[0]),
    .I1(_11534_[0]),
    .S(_03100_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17811_ (.A1(_11522_[0]),
    .A2(_03100_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_258_clk_i_regs (.I(clknet_6_41__leaf_clk_i_regs),
    .Z(clknet_leaf_258_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17813_ (.A1(_11514_[0]),
    .A2(_03114_),
    .B(_06388_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17814_ (.A1(_06388_),
    .A2(_03140_),
    .B1(_03141_),
    .B2(_03143_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17815_ (.I0(_11485_[0]),
    .I1(_11477_[0]),
    .I2(_11554_[0]),
    .I3(_11562_[0]),
    .S0(_06388_),
    .S1(_03100_),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_260_clk_i_regs (.I(clknet_6_32__leaf_clk_i_regs),
    .Z(clknet_leaf_260_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _17817_ (.I0(_03138_),
    .I1(_03139_),
    .I2(_03144_),
    .I3(_03145_),
    .S0(_03111_),
    .S1(net3207),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17818_ (.A1(_03127_),
    .A2(_03147_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17819_ (.A1(_03137_),
    .A2(_03148_),
    .B(_03093_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17820_ (.A1(_03091_),
    .A2(_03130_),
    .A3(_03149_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17821_ (.A1(net3126),
    .A2(net3160),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _17822_ (.A1(net3657),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A3(_08471_),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_262_clk_i_regs (.I(clknet_6_41__leaf_clk_i_regs),
    .Z(clknet_leaf_262_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17824_ (.A1(net3417),
    .A2(_03152_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_263_clk_i_regs (.I(clknet_6_34__leaf_clk_i_regs),
    .Z(clknet_leaf_263_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17826_ (.I0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .I1(_03151_),
    .S(_03154_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_264_clk_i_regs (.I(clknet_6_34__leaf_clk_i_regs),
    .Z(clknet_leaf_264_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17828_ (.A1(_03132_),
    .A2(_03133_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17829_ (.A1(_03158_),
    .A2(_03134_),
    .Z(_03159_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _17830_ (.A1(_06895_),
    .A2(_06918_),
    .A3(_03100_),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _17831_ (.A1(_08201_),
    .A2(_08216_),
    .A3(_03114_),
    .Z(_03161_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17832_ (.A1(_03160_),
    .A2(_03161_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17833_ (.A1(_11414_[0]),
    .A2(_03110_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_265_clk_i_regs (.I(clknet_6_34__leaf_clk_i_regs),
    .Z(clknet_leaf_265_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17835_ (.A1(_03163_),
    .A2(net3207),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17836_ (.A1(_06388_),
    .A2(_03162_),
    .A3(_03165_),
    .B(_03135_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17837_ (.I0(_11433_[0]),
    .I1(_11606_[0]),
    .S(_03100_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17838_ (.I0(_11449_[0]),
    .I1(_11590_[0]),
    .S(_03100_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17839_ (.I0(_11441_[0]),
    .I1(_11598_[0]),
    .S(_03100_),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17840_ (.I0(_11457_[0]),
    .I1(_11582_[0]),
    .S(_03100_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _17841_ (.I0(_03167_),
    .I1(_03168_),
    .I2(_03169_),
    .I3(_03170_),
    .S0(net3207),
    .S1(net3253),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _17842_ (.I0(_11402_[0]),
    .I1(_11409_[0]),
    .I2(_11638_[0]),
    .I3(_11630_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17843_ (.I0(_11417_[0]),
    .I1(net3252),
    .I2(_11622_[0]),
    .I3(_11614_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17844_ (.I0(_03172_),
    .I1(_03173_),
    .S(net3207),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17845_ (.I0(_03171_),
    .I1(_03174_),
    .S(_03111_),
    .Z(_03175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17846_ (.I0(_03166_),
    .I1(_03175_),
    .S(_03093_),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17847_ (.I0(_03159_),
    .I1(_03176_),
    .S(_03127_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17848_ (.I(_11463_[0]),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17849_ (.A1(_11004_[0]),
    .A2(_09742_),
    .B(_01922_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _17850_ (.A1(net3383),
    .A2(_07294_),
    .A3(_03179_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _17851_ (.A1(net3383),
    .A2(_07000_),
    .A3(_07294_),
    .A4(_01953_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17852_ (.I(_03181_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _17853_ (.A1(net3383),
    .A2(_07294_),
    .A3(_03179_),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17854_ (.A1(_11004_[0]),
    .A2(_01921_),
    .Z(_03184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17855_ (.I0(_11012_[0]),
    .I1(_03184_),
    .S(_01931_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17856_ (.A1(_07003_),
    .A2(_03185_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17857_ (.A1(_03182_),
    .A2(_03183_),
    .A3(_03186_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17858_ (.A1(_03178_),
    .A2(_03180_),
    .B1(_03187_),
    .B2(_11460_[0]),
    .C1(_11459_[0]),
    .C2(_03181_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17859_ (.A1(_01923_),
    .A2(_07004_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _17860_ (.A1(_01921_),
    .A2(_01931_),
    .A3(_07003_),
    .A4(_03189_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_266_clk_i_regs (.I(clknet_6_44__leaf_clk_i_regs),
    .Z(clknet_leaf_266_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17862_ (.A1(net179),
    .A2(_03190_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17863_ (.A1(net3215),
    .A2(_01916_),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17864_ (.A1(_09742_),
    .A2(_03193_),
    .B(_01948_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17865_ (.A1(_07295_),
    .A2(_03194_),
    .B(_01956_),
    .C(_01920_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17866_ (.A1(_01952_),
    .A2(_01953_),
    .B(_03089_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17867_ (.A1(_03186_),
    .A2(_03190_),
    .A3(_03196_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _17868_ (.A1(_03195_),
    .A2(_03181_),
    .A3(_03180_),
    .A4(_03197_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _17869_ (.A1(net3374),
    .A2(_03198_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17870_ (.A1(_03188_),
    .A2(_03192_),
    .B(_03199_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17871_ (.A1(net3373),
    .A2(_03156_),
    .B1(_03114_),
    .B2(_03177_),
    .C(_03200_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17872_ (.A1(_08265_),
    .A2(_03150_),
    .A3(_03201_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17873_ (.A1(_06718_),
    .A2(_09611_),
    .B(_03202_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17874_ (.A1(net263),
    .A2(_08351_),
    .A3(_08348_),
    .A4(_08349_),
    .Z(_03204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17875_ (.A1(_08352_),
    .A2(_03204_),
    .B(_08356_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _17876_ (.A1(_08332_),
    .A2(_08341_),
    .A3(_08347_),
    .A4(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17877_ (.A1(_11410_[0]),
    .A2(_08274_),
    .A3(_08287_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17878_ (.I(_08324_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _17879_ (.A1(_08305_),
    .A2(_08306_),
    .A3(_08311_),
    .B1(_08299_),
    .B2(_03208_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17880_ (.A1(_06530_),
    .A2(_08299_),
    .A3(_08303_),
    .B(_11410_[0]),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17881_ (.A1(_06388_),
    .A2(net485),
    .B(_11410_[0]),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17882_ (.A1(_08896_),
    .A2(_03209_),
    .B(_03210_),
    .C(_03211_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17883_ (.A1(_03207_),
    .A2(_03212_),
    .B(_11418_[0]),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17884_ (.A1(_03206_),
    .A2(_03213_),
    .B(_08950_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17885_ (.A1(_06323_),
    .A2(_06346_),
    .B(_06393_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17886_ (.I(_03215_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _17887_ (.A1(_06782_),
    .A2(_08404_),
    .A3(_08365_),
    .A4(_01967_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17888_ (.A1(_03214_),
    .A2(_03216_),
    .B(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_269_clk_i_regs (.I(clknet_6_44__leaf_clk_i_regs),
    .Z(clknet_leaf_269_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place3096 (.I(_03745_),
    .Z(net3096));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17891_ (.I0(_03088_),
    .I1(_03203_),
    .S(_03218_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_276_clk_i_regs (.I(clknet_6_43__leaf_clk_i_regs),
    .Z(clknet_leaf_276_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17893_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _17894_ (.A1(net25),
    .A2(\load_store_unit_i.lsu_err_q ),
    .A3(\load_store_unit_i.data_we_q ),
    .A4(_08396_),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17895_ (.A1(_08326_),
    .A2(_08358_),
    .B(_08373_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _17896_ (.A1(_11154_[0]),
    .A2(_08359_),
    .A3(_08364_),
    .A4(_09586_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _17897_ (.A1(_03226_),
    .A2(_08405_),
    .A3(_01967_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _17898_ (.A1(_03225_),
    .A2(_03215_),
    .B(_03227_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17899_ (.A1(_03224_),
    .A2(_03228_),
    .B(_06739_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17900_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .Z(_03230_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17901_ (.A1(_03229_),
    .A2(_03230_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17902_ (.A1(_03223_),
    .A2(_03231_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_277_clk_i_regs (.I(clknet_6_43__leaf_clk_i_regs),
    .Z(clknet_leaf_277_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17904_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .I1(net3090),
    .S(_03232_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_278_clk_i_regs (.I(clknet_6_43__leaf_clk_i_regs),
    .Z(clknet_leaf_278_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_280_clk_i_regs (.I(clknet_6_46__leaf_clk_i_regs),
    .Z(clknet_leaf_280_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_281_clk_i_regs (.I(clknet_6_43__leaf_clk_i_regs),
    .Z(clknet_leaf_281_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17908_ (.I0(net58),
    .I1(\load_store_unit_i.rdata_q[9] ),
    .I2(\load_store_unit_i.rdata_q[17] ),
    .I3(net38),
    .S0(net3471),
    .S1(net3470),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_283_clk_i_regs (.I(clknet_6_46__leaf_clk_i_regs),
    .Z(clknet_leaf_283_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17910_ (.I0(net44),
    .I1(net38),
    .S(net3471),
    .Z(_03239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17911_ (.I0(net58),
    .I1(net35),
    .S(net3471),
    .Z(_03240_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_282_clk_i_regs (.I(clknet_6_46__leaf_clk_i_regs),
    .Z(clknet_leaf_282_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17913_ (.I0(_03239_),
    .I1(_03240_),
    .S(_03076_),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17914_ (.A1(_03218_),
    .A2(_03086_),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17915_ (.A1(_03079_),
    .A2(_03237_),
    .B1(_03242_),
    .B2(\load_store_unit_i.data_type_q[2] ),
    .C(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _17916_ (.A1(_11004_[0]),
    .A2(_03089_),
    .A3(_03090_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_284_clk_i_regs (.I(clknet_6_43__leaf_clk_i_regs),
    .Z(clknet_leaf_284_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_285_clk_i_regs (.I(clknet_6_43__leaf_clk_i_regs),
    .Z(clknet_leaf_285_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17919_ (.A1(_11418_[0]),
    .A2(_03092_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_286_clk_i_regs (.I(clknet_6_43__leaf_clk_i_regs),
    .Z(clknet_leaf_286_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_287_clk_i_regs (.I(clknet_6_42__leaf_clk_i_regs),
    .Z(clknet_leaf_287_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17922_ (.I0(_11494_[0]),
    .I1(_11481_[0]),
    .I2(_11550_[0]),
    .I3(_11558_[0]),
    .S0(net3253),
    .S1(_03114_),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17923_ (.I0(_11465_[0]),
    .I1(_11473_[0]),
    .I2(_11574_[0]),
    .I3(_11566_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17924_ (.I0(_03251_),
    .I1(_03252_),
    .S(net3207),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17925_ (.A1(net3253),
    .A2(_03114_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17926_ (.I0(_11518_[0]),
    .I1(_11526_[0]),
    .S(_03254_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17927_ (.I0(_11502_[0]),
    .I1(_11542_[0]),
    .S(_03114_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17928_ (.I0(_11510_[0]),
    .I1(_11534_[0]),
    .S(_03114_),
    .Z(_03257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17929_ (.I0(_03256_),
    .I1(_03257_),
    .S(_06388_),
    .Z(_03258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17930_ (.I0(_03255_),
    .I1(_03258_),
    .S(net3207),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17931_ (.I0(_03253_),
    .I1(_03259_),
    .S(_03111_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17932_ (.I0(_11494_[0]),
    .I1(_11481_[0]),
    .I2(_11550_[0]),
    .I3(_11558_[0]),
    .S0(_06388_),
    .S1(_03100_),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17933_ (.I0(_11502_[0]),
    .I1(_11542_[0]),
    .S(_03100_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17934_ (.I0(_03262_),
    .I1(_03140_),
    .S(net3253),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_288_clk_i_regs (.I(clknet_6_42__leaf_clk_i_regs),
    .Z(clknet_leaf_288_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17936_ (.I0(_11449_[0]),
    .I1(_11457_[0]),
    .I2(_11590_[0]),
    .I3(_11582_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17937_ (.I0(_11465_[0]),
    .I1(_11473_[0]),
    .I2(_11574_[0]),
    .I3(_11566_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17938_ (.I0(_03261_),
    .I1(_03263_),
    .I2(_03265_),
    .I3(_03266_),
    .S0(net3207),
    .S1(_03111_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17939_ (.A1(_03093_),
    .A2(_03267_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17940_ (.A1(_03248_),
    .A2(_03260_),
    .B(_03268_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_289_clk_i_regs (.I(clknet_6_42__leaf_clk_i_regs),
    .Z(clknet_leaf_289_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17942_ (.I0(_11417_[0]),
    .I1(_11622_[0]),
    .S(_03100_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17943_ (.I0(net3252),
    .I1(_11614_[0]),
    .S(_03100_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17944_ (.I0(_11394_[0]),
    .I1(_06440_),
    .S(net299),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17945_ (.I0(_03167_),
    .I1(_03169_),
    .I2(_03271_),
    .I3(_03272_),
    .S0(net3253),
    .S1(_03273_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17946_ (.A1(_03163_),
    .A2(_03274_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_294_clk_i_regs (.I(clknet_6_42__leaf_clk_i_regs),
    .Z(clknet_leaf_294_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17948_ (.A1(_03273_),
    .A2(_03172_),
    .Z(_03277_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17949_ (.A1(_06388_),
    .A2(_03162_),
    .B(_03273_),
    .C(_03135_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17950_ (.A1(_03111_),
    .A2(_03277_),
    .A3(_03278_),
    .Z(_03279_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _17951_ (.A1(_03275_),
    .A2(_03279_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17952_ (.A1(_03131_),
    .A2(_03135_),
    .Z(_03281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17953_ (.A1(_03248_),
    .A2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17954_ (.A1(_03127_),
    .A2(_03248_),
    .A3(_03280_),
    .B(_03282_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17955_ (.A1(_03127_),
    .A2(_03269_),
    .B(_03283_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_292_clk_i_regs (.I(clknet_6_42__leaf_clk_i_regs),
    .Z(clknet_leaf_292_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17957_ (.I0(_11445_[0]),
    .I1(_11453_[0]),
    .I2(_11594_[0]),
    .I3(_11586_[0]),
    .S0(net3253),
    .S1(_03100_),
    .Z(_03286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17958_ (.I0(_03139_),
    .I1(_03286_),
    .S(_03273_),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17959_ (.I0(_11421_[0]),
    .I1(_11437_[0]),
    .I2(_11618_[0]),
    .I3(_11602_[0]),
    .S0(net3207),
    .S1(_03100_),
    .Z(_03288_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17960_ (.I0(_11413_[0]),
    .I1(_11429_[0]),
    .I2(_11626_[0]),
    .I3(_11610_[0]),
    .S0(net3207),
    .S1(_03100_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17961_ (.I0(_03288_),
    .I1(_03289_),
    .S(_06388_),
    .Z(_03290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17962_ (.I0(_03287_),
    .I1(_03290_),
    .S(_03111_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17963_ (.A1(_03163_),
    .A2(net3207),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17964_ (.I0(_03135_),
    .I1(_03106_),
    .S(_03292_),
    .Z(_03293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17965_ (.I0(_03291_),
    .I1(_03293_),
    .S(_03248_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17966_ (.A1(_03131_),
    .A2(_03159_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17967_ (.A1(_03131_),
    .A2(_03294_),
    .B(_03295_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_295_clk_i_regs (.I(clknet_6_15__leaf_clk_i_regs),
    .Z(clknet_leaf_295_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _17969_ (.A1(net3374),
    .A2(_03198_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_296_clk_i_regs (.I(clknet_6_14__leaf_clk_i_regs),
    .Z(clknet_leaf_296_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17971_ (.A1(net180),
    .A2(_03190_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_297_clk_i_regs (.I(clknet_6_14__leaf_clk_i_regs),
    .Z(clknet_leaf_297_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_304_clk_i_regs (.I(clknet_6_40__leaf_clk_i_regs),
    .Z(clknet_leaf_304_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17974_ (.A1(_11471_[0]),
    .A2(_03183_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17975_ (.A1(_11467_[0]),
    .A2(_03181_),
    .B1(_03187_),
    .B2(_11468_[0]),
    .C(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17976_ (.A1(_03300_),
    .A2(_03304_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17977_ (.I(_11236_[0]),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17978_ (.A1(net3161),
    .A2(_11227_[0]),
    .B(_11226_[0]),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17979_ (.I(_11235_[0]),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17980_ (.A1(_03306_),
    .A2(_03307_),
    .B(_03308_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17981_ (.A1(net3157),
    .A2(net3130),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17982_ (.I0(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .I1(_03310_),
    .S(_03154_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17983_ (.A1(_03298_),
    .A2(_03305_),
    .B1(_03311_),
    .B2(net3370),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17984_ (.A1(_09626_),
    .A2(_03218_),
    .A3(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17985_ (.A1(_03245_),
    .A2(_03284_),
    .B1(_03296_),
    .B2(_03114_),
    .C(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _17986_ (.A1(_03244_),
    .A2(_03314_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_299_clk_i_regs (.I(clknet_6_15__leaf_clk_i_regs),
    .Z(clknet_leaf_299_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17988_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .I1(_03315_),
    .S(_03232_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17989_ (.A1(_03245_),
    .A2(_03282_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17990_ (.I0(_03138_),
    .I1(_03145_),
    .S(_03273_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17991_ (.I0(_03287_),
    .I1(_03318_),
    .S(_03163_),
    .Z(_03319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17992_ (.I0(_03120_),
    .I1(_03122_),
    .S(net3253),
    .Z(_03320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17993_ (.I0(_03144_),
    .I1(_03320_),
    .S(net3207),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17994_ (.I0(_11494_[0]),
    .I1(_11550_[0]),
    .S(_03114_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17995_ (.I0(_03256_),
    .I1(_03322_),
    .S(net3253),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17996_ (.I0(_11481_[0]),
    .I1(_11473_[0]),
    .I2(_11558_[0]),
    .I3(_11566_[0]),
    .S0(net3253),
    .S1(_03114_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17997_ (.A1(net3207),
    .A2(_03324_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17998_ (.A1(_03273_),
    .A2(_03323_),
    .B(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_303_clk_i_regs (.I(clknet_6_15__leaf_clk_i_regs),
    .Z(clknet_leaf_303_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18000_ (.I0(_03321_),
    .I1(_03326_),
    .S(_03163_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18001_ (.I0(_03319_),
    .I1(_03328_),
    .S(_03093_),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18002_ (.I0(_03135_),
    .I1(_03106_),
    .S(net3207),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18003_ (.I0(_03290_),
    .I1(_03330_),
    .S(_03111_),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18004_ (.A1(_03093_),
    .A2(_03331_),
    .Z(_03332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18005_ (.I0(_03329_),
    .I1(_03332_),
    .S(_03131_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_301_clk_i_regs (.I(clknet_6_15__leaf_clk_i_regs),
    .Z(clknet_leaf_301_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_302_clk_i_regs (.I(clknet_6_15__leaf_clk_i_regs),
    .Z(clknet_leaf_302_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_306_clk_i_regs (.I(clknet_6_15__leaf_clk_i_regs),
    .Z(clknet_leaf_306_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18009_ (.A1(_03306_),
    .A2(_09859_[0]),
    .B(_03308_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18010_ (.A1(_11245_[0]),
    .A2(_03337_),
    .B(net3158),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18011_ (.A1(net3156),
    .A2(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18012_ (.I0(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .I1(_03339_),
    .S(_03154_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18013_ (.A1(net3370),
    .A2(_03340_),
    .B(_06718_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_307_clk_i_regs (.I(clknet_6_13__leaf_clk_i_regs),
    .Z(clknet_leaf_307_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_308_clk_i_regs (.I(clknet_6_13__leaf_clk_i_regs),
    .Z(clknet_leaf_308_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18016_ (.A1(_11475_[0]),
    .A2(_03181_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18017_ (.A1(_11479_[0]),
    .A2(_03183_),
    .B(_03341_),
    .C(_03344_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18018_ (.A1(net151),
    .A2(_03190_),
    .B1(_03187_),
    .B2(_11476_[0]),
    .C(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18019_ (.A1(_03114_),
    .A2(_03137_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18020_ (.A1(_03160_),
    .A2(_03161_),
    .B(_06388_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18021_ (.A1(_03348_),
    .A2(net3207),
    .B(_03163_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18022_ (.A1(_03165_),
    .A2(_03172_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18023_ (.A1(_03135_),
    .A2(_03349_),
    .B(_03350_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18024_ (.I0(_03266_),
    .I1(_03265_),
    .S(_03273_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18025_ (.I0(_03352_),
    .I1(_03274_),
    .S(_03111_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18026_ (.I0(_03351_),
    .I1(_03353_),
    .S(_03093_),
    .Z(_03354_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18027_ (.A1(_03131_),
    .A2(_03354_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18028_ (.A1(_03347_),
    .A2(_03355_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18029_ (.A1(_03317_),
    .A2(_03333_),
    .B(_03346_),
    .C(_03356_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_309_clk_i_regs (.I(clknet_6_12__leaf_clk_i_regs),
    .Z(clknet_leaf_309_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18031_ (.A1(_06718_),
    .A2(_09023_),
    .B1(_03199_),
    .B2(_03341_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18032_ (.A1(_03357_),
    .A2(_03359_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_310_clk_i_regs (.I(clknet_6_15__leaf_clk_i_regs),
    .Z(clknet_leaf_310_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_311_clk_i_regs (.I(clknet_6_12__leaf_clk_i_regs),
    .Z(clknet_leaf_311_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18035_ (.I0(net28),
    .I1(\load_store_unit_i.rdata_q[10] ),
    .I2(\load_store_unit_i.rdata_q[18] ),
    .I3(net49),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(net3470),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18036_ (.I0(net45),
    .I1(net49),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18037_ (.I0(net28),
    .I1(net36),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18038_ (.I0(_03364_),
    .I1(_03365_),
    .S(_03076_),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18039_ (.A1(net3400),
    .A2(_03363_),
    .B1(_03366_),
    .B2(\load_store_unit_i.data_type_q[2] ),
    .C(_03243_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18040_ (.A1(_03218_),
    .A2(_03360_),
    .B(_03367_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_312_clk_i_regs (.I(clknet_6_12__leaf_clk_i_regs),
    .Z(clknet_leaf_312_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18042_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .I1(net3089),
    .S(_03232_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18043_ (.I0(_03261_),
    .I1(_03266_),
    .S(_03273_),
    .Z(_03370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18044_ (.I0(_03263_),
    .I1(_03255_),
    .S(net3207),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18045_ (.I0(_03251_),
    .I1(_03258_),
    .S(_03273_),
    .Z(_03372_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18046_ (.I0(_03171_),
    .I1(_03370_),
    .I2(_03371_),
    .I3(_03372_),
    .S0(_03163_),
    .S1(_03093_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_317_clk_i_regs (.I(clknet_6_14__leaf_clk_i_regs),
    .Z(clknet_leaf_317_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18048_ (.A1(_06388_),
    .A2(_03162_),
    .A3(_03273_),
    .B(_03135_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18049_ (.I0(_03174_),
    .I1(_03375_),
    .S(_03111_),
    .Z(_03376_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18050_ (.A1(_03127_),
    .A2(_03248_),
    .A3(_03376_),
    .Z(_03377_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18051_ (.A1(_03131_),
    .A2(_03373_),
    .B(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18052_ (.A1(_03317_),
    .A2(_03378_),
    .Z(_03379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18053_ (.I0(_03139_),
    .I1(_03145_),
    .S(net3207),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18054_ (.I0(_03104_),
    .I1(_03380_),
    .S(_03163_),
    .Z(_03381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18055_ (.I0(_03135_),
    .I1(_03109_),
    .S(_03163_),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18056_ (.I0(_03381_),
    .I1(_03382_),
    .S(_03248_),
    .Z(_03383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18057_ (.A1(_03127_),
    .A2(_03383_),
    .Z(_03384_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18058_ (.A1(_03100_),
    .A2(_03281_),
    .A3(_03384_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_319_clk_i_regs (.I(clknet_6_10__leaf_clk_i_regs),
    .Z(clknet_leaf_319_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_320_clk_i_regs (.I(clknet_6_11__leaf_clk_i_regs),
    .Z(clknet_leaf_320_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18061_ (.A1(_11484_[0]),
    .A2(_03187_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18062_ (.A1(_11483_[0]),
    .A2(_03181_),
    .B1(_03190_),
    .B2(net152),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18063_ (.A1(_11487_[0]),
    .A2(_03183_),
    .B(_03388_),
    .C(_03389_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18064_ (.I(_11252_[0]),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18065_ (.A1(net3157),
    .A2(net3130),
    .B(net3159),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18066_ (.I(_11251_[0]),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18067_ (.A1(net3155),
    .A2(_03392_),
    .B(net3154),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _18068_ (.A1(net3152),
    .A2(_03394_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18069_ (.I0(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .I1(_03395_),
    .S(_03152_),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18070_ (.A1(net3647),
    .A2(_03396_),
    .Z(_03397_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18071_ (.A1(net3371),
    .A2(_03397_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18072_ (.A1(_07282_),
    .A2(_02906_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18073_ (.A1(_03298_),
    .A2(_03390_),
    .B1(_03398_),
    .B2(_03399_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18074_ (.A1(_09064_),
    .A2(net3190),
    .A3(_03385_),
    .A4(_03400_),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18075_ (.I0(net29),
    .I1(\load_store_unit_i.rdata_q[11] ),
    .I2(\load_store_unit_i.rdata_q[19] ),
    .I3(net52),
    .S0(net3471),
    .S1(net3470),
    .Z(_03402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18076_ (.I0(net46),
    .I1(net52),
    .S(net3471),
    .Z(_03403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18077_ (.I0(net29),
    .I1(net37),
    .S(net3471),
    .Z(_03404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18078_ (.I0(_03403_),
    .I1(_03404_),
    .S(_03076_),
    .Z(_03405_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18079_ (.A1(net3400),
    .A2(_03402_),
    .B1(_03405_),
    .B2(\load_store_unit_i.data_type_q[2] ),
    .C(_03243_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18080_ (.A1(_03379_),
    .A2(_03401_),
    .B(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_322_clk_i_regs (.I(clknet_6_14__leaf_clk_i_regs),
    .Z(clknet_leaf_322_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18082_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .I1(net3093),
    .S(_03232_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18083_ (.I0(net47),
    .I1(net53),
    .S(net3471),
    .Z(_03409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18084_ (.I0(net30),
    .I1(net39),
    .S(net3471),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18085_ (.I0(_03409_),
    .I1(_03410_),
    .S(_03076_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18086_ (.I0(net30),
    .I1(\load_store_unit_i.rdata_q[12] ),
    .I2(\load_store_unit_i.rdata_q[20] ),
    .I3(net53),
    .S0(net3471),
    .S1(net3470),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18087_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_03411_),
    .B1(_03412_),
    .B2(_03079_),
    .C(_03086_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18088_ (.A1(_03338_),
    .A2(_03391_),
    .B(_03393_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18089_ (.A1(net3152),
    .A2(_03414_),
    .B(net3153),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18090_ (.A1(net3150),
    .A2(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18091_ (.I0(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .I1(_03416_),
    .S(_03152_),
    .Z(_03417_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18092_ (.A1(net3417),
    .A2(_03417_),
    .Z(_03418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18093_ (.A1(net3647),
    .A2(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .B(_03418_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18094_ (.A1(net3374),
    .A2(_03419_),
    .B(_08265_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18095_ (.A1(_11491_[0]),
    .A2(_03183_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18096_ (.A1(_11495_[0]),
    .A2(net3206),
    .B(_03420_),
    .C(_03421_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18097_ (.A1(net153),
    .A2(_03190_),
    .B1(_03187_),
    .B2(_11492_[0]),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18098_ (.A1(_03093_),
    .A2(_03163_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18099_ (.I0(_03135_),
    .I1(_03109_),
    .S(_03424_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18100_ (.I0(_11518_[0]),
    .I1(_11526_[0]),
    .S(_03114_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18101_ (.I0(_03426_),
    .I1(_03256_),
    .I2(_03257_),
    .I3(_03322_),
    .S0(net3207),
    .S1(net3253),
    .Z(_03427_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18102_ (.A1(_03273_),
    .A2(_03138_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18103_ (.A1(net3207),
    .A2(_03144_),
    .B(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18104_ (.I0(_03427_),
    .I1(_03429_),
    .S(_03111_),
    .Z(_03430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18105_ (.A1(_03248_),
    .A2(_03381_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18106_ (.A1(_03248_),
    .A2(_03430_),
    .B(_03431_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18107_ (.I0(_03425_),
    .I1(_03432_),
    .S(_03127_),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18108_ (.A1(_03091_),
    .A2(_03433_),
    .Z(_03434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18109_ (.I0(_03171_),
    .I1(_03370_),
    .S(_03163_),
    .Z(_03435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18110_ (.I0(_03435_),
    .I1(_03376_),
    .S(_03248_),
    .Z(_03436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18111_ (.I0(_03159_),
    .I1(_03436_),
    .S(_03127_),
    .Z(_03437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18112_ (.A1(_03114_),
    .A2(_03437_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18113_ (.A1(_03422_),
    .A2(_03423_),
    .A3(_03434_),
    .A4(_03438_),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_324_clk_i_regs (.I(clknet_6_14__leaf_clk_i_regs),
    .Z(clknet_leaf_324_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _18115_ (.A1(_08265_),
    .A2(_09094_),
    .B1(_03298_),
    .B2(_03420_),
    .C(net3190),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _18116_ (.A1(_03218_),
    .A2(_03413_),
    .B1(_03439_),
    .B2(_03441_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3094 (.I(_08254_),
    .Z(net3094));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18118_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .I1(_03442_),
    .S(_03232_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18119_ (.I0(_03261_),
    .I1(_03263_),
    .I2(_03255_),
    .I3(_03258_),
    .S0(net3207),
    .S1(_03163_),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _18120_ (.I0(_03159_),
    .I1(_03351_),
    .I2(_03353_),
    .I3(_03444_),
    .S0(_03093_),
    .S1(_03127_),
    .Z(_03445_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18121_ (.A1(_03245_),
    .A2(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18122_ (.I0(_03319_),
    .I1(_03331_),
    .S(_03248_),
    .Z(_03447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18123_ (.A1(_03127_),
    .A2(_03447_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_325_clk_i_regs (.I(clknet_6_14__leaf_clk_i_regs),
    .Z(clknet_leaf_325_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18125_ (.A1(_11503_[0]),
    .A2(net3206),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18126_ (.A1(_11499_[0]),
    .A2(_03183_),
    .B(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18127_ (.A1(net154),
    .A2(_03190_),
    .B1(_03187_),
    .B2(_11500_[0]),
    .C(_03451_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18128_ (.A1(_11245_[0]),
    .A2(_03309_),
    .B(_11251_[0]),
    .C(_11244_[0]),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18129_ (.A1(_11252_[0]),
    .A2(_11251_[0]),
    .B(_11256_[0]),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18130_ (.I(net3153),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18131_ (.A1(net3111),
    .A2(net3129),
    .B(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18132_ (.A1(net3150),
    .A2(_03456_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18133_ (.A1(net3151),
    .A2(_03457_),
    .Z(_03458_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _18134_ (.A1(net3124),
    .A2(_03458_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18135_ (.I0(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .I1(_03459_),
    .S(_03154_),
    .Z(_03460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18136_ (.A1(net3371),
    .A2(_03460_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18137_ (.A1(_03199_),
    .A2(_03452_),
    .B(_03461_),
    .C(_09115_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18138_ (.A1(_03214_),
    .A2(_03216_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18139_ (.A1(_03463_),
    .A2(_03217_),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18140_ (.A1(_03347_),
    .A2(_03448_),
    .B(_03462_),
    .C(_03464_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18141_ (.I0(net31),
    .I1(\load_store_unit_i.rdata_q[13] ),
    .I2(\load_store_unit_i.rdata_q[21] ),
    .I3(net54),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(net3470),
    .Z(_03466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18142_ (.I0(net48),
    .I1(net54),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18143_ (.I0(net31),
    .I1(net40),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18144_ (.I0(_03467_),
    .I1(_03468_),
    .S(_03076_),
    .Z(_03469_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18145_ (.A1(net3400),
    .A2(_03466_),
    .B1(_03469_),
    .B2(\load_store_unit_i.data_type_q[2] ),
    .C(_03243_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18146_ (.A1(_03446_),
    .A2(_03465_),
    .B(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_330_clk_i_regs (.I(clknet_6_11__leaf_clk_i_regs),
    .Z(clknet_leaf_330_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18148_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .I1(net3088),
    .S(_03232_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18149_ (.I0(_03318_),
    .I1(_03321_),
    .S(_03163_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18150_ (.I0(_03291_),
    .I1(_03473_),
    .S(_03093_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18151_ (.A1(_03248_),
    .A2(_03165_),
    .A3(_03106_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18152_ (.A1(_03093_),
    .A2(_03292_),
    .B(_03135_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18153_ (.A1(_03127_),
    .A2(_03475_),
    .A3(_03476_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18154_ (.A1(_03127_),
    .A2(_03474_),
    .B(_03477_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18155_ (.A1(_03245_),
    .A2(_03478_),
    .Z(_03479_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18156_ (.A1(net364),
    .A2(_03190_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18157_ (.A1(_03131_),
    .A2(_03248_),
    .A3(_03267_),
    .Z(_03481_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18158_ (.A1(_03131_),
    .A2(_03093_),
    .A3(_03275_),
    .A4(_03279_),
    .Z(_03482_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18159_ (.A1(_03481_),
    .A2(_03482_),
    .Z(_03483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18160_ (.A1(_11511_[0]),
    .A2(net3206),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18161_ (.A1(_11507_[0]),
    .A2(_03183_),
    .B(_03484_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18162_ (.A1(_11508_[0]),
    .A2(_03187_),
    .B1(_03347_),
    .B2(_03483_),
    .C(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18163_ (.A1(_03480_),
    .A2(_03486_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18164_ (.A1(_03479_),
    .A2(_03487_),
    .B(_03298_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_327_clk_i_regs (.I(clknet_6_14__leaf_clk_i_regs),
    .Z(clknet_leaf_327_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18166_ (.A1(net3150),
    .A2(net3151),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18167_ (.A1(net3124),
    .A2(_03490_),
    .B(net3125),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18168_ (.A1(net3153),
    .A2(net3151),
    .A3(net3125),
    .Z(_03492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18169_ (.A1(net3152),
    .A2(_03414_),
    .B(_03492_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18170_ (.A1(_03491_),
    .A2(_03493_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18171_ (.A1(net3122),
    .A2(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_332_clk_i_regs (.I(clknet_6_11__leaf_clk_i_regs),
    .Z(clknet_leaf_332_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18173_ (.I0(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .I1(_03495_),
    .S(_03152_),
    .Z(_03497_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18174_ (.A1(net3647),
    .A2(_03497_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18175_ (.A1(net3417),
    .A2(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .B(net3371),
    .C(_03498_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _18176_ (.A1(_09129_),
    .A2(net3190),
    .A3(_03499_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18177_ (.I0(net32),
    .I1(\load_store_unit_i.rdata_q[14] ),
    .I2(\load_store_unit_i.rdata_q[22] ),
    .I3(net55),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(net3470),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18178_ (.I0(net50),
    .I1(net55),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18179_ (.I0(net32),
    .I1(net41),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18180_ (.I0(_03502_),
    .I1(_03503_),
    .S(_03076_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18181_ (.A1(net3400),
    .A2(_03501_),
    .B1(_03504_),
    .B2(\load_store_unit_i.data_type_q[2] ),
    .C(_03243_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18182_ (.A1(_03488_),
    .A2(_03500_),
    .B(_03505_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_331_clk_i_regs (.I(clknet_6_11__leaf_clk_i_regs),
    .Z(clknet_leaf_331_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18184_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .I1(net3082),
    .S(net3185),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18185_ (.A1(_11519_[0]),
    .A2(net3206),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18186_ (.A1(_11515_[0]),
    .A2(_03183_),
    .B(_03508_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18187_ (.A1(net156),
    .A2(_03190_),
    .B1(_03187_),
    .B2(_11516_[0]),
    .C(_03509_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18188_ (.A1(_03199_),
    .A2(_03510_),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18189_ (.A1(net3647),
    .A2(net3371),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18190_ (.A1(_11279_[0]),
    .A2(_11273_[0]),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18191_ (.A1(net3149),
    .A2(net3118),
    .A3(net3109),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18192_ (.I(net3120),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18193_ (.A1(net3123),
    .A2(_11264_[0]),
    .B(_11272_[0]),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18194_ (.I(_11278_[0]),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18195_ (.A1(_03515_),
    .A2(_03516_),
    .B(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18196_ (.A1(_11265_[0]),
    .A2(_11288_[0]),
    .A3(_11255_[0]),
    .A4(_03513_),
    .Z(_03519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18197_ (.A1(net3117),
    .A2(_03518_),
    .B(_03519_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18198_ (.A1(_03453_),
    .A2(_03454_),
    .A3(_03514_),
    .B(_03520_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18199_ (.A1(_03457_),
    .A2(net3110),
    .B(net3103),
    .C(net3118),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18200_ (.A1(net3100),
    .A2(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18201_ (.I0(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .I1(_03523_),
    .S(_03152_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18202_ (.A1(net3647),
    .A2(_03524_),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18203_ (.A1(net3371),
    .A2(_03525_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18204_ (.A1(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .A2(_03512_),
    .B(_03526_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18205_ (.A1(_09147_),
    .A2(net3190),
    .A3(_03511_),
    .A4(_03527_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18206_ (.I0(_03370_),
    .I1(_03371_),
    .S(_03163_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _18207_ (.I0(_03159_),
    .I1(_03166_),
    .I2(_03175_),
    .I3(_03529_),
    .S0(_03093_),
    .S1(_03127_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18208_ (.I0(_03113_),
    .I1(_03147_),
    .S(_03093_),
    .Z(_03531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18209_ (.A1(_03127_),
    .A2(_03531_),
    .B(_03281_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18210_ (.A1(_03245_),
    .A2(_03530_),
    .B1(_03532_),
    .B2(_03114_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18211_ (.I0(net33),
    .I1(\load_store_unit_i.rdata_q[15] ),
    .I2(\load_store_unit_i.rdata_q[23] ),
    .I3(net56),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18212_ (.I0(net51),
    .I1(net56),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18213_ (.I0(net33),
    .I1(net42),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18214_ (.I0(_03535_),
    .I1(_03536_),
    .S(_03076_),
    .Z(_03537_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18215_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_03537_),
    .Z(_03538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18216_ (.A1(net3400),
    .A2(_03534_),
    .B(_03538_),
    .C(_03243_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18217_ (.A1(_03528_),
    .A2(_03533_),
    .B(_03539_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_334_clk_i_regs (.I(clknet_6_11__leaf_clk_i_regs),
    .Z(clknet_leaf_334_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18219_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .I1(net3081),
    .S(net3185),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18220_ (.A1(_11527_[0]),
    .A2(net3206),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18221_ (.A1(_11523_[0]),
    .A2(_03183_),
    .B(_03542_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18222_ (.A1(net402),
    .A2(_03190_),
    .B1(_03187_),
    .B2(_11524_[0]),
    .C(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _18223_ (.A1(net3657),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A3(_08471_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_335_clk_i_regs (.I(clknet_6_11__leaf_clk_i_regs),
    .Z(clknet_leaf_335_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18225_ (.A1(_11184_[0]),
    .A2(_03545_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18226_ (.A1(net3108),
    .A2(_03494_),
    .B(_03517_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18227_ (.A1(net3117),
    .A2(_03548_),
    .B(net3119),
    .C(net3115),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18228_ (.A1(net3121),
    .A2(net3117),
    .A3(net560),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18229_ (.A1(net3117),
    .A2(net3115),
    .A3(_11278_[0]),
    .Z(_03551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18230_ (.A1(net3115),
    .A2(net3119),
    .B(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18231_ (.A1(_03493_),
    .A2(_03491_),
    .A3(_03550_),
    .B(_03552_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _18232_ (.A1(_03545_),
    .A2(_03549_),
    .A3(net3099),
    .Z(_03554_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18233_ (.A1(_03547_),
    .A2(_03554_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18234_ (.A1(net3417),
    .A2(_03555_),
    .B(net3374),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18235_ (.A1(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .A2(_03512_),
    .B(_03556_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18236_ (.A1(_03199_),
    .A2(_03544_),
    .B(_03557_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18237_ (.A1(_09173_),
    .A2(_03464_),
    .A3(_03558_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18238_ (.A1(_03114_),
    .A2(_03530_),
    .B1(_03532_),
    .B2(_03245_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_338_clk_i_regs (.I(clknet_6_11__leaf_clk_i_regs),
    .Z(clknet_leaf_338_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18240_ (.I0(net34),
    .I1(net27),
    .I2(\load_store_unit_i.rdata_q[16] ),
    .I3(net57),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(net3471),
    .Z(_03562_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18241_ (.A1(\load_store_unit_i.data_sign_ext_q ),
    .A2(_03538_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _18242_ (.A1(_03218_),
    .A2(_03086_),
    .A3(_03563_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_339_clk_i_regs (.I(clknet_6_10__leaf_clk_i_regs),
    .Z(clknet_leaf_339_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18244_ (.A1(net3400),
    .A2(_03562_),
    .B(_03564_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18245_ (.A1(_03559_),
    .A2(_03560_),
    .B(_03566_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_342_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_342_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3093 (.I(_03407_),
    .Z(net3093));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18248_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .I1(net3056),
    .S(_03232_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18249_ (.I0(net35),
    .I1(net38),
    .I2(\load_store_unit_i.rdata_q[17] ),
    .I3(net58),
    .S0(net3470),
    .S1(net3471),
    .Z(_03570_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18250_ (.A1(_03079_),
    .A2(_03570_),
    .B(_03564_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18251_ (.A1(_03114_),
    .A2(_03478_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18252_ (.A1(_03137_),
    .A2(_03245_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18253_ (.A1(_03483_),
    .A2(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18254_ (.A1(net3119),
    .A2(net3100),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18255_ (.A1(net477),
    .A2(_03575_),
    .B(net3116),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18256_ (.A1(net3113),
    .A2(_03576_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18257_ (.I0(_11187_[0]),
    .I1(_03577_),
    .S(_03152_),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18258_ (.A1(net3647),
    .A2(_03578_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18259_ (.A1(net3371),
    .A2(_03579_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18260_ (.A1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .A2(_03512_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18261_ (.I(_11531_[0]),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18262_ (.A1(_03582_),
    .A2(_03180_),
    .B1(_03187_),
    .B2(_11532_[0]),
    .C1(_11535_[0]),
    .C2(net3206),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18263_ (.A1(net158),
    .A2(_03190_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18264_ (.A1(_03583_),
    .A2(_03584_),
    .B(_03199_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18265_ (.A1(_03580_),
    .A2(_03581_),
    .B(_03585_),
    .C(_09193_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18266_ (.A1(_03218_),
    .A2(_03572_),
    .A3(_03574_),
    .A4(_03586_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18267_ (.A1(_03587_),
    .A2(_03571_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_343_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_343_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18269_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .I1(_03588_),
    .S(net3185),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18270_ (.I0(_11457_[0]),
    .I1(_11465_[0]),
    .I2(_11582_[0]),
    .I3(_11574_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18271_ (.I0(_03324_),
    .I1(_03590_),
    .S(net3207),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18272_ (.I0(net3252),
    .I1(_11433_[0]),
    .I2(_11614_[0]),
    .I3(_11606_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18273_ (.I0(_11441_[0]),
    .I1(_11449_[0]),
    .I2(_11598_[0]),
    .I3(_11590_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18274_ (.I0(_03592_),
    .I1(_03593_),
    .S(_03273_),
    .Z(_03594_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18275_ (.I0(_03591_),
    .I1(_03429_),
    .I2(_03594_),
    .I3(_03427_),
    .S0(_03248_),
    .S1(_03163_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18276_ (.I(_03595_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18277_ (.I0(_03383_),
    .I1(_03596_),
    .S(_03127_),
    .Z(_03597_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18278_ (.A1(_03091_),
    .A2(_03597_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18279_ (.I(_03376_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18280_ (.A1(_03127_),
    .A2(_03093_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18281_ (.I0(_03135_),
    .I1(_03599_),
    .S(_03600_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18282_ (.A1(_11431_[0]),
    .A2(_03183_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18283_ (.A1(_11427_[0]),
    .A2(_03181_),
    .B1(_03187_),
    .B2(_11428_[0]),
    .C(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18284_ (.A1(net175),
    .A2(_03190_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18285_ (.A1(_03100_),
    .A2(_03601_),
    .B(_03603_),
    .C(_03604_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18286_ (.I0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .I1(_11201_[0]),
    .S(_03154_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18287_ (.A1(_03298_),
    .A2(_03605_),
    .B1(_03606_),
    .B2(net3370),
    .C(_09507_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18288_ (.A1(_03598_),
    .A2(_03607_),
    .Z(_03608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _18289_ (.I(net3471),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18290_ (.A1(net3470),
    .A2(_03609_),
    .A3(net39),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18291_ (.A1(_03076_),
    .A2(net3471),
    .A3(net30),
    .Z(_03611_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18292_ (.A1(_03610_),
    .A2(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18293_ (.A1(_03076_),
    .A2(net3471),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18294_ (.A1(net3470),
    .A2(_03609_),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18295_ (.A1(\load_store_unit_i.rdata_q[4] ),
    .A2(_03613_),
    .B1(_03614_),
    .B2(\load_store_unit_i.rdata_q[12] ),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18296_ (.I0(_03612_),
    .I1(_03615_),
    .S(_03079_),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18297_ (.I(\load_store_unit_i.data_type_q[2] ),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18298_ (.A1(_03617_),
    .A2(\load_store_unit_i.data_type_q[1] ),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18299_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net47),
    .B1(_03618_),
    .B2(\load_store_unit_i.rdata_q[20] ),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _18300_ (.A1(net3470),
    .A2(net3471),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18301_ (.A1(_03619_),
    .A2(_03620_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_347_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_347_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18303_ (.A1(_03076_),
    .A2(_03609_),
    .A3(net53),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18304_ (.A1(_03228_),
    .A2(_03616_),
    .A3(_03621_),
    .A4(_03623_),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18305_ (.A1(_03218_),
    .A2(_03608_),
    .B(_03624_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_348_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_348_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18307_ (.A1(_03224_),
    .A2(_03228_),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18308_ (.A1(_03223_),
    .A2(_03627_),
    .Z(_03628_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18309_ (.A1(_06740_),
    .A2(_03628_),
    .Z(_03629_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_349_clk_i_regs (.I(clknet_6_10__leaf_clk_i_regs),
    .Z(clknet_leaf_349_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18311_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .I1(_03625_),
    .S(_03629_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18312_ (.A1(_11539_[0]),
    .A2(_03183_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18313_ (.A1(_11543_[0]),
    .A2(net3206),
    .B1(_03187_),
    .B2(_11540_[0]),
    .C(_03631_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18314_ (.A1(net361),
    .A2(_03190_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18315_ (.A1(_03632_),
    .A2(_03633_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18316_ (.A1(_03114_),
    .A2(_03445_),
    .B1(_03634_),
    .B2(_03298_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18317_ (.I(_09209_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18318_ (.A1(_03448_),
    .A2(_03573_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18319_ (.A1(net3116),
    .A2(net3099),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18320_ (.A1(net3113),
    .A2(_03638_),
    .B(net3114),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18321_ (.A1(net3112),
    .A2(_03639_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18322_ (.I0(_11189_[0]),
    .I1(_03640_),
    .S(_03152_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18323_ (.A1(net3647),
    .A2(_03641_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18324_ (.A1(net3417),
    .A2(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .B(net3371),
    .C(_03642_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18325_ (.A1(_03636_),
    .A2(net3190),
    .A3(_03637_),
    .A4(_03643_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18326_ (.I0(net36),
    .I1(net49),
    .I2(\load_store_unit_i.rdata_q[18] ),
    .I3(net28),
    .S0(net3470),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03645_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18327_ (.A1(net3400),
    .A2(_03645_),
    .B(_03564_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18328_ (.A1(_03635_),
    .A2(_03644_),
    .B(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_350_clk_i_regs (.I(clknet_6_10__leaf_clk_i_regs),
    .Z(clknet_leaf_350_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18330_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .I1(net3067),
    .S(_03232_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18331_ (.I0(net37),
    .I1(net52),
    .I2(\load_store_unit_i.rdata_q[19] ),
    .I3(net29),
    .S0(net3470),
    .S1(net3471),
    .Z(_03649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18332_ (.A1(_03079_),
    .A2(_03649_),
    .B(_03564_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18333_ (.A1(_03100_),
    .A2(_03433_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18334_ (.A1(_03245_),
    .A2(_03437_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18335_ (.A1(_11551_[0]),
    .A2(net3206),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18336_ (.A1(_11547_[0]),
    .A2(_03183_),
    .B(_03653_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18337_ (.A1(net160),
    .A2(_03190_),
    .B1(_03187_),
    .B2(_11548_[0]),
    .C(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18338_ (.A1(_03199_),
    .A2(_03655_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18339_ (.I(_11300_[0]),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18340_ (.A1(_11287_[0]),
    .A2(_11289_[0]),
    .A3(_11294_[0]),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18341_ (.A1(_11290_[0]),
    .A2(_11289_[0]),
    .A3(_11294_[0]),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18342_ (.A1(_11295_[0]),
    .A2(_11294_[0]),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18343_ (.A1(_03659_),
    .A2(_03660_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18344_ (.A1(net3100),
    .A2(net3107),
    .B(net3102),
    .C(net3112),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18345_ (.A1(_03657_),
    .A2(_03662_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18346_ (.A1(net3148),
    .A2(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18347_ (.I0(_11197_[0]),
    .I1(_03664_),
    .S(_03152_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18348_ (.A1(net3647),
    .A2(_03665_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18349_ (.A1(net3417),
    .A2(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .B(net3371),
    .C(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18350_ (.A1(_09227_),
    .A2(net3190),
    .A3(_03656_),
    .A4(_03667_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _18351_ (.A1(_03651_),
    .A2(_03652_),
    .A3(_03668_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18352_ (.A1(_03650_),
    .A2(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_352_clk_i_regs (.I(clknet_6_11__leaf_clk_i_regs),
    .Z(clknet_leaf_352_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18354_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .I1(net3066),
    .S(_03232_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18355_ (.I0(net39),
    .I1(net53),
    .I2(\load_store_unit_i.rdata_q[20] ),
    .I3(net30),
    .S0(net3470),
    .S1(net3471),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18356_ (.A1(_03079_),
    .A2(_03672_),
    .B(_03564_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18357_ (.I(_09261_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18358_ (.A1(_03137_),
    .A2(_03245_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18359_ (.A1(_03114_),
    .A2(_03282_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18360_ (.A1(_11559_[0]),
    .A2(net3206),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18361_ (.A1(_11555_[0]),
    .A2(_03183_),
    .B(_03677_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18362_ (.A1(net161),
    .A2(_03190_),
    .B1(_03187_),
    .B2(_11556_[0]),
    .C(_03678_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18363_ (.A1(_03384_),
    .A2(_03675_),
    .B1(_03676_),
    .B2(_03378_),
    .C(_03679_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18364_ (.A1(_03298_),
    .A2(_03680_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18365_ (.I(_11306_[0]),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _18366_ (.A1(net3116),
    .A2(net3114),
    .A3(_11300_[0]),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18367_ (.A1(_11300_[0]),
    .A2(_03660_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18368_ (.A1(net3112),
    .A2(_11300_[0]),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18369_ (.A1(_03684_),
    .A2(_03685_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18370_ (.A1(net3099),
    .A2(_03683_),
    .B(net3101),
    .C(net3148),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18371_ (.A1(_03682_),
    .A2(_03687_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18372_ (.A1(net3146),
    .A2(_03688_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18373_ (.I0(_11201_[0]),
    .I1(_03689_),
    .S(_03152_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18374_ (.A1(net3647),
    .A2(_03690_),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18375_ (.A1(net3417),
    .A2(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .B(net3371),
    .C(_03691_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18376_ (.A1(_03674_),
    .A2(net3190),
    .A3(_03681_),
    .A4(_03692_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18377_ (.A1(_03673_),
    .A2(_03693_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_356_clk_i_regs (.I(clknet_6_9__leaf_clk_i_regs),
    .Z(clknet_leaf_356_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18379_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .I1(net3065),
    .S(_03232_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18380_ (.I(_11210_[0]),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18381_ (.I(net3147),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18382_ (.A1(_11301_[0]),
    .A2(_11307_[0]),
    .A3(_11313_[0]),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18383_ (.A1(_03658_),
    .A2(_03521_),
    .B(_03661_),
    .C(_03698_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18384_ (.A1(net3146),
    .A2(_11306_[0]),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18385_ (.A1(net3148),
    .A2(net3146),
    .A3(_11300_[0]),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _18386_ (.A1(_03697_),
    .A2(net3098),
    .A3(net3128),
    .A4(net3106),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18387_ (.A1(net3144),
    .A2(_03702_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18388_ (.I0(_03696_),
    .I1(_03703_),
    .S(_03152_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18389_ (.A1(net3417),
    .A2(_03704_),
    .B(net3375),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _18390_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(_03512_),
    .B(_03705_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18391_ (.A1(net3374),
    .A2(_03190_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18392_ (.I(_11563_[0]),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18393_ (.A1(_03708_),
    .A2(_03180_),
    .B1(_03187_),
    .B2(_11564_[0]),
    .C1(_11567_[0]),
    .C2(net3206),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18394_ (.A1(_03199_),
    .A2(_03709_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18395_ (.A1(net162),
    .A2(_03707_),
    .B(_03710_),
    .C(_09276_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18396_ (.A1(_03333_),
    .A2(_03676_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18397_ (.A1(_03355_),
    .A2(_03573_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18398_ (.A1(net3190),
    .A2(_03711_),
    .A3(_03712_),
    .A4(_03713_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18399_ (.I0(net40),
    .I1(net54),
    .I2(\load_store_unit_i.rdata_q[21] ),
    .I3(net31),
    .S0(net3470),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18400_ (.A1(net3400),
    .A2(_03715_),
    .B(_03564_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18401_ (.A1(_03706_),
    .A2(_03714_),
    .B(_03716_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_359_clk_i_regs (.I(clknet_6_9__leaf_clk_i_regs),
    .Z(clknet_leaf_359_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18403_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .I1(net3080),
    .S(_03232_),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18404_ (.I(_09292_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18405_ (.I(_11571_[0]),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18406_ (.A1(_03720_),
    .A2(_03180_),
    .B1(_03187_),
    .B2(_11572_[0]),
    .C1(_11575_[0]),
    .C2(net3206),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18407_ (.A1(net163),
    .A2(_03190_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18408_ (.A1(_03721_),
    .A2(_03722_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18409_ (.A1(_03245_),
    .A2(_03296_),
    .B1(_03723_),
    .B2(_03298_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18410_ (.A1(_03114_),
    .A2(_03284_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18411_ (.A1(_03719_),
    .A2(net3190),
    .A3(_03724_),
    .A4(_03725_),
    .Z(_03726_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18412_ (.I(net3145),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18413_ (.A1(net3148),
    .A2(net3146),
    .A3(_11319_[0]),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18414_ (.A1(_03553_),
    .A2(_03683_),
    .B(_03686_),
    .C(_03728_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18415_ (.A1(net3143),
    .A2(net3147),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18416_ (.A1(net3146),
    .A2(net3143),
    .A3(_11306_[0]),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18417_ (.A1(_03727_),
    .A2(_03729_),
    .A3(_03730_),
    .A4(_03731_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18418_ (.A1(net3141),
    .A2(_03732_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18419_ (.I0(_11221_[0]),
    .I1(_03733_),
    .S(_03152_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18420_ (.A1(net3647),
    .A2(_03734_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _18421_ (.A1(net3417),
    .A2(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .B(net3371),
    .C(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18422_ (.I0(net41),
    .I1(net55),
    .I2(\load_store_unit_i.rdata_q[22] ),
    .I3(net32),
    .S0(net3470),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18423_ (.A1(net3400),
    .A2(_03737_),
    .B(_03564_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18424_ (.A1(_03726_),
    .A2(_03736_),
    .B(_03738_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_360_clk_i_regs (.I(clknet_6_9__leaf_clk_i_regs),
    .Z(clknet_leaf_360_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18426_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .I1(net3076),
    .S(_03232_),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18427_ (.I0(net42),
    .I1(net56),
    .I2(\load_store_unit_i.rdata_q[23] ),
    .I3(net33),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18428_ (.A1(net3400),
    .A2(_03741_),
    .B(_03564_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18429_ (.I(_09309_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18430_ (.A1(_11312_[0]),
    .A2(_11318_[0]),
    .A3(_11324_[0]),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18431_ (.A1(_03699_),
    .A2(_03700_),
    .A3(_03701_),
    .A4(_03744_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18432_ (.A1(_11325_[0]),
    .A2(_11324_[0]),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _18433_ (.A1(net3143),
    .A2(_11318_[0]),
    .A3(_11324_[0]),
    .B(_03746_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18434_ (.A1(net3096),
    .A2(net3105),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18435_ (.A1(net585),
    .A2(net3139),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18436_ (.I0(_09860_[0]),
    .I1(_03749_),
    .S(_03152_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18437_ (.I0(_07862_),
    .I1(_03750_),
    .S(net3417),
    .Z(_03751_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18438_ (.A1(_03751_),
    .A2(net3374),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18439_ (.A1(_03177_),
    .A2(_03245_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18440_ (.A1(_11583_[0]),
    .A2(net3206),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18441_ (.A1(_11579_[0]),
    .A2(_03183_),
    .B(_03754_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18442_ (.A1(net373),
    .A2(_03190_),
    .B1(_03187_),
    .B2(_11580_[0]),
    .C(_03755_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18443_ (.A1(_03100_),
    .A2(_03130_),
    .A3(_03149_),
    .B(_03756_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18444_ (.A1(_03753_),
    .A2(_03757_),
    .B(_03298_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18445_ (.A1(_03752_),
    .A2(net3190),
    .A3(_03743_),
    .A4(_03758_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18446_ (.A1(_03759_),
    .A2(_03742_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_361_clk_i_regs (.I(clknet_6_9__leaf_clk_i_regs),
    .Z(clknet_leaf_361_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18448_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .I1(net737),
    .S(net3185),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18449_ (.I0(_03074_),
    .I1(_03075_),
    .S(\load_store_unit_i.rdata_offset_q[1] ),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18450_ (.A1(_03079_),
    .A2(_03762_),
    .B(_03564_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18451_ (.A1(net3145),
    .A2(net3142),
    .A3(net3140),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18452_ (.A1(_03729_),
    .A2(_03730_),
    .A3(_03731_),
    .A4(_03764_),
    .Z(_03765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18453_ (.A1(net3139),
    .A2(net3127),
    .B(net3140),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18454_ (.A1(_03765_),
    .A2(_03766_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18455_ (.A1(net3137),
    .A2(_03767_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18456_ (.I0(_03151_),
    .I1(_03768_),
    .S(_03152_),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18457_ (.I0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .I1(_03769_),
    .S(net3417),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18458_ (.I0(_11449_[0]),
    .I1(_11457_[0]),
    .I2(_11590_[0]),
    .I3(_11582_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18459_ (.I0(_03252_),
    .I1(_03771_),
    .S(net3207),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18460_ (.I0(_03372_),
    .I1(_03772_),
    .S(_03163_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18461_ (.I0(_03529_),
    .I1(_03773_),
    .S(_03093_),
    .Z(_03774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18462_ (.I0(_03176_),
    .I1(_03774_),
    .S(_03127_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18463_ (.A1(_03159_),
    .A2(_03248_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18464_ (.A1(_03131_),
    .A2(_03776_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18465_ (.A1(_03248_),
    .A2(_03113_),
    .B(_03777_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18466_ (.A1(_11591_[0]),
    .A2(net3206),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18467_ (.A1(_11587_[0]),
    .A2(_03183_),
    .B(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18468_ (.A1(_11588_[0]),
    .A2(_03187_),
    .B1(_03573_),
    .B2(_03778_),
    .C(_03780_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18469_ (.A1(net376),
    .A2(_03707_),
    .B(_09329_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18470_ (.A1(_03199_),
    .A2(_03781_),
    .B(_03782_),
    .C(net3190),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _18471_ (.A1(net3370),
    .A2(_03770_),
    .B1(_03775_),
    .B2(_03114_),
    .C(_03783_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18472_ (.A1(_03763_),
    .A2(_03784_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_364_clk_i_regs (.I(clknet_6_6__leaf_clk_i_regs),
    .Z(clknet_leaf_364_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18474_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .I1(net3063),
    .S(_03232_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18475_ (.A1(_06718_),
    .A2(_03218_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18476_ (.I0(_03239_),
    .I1(_03240_),
    .S(net3470),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18477_ (.A1(net3400),
    .A2(_03788_),
    .B(_03564_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18478_ (.A1(_09346_),
    .A2(_03787_),
    .B(_03789_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18479_ (.I(_03310_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18480_ (.I(net3138),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18481_ (.A1(net3139),
    .A2(_03748_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18482_ (.A1(net3140),
    .A2(_03793_),
    .B(net3137),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18483_ (.A1(_03794_),
    .A2(_03792_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18484_ (.A1(_03795_),
    .A2(net3135),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18485_ (.I0(_03791_),
    .I1(_03796_),
    .S(_03152_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18486_ (.I0(_07960_),
    .I1(_03797_),
    .S(net3417),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18487_ (.A1(net3375),
    .A2(_03798_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18488_ (.I0(_03159_),
    .I1(_03280_),
    .S(_03600_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18489_ (.I(_11595_[0]),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18490_ (.A1(_03801_),
    .A2(_03180_),
    .B1(_03187_),
    .B2(_11596_[0]),
    .C1(_11599_[0]),
    .C2(net3206),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18491_ (.A1(_03199_),
    .A2(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18492_ (.A1(net289),
    .A2(_03707_),
    .B1(_03800_),
    .B2(_03245_),
    .C(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18493_ (.A1(_03273_),
    .A2(_03590_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18494_ (.A1(net3207),
    .A2(_03593_),
    .B(_03805_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18495_ (.I0(_03326_),
    .I1(_03806_),
    .S(_03163_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18496_ (.I0(_03473_),
    .I1(_03807_),
    .S(_03093_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18497_ (.I0(_03294_),
    .I1(_03808_),
    .S(_03127_),
    .Z(_03809_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18498_ (.A1(_03100_),
    .A2(_03809_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18499_ (.A1(_08265_),
    .A2(_03218_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _18500_ (.A1(_03799_),
    .A2(_03804_),
    .A3(_03810_),
    .A4(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18501_ (.A1(_03790_),
    .A2(_03812_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_365_clk_i_regs (.I(clknet_6_9__leaf_clk_i_regs),
    .Z(clknet_leaf_365_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18503_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .I1(net584),
    .S(_03232_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18504_ (.A1(_03248_),
    .A2(_03331_),
    .B(_03777_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18505_ (.A1(_11604_[0]),
    .A2(_03187_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18506_ (.A1(_11607_[0]),
    .A2(net3206),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18507_ (.A1(_11603_[0]),
    .A2(_03183_),
    .B(_03816_),
    .C(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18508_ (.A1(net167),
    .A2(_03190_),
    .B1(_03573_),
    .B2(_03815_),
    .C(_03818_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18509_ (.I0(_11433_[0]),
    .I1(_11441_[0]),
    .I2(_11606_[0]),
    .I3(_11598_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18510_ (.I0(_03771_),
    .I1(_03820_),
    .S(net3207),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18511_ (.I0(_03253_),
    .I1(_03821_),
    .S(_03163_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18512_ (.I0(_03444_),
    .I1(_03822_),
    .S(_03093_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18513_ (.I0(_03354_),
    .I1(_03823_),
    .S(_03127_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18514_ (.A1(_03114_),
    .A2(_03824_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18515_ (.A1(_03819_),
    .A2(_03825_),
    .B(_03199_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18516_ (.A1(net3137),
    .A2(net3135),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18517_ (.A1(net3135),
    .A2(net3138),
    .B(_11342_[0]),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _18518_ (.A1(_03827_),
    .A2(_03766_),
    .A3(_03765_),
    .B(_03828_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _18519_ (.A1(net3132),
    .A2(_03829_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18520_ (.I0(_03339_),
    .I1(_03830_),
    .S(_03152_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _18521_ (.I0(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .I1(_03831_),
    .S(net3417),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18522_ (.A1(net3370),
    .A2(_03832_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18523_ (.A1(_08265_),
    .A2(_09366_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _18524_ (.A1(_03833_),
    .A2(_03826_),
    .A3(_06718_),
    .B(_03834_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18525_ (.I0(_03364_),
    .I1(_03365_),
    .S(net3470),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18526_ (.A1(net3400),
    .A2(_03836_),
    .B(_03564_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18527_ (.A1(_03835_),
    .A2(_03218_),
    .B(_03837_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_368_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_368_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_371_clk_i_regs (.I(clknet_6_3__leaf_clk_i_regs),
    .Z(clknet_leaf_371_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18530_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .I1(net466),
    .S(_03232_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18531_ (.I(_09383_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18532_ (.I0(_03403_),
    .I1(_03404_),
    .S(net3470),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18533_ (.A1(net3400),
    .A2(_03842_),
    .B(_03564_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18534_ (.A1(_11331_[0]),
    .A2(net3136),
    .A3(net3134),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18535_ (.A1(_11337_[0]),
    .A2(_11343_[0]),
    .A3(_11330_[0]),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18536_ (.A1(net3134),
    .A2(_11336_[0]),
    .B(_03845_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _18537_ (.A1(_03844_),
    .A2(_03747_),
    .A3(_03745_),
    .B(_03846_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18538_ (.A1(_11342_[0]),
    .A2(_03847_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18539_ (.A1(_03848_),
    .A2(net3132),
    .B(net3133),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18540_ (.A1(net3131),
    .A2(_03849_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18541_ (.I0(_03395_),
    .I1(_03850_),
    .S(_03152_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _18542_ (.I0(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .I1(_03851_),
    .S(net3417),
    .Z(_03852_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18543_ (.A1(_03852_),
    .A2(net3370),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18544_ (.A1(_03100_),
    .A2(_03597_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18545_ (.I(_11611_[0]),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18546_ (.A1(_03855_),
    .A2(_03180_),
    .B1(_03187_),
    .B2(_11612_[0]),
    .C1(_11615_[0]),
    .C2(net3206),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18547_ (.A1(_03091_),
    .A2(_03601_),
    .B(_03856_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18548_ (.A1(net366),
    .A2(_03707_),
    .B1(_03857_),
    .B2(_03298_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18549_ (.A1(_03853_),
    .A2(_03811_),
    .A3(_03854_),
    .A4(_03858_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _18550_ (.A1(_03841_),
    .A2(_03787_),
    .B(_03843_),
    .C(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_373_clk_i_regs (.I(clknet_6_2__leaf_clk_i_regs),
    .Z(clknet_leaf_373_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18552_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .I1(net578),
    .S(_03232_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18553_ (.A1(_03609_),
    .A2(net54),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18554_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net48),
    .B1(_03618_),
    .B2(\load_store_unit_i.rdata_q[21] ),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18555_ (.A1(net3470),
    .A2(_03609_),
    .A3(net40),
    .Z(_03864_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18556_ (.A1(_03076_),
    .A2(\load_store_unit_i.rdata_offset_q[0] ),
    .A3(net31),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18557_ (.A1(_03864_),
    .A2(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18558_ (.A1(\load_store_unit_i.rdata_q[5] ),
    .A2(_03613_),
    .B1(_03614_),
    .B2(\load_store_unit_i.rdata_q[13] ),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18559_ (.I0(_03866_),
    .I1(_03867_),
    .S(net3400),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18560_ (.A1(net3470),
    .A2(_03862_),
    .B1(_03863_),
    .B2(_03620_),
    .C(_03868_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18561_ (.A1(_03347_),
    .A2(_03815_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18562_ (.A1(_11435_[0]),
    .A2(_03181_),
    .B1(_03190_),
    .B2(net176),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18563_ (.A1(_11436_[0]),
    .A2(_03187_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18564_ (.A1(_11439_[0]),
    .A2(_03183_),
    .B(_03871_),
    .C(_03872_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18565_ (.I0(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .I1(_11210_[0]),
    .S(_03154_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18566_ (.A1(_03298_),
    .A2(_03873_),
    .B1(_03874_),
    .B2(net3370),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18567_ (.A1(_03245_),
    .A2(_03824_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _18568_ (.A1(_09522_),
    .A2(_03870_),
    .A3(_03875_),
    .A4(_03876_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18569_ (.I0(_03869_),
    .I1(_03877_),
    .S(_03218_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_375_clk_i_regs (.I(clknet_6_2__leaf_clk_i_regs),
    .Z(clknet_leaf_375_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18571_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .I1(_03878_),
    .S(_03629_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18572_ (.I(_11354_[0]),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18573_ (.A1(net3132),
    .A2(_03829_),
    .Z(_03881_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18574_ (.A1(net3133),
    .A2(_03881_),
    .B(net3131),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18575_ (.A1(_03880_),
    .A2(_03882_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18576_ (.A1(_11361_[0]),
    .A2(_03883_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_376_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_376_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18578_ (.I0(_03416_),
    .I1(_03884_),
    .S(_03152_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18579_ (.A1(net3417),
    .A2(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _18580_ (.A1(net3647),
    .A2(_03886_),
    .B(_03887_),
    .C(net3371),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18581_ (.A1(_03127_),
    .A2(_03425_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18582_ (.I0(_11417_[0]),
    .I1(net3252),
    .I2(_11622_[0]),
    .I3(_11614_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18583_ (.I0(_03820_),
    .I1(_03890_),
    .S(net3207),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18584_ (.I0(_03372_),
    .I1(_03371_),
    .I2(_03891_),
    .I3(_03772_),
    .S0(_03111_),
    .S1(_03093_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18585_ (.I0(_03436_),
    .I1(_03892_),
    .S(_03127_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18586_ (.A1(_11620_[0]),
    .A2(_03187_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18587_ (.A1(_11623_[0]),
    .A2(net3206),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18588_ (.A1(_11619_[0]),
    .A2(_03183_),
    .B(_03894_),
    .C(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18589_ (.A1(_03573_),
    .A2(_03889_),
    .B1(_03893_),
    .B2(_03114_),
    .C(_03896_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18590_ (.A1(_03199_),
    .A2(_03897_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18591_ (.A1(net169),
    .A2(_03707_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18592_ (.A1(_09399_),
    .A2(net3190),
    .A3(_03898_),
    .A4(_03899_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18593_ (.I0(_03409_),
    .I1(_03410_),
    .S(net3470),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18594_ (.A1(_03079_),
    .A2(_03901_),
    .B(_03564_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18595_ (.A1(_03888_),
    .A2(_03900_),
    .B(_03902_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_378_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_378_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18597_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .I1(net3053),
    .S(_03232_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18598_ (.A1(_11342_[0]),
    .A2(_11348_[0]),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18599_ (.A1(_11349_[0]),
    .A2(net3133),
    .B1(_03905_),
    .B2(_03847_),
    .C(_11355_[0]),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18600_ (.A1(_03906_),
    .A2(_03880_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18601_ (.A1(_03907_),
    .A2(_11361_[0]),
    .B(_11360_[0]),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18602_ (.A1(_11367_[0]),
    .A2(_03908_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18603_ (.I0(_03459_),
    .I1(_03909_),
    .S(_03152_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _18604_ (.I0(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .I1(_03910_),
    .S(net3417),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18605_ (.A1(_03135_),
    .A2(_03349_),
    .B(_03350_),
    .C(_03248_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _18606_ (.A1(_03131_),
    .A2(_03776_),
    .A3(_03912_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18607_ (.A1(_11631_[0]),
    .A2(net3206),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18608_ (.A1(_11627_[0]),
    .A2(_03183_),
    .B(_03914_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18609_ (.A1(_11628_[0]),
    .A2(_03187_),
    .B1(_03573_),
    .B2(_03913_),
    .C(_03915_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18610_ (.I0(_11413_[0]),
    .I1(_11421_[0]),
    .I2(_11626_[0]),
    .I3(_11618_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18611_ (.A1(net3207),
    .A2(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18612_ (.A1(net3207),
    .A2(_03592_),
    .B(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18613_ (.I0(_03321_),
    .I1(_03326_),
    .I2(_03806_),
    .I3(_03919_),
    .S0(_03163_),
    .S1(_03093_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18614_ (.I0(_03447_),
    .I1(_03920_),
    .S(_03127_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18615_ (.A1(net337),
    .A2(_03707_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18616_ (.A1(_03199_),
    .A2(_03916_),
    .B1(_03921_),
    .B2(_03100_),
    .C(_03922_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18617_ (.A1(net3370),
    .A2(_03911_),
    .B(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _18618_ (.I0(_09417_),
    .I1(_03924_),
    .S(_08265_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18619_ (.I0(_03467_),
    .I1(_03468_),
    .S(net3470),
    .Z(_03926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18620_ (.A1(net3400),
    .A2(_03926_),
    .B(_03564_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18621_ (.A1(_03925_),
    .A2(net3190),
    .B(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_379_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_379_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18623_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .I1(net434),
    .S(_03232_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18624_ (.I0(_03502_),
    .I1(_03503_),
    .S(net3470),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18625_ (.A1(net3400),
    .A2(_03930_),
    .B(_03564_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18626_ (.I(_11373_[0]),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18627_ (.I(_11367_[0]),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18628_ (.A1(net3133),
    .A2(_11354_[0]),
    .A3(_11360_[0]),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18629_ (.A1(net3132),
    .A2(_03829_),
    .B(_03934_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18630_ (.A1(_11355_[0]),
    .A2(_11354_[0]),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18631_ (.A1(_11361_[0]),
    .A2(_03936_),
    .B(_11360_[0]),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18632_ (.I(_11366_[0]),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18633_ (.A1(_03935_),
    .A2(_03933_),
    .A3(_03937_),
    .B(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18634_ (.A1(_03932_),
    .A2(_03939_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18635_ (.I0(_03495_),
    .I1(_03940_),
    .S(_03152_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _18636_ (.I0(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .I1(_03941_),
    .S(net3417),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18637_ (.I0(_11402_[0]),
    .I1(_11409_[0]),
    .I2(_11638_[0]),
    .I3(_11630_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18638_ (.I0(_03890_),
    .I1(_03943_),
    .S(net3207),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18639_ (.I0(_03821_),
    .I1(_03944_),
    .S(_03163_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _18640_ (.I0(_03267_),
    .I1(_03280_),
    .I2(_03945_),
    .I3(_03260_),
    .S0(_03248_),
    .S1(_03127_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18641_ (.A1(_03114_),
    .A2(_03946_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18642_ (.I(_11635_[0]),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18643_ (.A1(_03948_),
    .A2(_03180_),
    .B1(_03187_),
    .B2(_11636_[0]),
    .C1(_11639_[0]),
    .C2(net3206),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _18644_ (.A1(_03131_),
    .A2(_03475_),
    .A3(_03476_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18645_ (.A1(_03137_),
    .A2(_03245_),
    .A3(_03950_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18646_ (.A1(_03949_),
    .A2(_03951_),
    .B(_03199_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18647_ (.A1(_09440_),
    .A2(_03464_),
    .A3(_03947_),
    .A4(_03952_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18648_ (.A1(net258),
    .A2(_03707_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _18649_ (.A1(_03942_),
    .A2(net3370),
    .B(_03953_),
    .C(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18650_ (.A1(_03955_),
    .A2(_03931_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_380_clk_i_regs (.I(clknet_6_8__leaf_clk_i_regs),
    .Z(clknet_leaf_380_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18652_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .I1(net556),
    .S(_03232_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18653_ (.I0(_03535_),
    .I1(_03536_),
    .S(\load_store_unit_i.rdata_offset_q[1] ),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18654_ (.A1(net3400),
    .A2(_03958_),
    .B(_03564_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18655_ (.I(_03166_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18656_ (.I0(_03135_),
    .I1(_03960_),
    .S(_03600_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18657_ (.I(_11140_[0]),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18658_ (.A1(_11144_[0]),
    .A2(_03181_),
    .B1(_03180_),
    .B2(_03962_),
    .C1(_11141_[0]),
    .C2(_03187_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18659_ (.A1(_03091_),
    .A2(_03961_),
    .B(_03963_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18660_ (.I0(_11395_[0]),
    .I1(_11402_[0]),
    .I2(_11143_[0]),
    .I3(_11638_[0]),
    .S0(_06388_),
    .S1(_03114_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18661_ (.A1(_03163_),
    .A2(_03273_),
    .A3(_03917_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18662_ (.A1(_03163_),
    .A2(_03594_),
    .B1(_03965_),
    .B2(_03165_),
    .C(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18663_ (.I0(_03125_),
    .I1(_03967_),
    .S(_03093_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18664_ (.I0(_03531_),
    .I1(_03968_),
    .S(_03127_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18665_ (.A1(_03100_),
    .A2(_03969_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18666_ (.A1(net296),
    .A2(_03707_),
    .B1(_03964_),
    .B2(_03298_),
    .C(_03970_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18667_ (.A1(_03545_),
    .A2(_03523_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18668_ (.A1(_03932_),
    .A2(_11379_[0]),
    .A3(_03545_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18669_ (.I(_11379_[0]),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18670_ (.A1(_03974_),
    .A2(_11372_[0]),
    .A3(_03545_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _18671_ (.A1(_11361_[0]),
    .A2(_11367_[0]),
    .A3(_03907_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _18672_ (.A1(_11367_[0]),
    .A2(_11360_[0]),
    .B(_03976_),
    .C(_11366_[0]),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18673_ (.I0(_03973_),
    .I1(_03975_),
    .S(_03977_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _18674_ (.A1(_11373_[0]),
    .A2(_03974_),
    .A3(_11372_[0]),
    .A4(_03545_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18675_ (.I(_11372_[0]),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _18676_ (.A1(_11379_[0]),
    .A2(_03980_),
    .A3(_03545_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _18677_ (.A1(_03972_),
    .A2(_03978_),
    .A3(_03979_),
    .A4(_03981_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18678_ (.A1(net3647),
    .A2(_08240_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _18679_ (.A1(_03982_),
    .A2(net3647),
    .B(_03983_),
    .C(net3371),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _18680_ (.A1(_03984_),
    .A2(_03971_),
    .A3(_03811_),
    .Z(_03985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _18681_ (.A1(_09454_),
    .A2(_03787_),
    .B(_03985_),
    .C(_03959_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_381_clk_i_regs (.I(clknet_6_2__leaf_clk_i_regs),
    .Z(clknet_leaf_381_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18683_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .I1(net459),
    .S(_03232_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18684_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net50),
    .B1(_03618_),
    .B2(\load_store_unit_i.rdata_q[22] ),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18685_ (.A1(net3470),
    .A2(_03609_),
    .A3(net41),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18686_ (.A1(net32),
    .A2(_03613_),
    .B(_03989_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18687_ (.A1(\load_store_unit_i.rdata_q[6] ),
    .A2(_03613_),
    .B1(_03614_),
    .B2(\load_store_unit_i.rdata_q[14] ),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18688_ (.I0(_03990_),
    .I1(_03991_),
    .S(net3400),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18689_ (.A1(_03609_),
    .A2(_03988_),
    .B(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18690_ (.I(_03992_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18691_ (.I0(net55),
    .I1(_03994_),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18692_ (.I0(_03993_),
    .I1(_03995_),
    .S(_03076_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18693_ (.I0(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .I1(_11221_[0]),
    .S(_03154_),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18694_ (.A1(net3371),
    .A2(_03997_),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18695_ (.A1(_03091_),
    .A2(_03809_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18696_ (.A1(_11444_[0]),
    .A2(_03187_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18697_ (.A1(_11443_[0]),
    .A2(net3206),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18698_ (.A1(_11447_[0]),
    .A2(_03183_),
    .B(_04000_),
    .C(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18699_ (.A1(net177),
    .A2(_03190_),
    .B1(_03114_),
    .B2(_03800_),
    .C(_04002_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18700_ (.A1(_03199_),
    .A2(_04003_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18701_ (.A1(_09540_),
    .A2(_03998_),
    .A3(_03999_),
    .A4(_04004_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18702_ (.I0(_03996_),
    .I1(_04005_),
    .S(_03218_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_385_clk_i_regs (.I(clknet_6_2__leaf_clk_i_regs),
    .Z(clknet_leaf_385_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18704_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .I1(_04006_),
    .S(net3184),
    .Z(_00539_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18705_ (.A1(_03609_),
    .A2(_03617_),
    .A3(\load_store_unit_i.rdata_q[15] ),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18706_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(\load_store_unit_i.rdata_q[23] ),
    .B(_04008_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18707_ (.A1(_03609_),
    .A2(net42),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18708_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(\load_store_unit_i.rdata_q[23] ),
    .B1(net51),
    .B2(\load_store_unit_i.data_type_q[1] ),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _18709_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(_04009_),
    .B1(_04010_),
    .B2(net3400),
    .C1(_04011_),
    .C2(_03609_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18710_ (.I0(net33),
    .I1(\load_store_unit_i.rdata_q[7] ),
    .S(net3400),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18711_ (.I0(net56),
    .I1(_04013_),
    .S(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(_04014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18712_ (.I0(_04012_),
    .I1(_04014_),
    .S(_03076_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18713_ (.I0(_07175_),
    .I1(_09860_[0]),
    .S(_03154_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18714_ (.A1(_11451_[0]),
    .A2(net3206),
    .B1(_03190_),
    .B2(net178),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18715_ (.A1(_11455_[0]),
    .A2(_03183_),
    .B(_04017_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18716_ (.A1(_11452_[0]),
    .A2(_03187_),
    .B(_04018_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18717_ (.A1(_08233_),
    .A2(_04016_),
    .B1(_04019_),
    .B2(_03199_),
    .C(_08265_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18718_ (.A1(_03245_),
    .A2(_03775_),
    .B1(_03778_),
    .B2(_03347_),
    .C(_04020_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18719_ (.A1(_06718_),
    .A2(_09591_),
    .B(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18720_ (.I0(_04015_),
    .I1(_04022_),
    .S(_03218_),
    .Z(_04023_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_384_clk_i_regs (.I(clknet_6_2__leaf_clk_i_regs),
    .Z(clknet_leaf_384_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18722_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .I1(_04023_),
    .S(net3184),
    .Z(_00540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18723_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .I1(net3090),
    .S(net3184),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18724_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .I1(_03315_),
    .S(net3184),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18725_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .I1(net3089),
    .S(net3184),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18726_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .I1(net3093),
    .S(net3184),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_383_clk_i_regs (.I(clknet_6_2__leaf_clk_i_regs),
    .Z(clknet_leaf_383_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18728_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .I1(_03442_),
    .S(_03629_),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18729_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .I1(net3088),
    .S(_03629_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18730_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .I1(net3082),
    .S(_03629_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18731_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .I1(net3081),
    .S(_03629_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18732_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .I1(net3056),
    .S(_03629_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18733_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .I1(_03588_),
    .S(_03629_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18734_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .I1(net3067),
    .S(_03629_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18735_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .I1(net3066),
    .S(_03629_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18736_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .I1(net3065),
    .S(_03629_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18737_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .I1(net3080),
    .S(_03629_),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3090 (.I(_03221_),
    .Z(net3090));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18739_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .I1(net3076),
    .S(_03629_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18740_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .I1(net738),
    .S(_03629_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18741_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .I1(net3063),
    .S(_03629_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18742_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .I1(net3051),
    .S(_03629_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18743_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .I1(net466),
    .S(_03629_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18744_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .I1(net578),
    .S(_03629_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18745_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .I1(net3053),
    .S(_03629_),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18746_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .I1(net291),
    .S(_03629_),
    .Z(_00562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18747_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .I1(net555),
    .S(_03629_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18748_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .I1(net385),
    .S(_03629_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18749_ (.I(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18750_ (.A1(_04027_),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18751_ (.A1(_06737_),
    .A2(_03627_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18752_ (.A1(_04028_),
    .A2(_04029_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_393_clk_i_regs (.I(clknet_6_0__leaf_clk_i_regs),
    .Z(clknet_leaf_393_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18754_ (.A1(_03609_),
    .A2(net27),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18755_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net43),
    .B1(_03618_),
    .B2(\load_store_unit_i.rdata_q[16] ),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18756_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_03609_),
    .A3(net34),
    .Z(_04034_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18757_ (.A1(_03076_),
    .A2(net3471),
    .A3(net57),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18758_ (.A1(_04034_),
    .A2(_04035_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18759_ (.A1(\load_store_unit_i.rdata_q[0] ),
    .A2(_03613_),
    .B1(_03614_),
    .B2(\load_store_unit_i.rdata_q[8] ),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18760_ (.I0(_04036_),
    .I1(_04037_),
    .S(_03079_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18761_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_04032_),
    .B1(_03620_),
    .B2(_04033_),
    .C(_04038_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _18762_ (.A1(_08442_),
    .A2(_08444_),
    .A3(_01947_),
    .A4(_01957_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18763_ (.A1(_08445_),
    .A2(_01950_),
    .B(_04040_),
    .C(_03195_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18764_ (.I0(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .I1(_11184_[0]),
    .S(_03154_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18765_ (.A1(net3370),
    .A2(_04042_),
    .B(_06718_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18766_ (.A1(_11397_[0]),
    .A2(net3206),
    .B1(_03190_),
    .B2(\alu_adder_result_ex[0] ),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18767_ (.A1(_11400_[0]),
    .A2(_03183_),
    .B(_04044_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18768_ (.A1(_11398_[0]),
    .A2(_03187_),
    .B(_04045_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18769_ (.A1(_03091_),
    .A2(_03969_),
    .B1(_03961_),
    .B2(_03100_),
    .C(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18770_ (.A1(_03298_),
    .A2(_04047_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18771_ (.A1(_04041_),
    .A2(_04043_),
    .A3(_04048_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18772_ (.A1(_06718_),
    .A2(_08943_),
    .B(_03464_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _18773_ (.A1(_03228_),
    .A2(_04039_),
    .B1(_04049_),
    .B2(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_389_clk_i_regs (.I(clknet_6_2__leaf_clk_i_regs),
    .Z(clknet_leaf_389_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18775_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .A2(net3183),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18776_ (.A1(net3183),
    .A2(net3060),
    .B(_04053_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _18777_ (.A1(_03114_),
    .A2(_03137_),
    .A3(_03950_),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18778_ (.A1(_11404_[0]),
    .A2(_03181_),
    .B1(_03190_),
    .B2(\alu_adder_result_ex[1] ),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18779_ (.A1(_11407_[0]),
    .A2(_03183_),
    .B(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18780_ (.A1(_11405_[0]),
    .A2(_03187_),
    .B(_04054_),
    .C(_04056_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18781_ (.I0(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .I1(_11187_[0]),
    .S(_03154_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18782_ (.A1(net3370),
    .A2(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18783_ (.A1(_03199_),
    .A2(_04057_),
    .B(_04059_),
    .C(_09243_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18784_ (.A1(_03245_),
    .A2(_03946_),
    .B(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18785_ (.A1(net3470),
    .A2(_03609_),
    .A3(net35),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18786_ (.A1(_03076_),
    .A2(net3471),
    .A3(net58),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18787_ (.A1(_04062_),
    .A2(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18788_ (.A1(\load_store_unit_i.rdata_q[1] ),
    .A2(_03613_),
    .B1(_03614_),
    .B2(\load_store_unit_i.rdata_q[9] ),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18789_ (.I0(_04064_),
    .I1(_04065_),
    .S(_03079_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18790_ (.A1(_03076_),
    .A2(_03609_),
    .A3(net38),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18791_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net44),
    .B1(_03618_),
    .B2(\load_store_unit_i.rdata_q[17] ),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18792_ (.A1(_03620_),
    .A2(_04068_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18793_ (.A1(_03228_),
    .A2(_04066_),
    .A3(_04067_),
    .A4(_04069_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18794_ (.A1(_03218_),
    .A2(_04061_),
    .B(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_386_clk_i_regs (.I(clknet_6_2__leaf_clk_i_regs),
    .Z(clknet_leaf_386_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18796_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .I1(_04071_),
    .S(_04030_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18797_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net45),
    .B1(_03618_),
    .B2(\load_store_unit_i.rdata_q[18] ),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18798_ (.A1(_03076_),
    .A2(_03609_),
    .A3(net49),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18799_ (.A1(net3470),
    .A2(_03609_),
    .A3(net36),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18800_ (.A1(_03076_),
    .A2(\load_store_unit_i.rdata_offset_q[0] ),
    .A3(net28),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18801_ (.A1(_04075_),
    .A2(_04076_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18802_ (.A1(\load_store_unit_i.rdata_q[2] ),
    .A2(_03613_),
    .B1(_03614_),
    .B2(\load_store_unit_i.rdata_q[10] ),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18803_ (.I0(_04077_),
    .I1(_04078_),
    .S(net3400),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18804_ (.A1(_03620_),
    .A2(_04073_),
    .B(_04074_),
    .C(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18805_ (.A1(_11412_[0]),
    .A2(_03187_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18806_ (.A1(_11411_[0]),
    .A2(_03181_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18807_ (.A1(_11415_[0]),
    .A2(_03183_),
    .B(_04081_),
    .C(_04082_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18808_ (.A1(net171),
    .A2(_03190_),
    .B1(_03347_),
    .B2(_03913_),
    .C(_04083_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18809_ (.A1(_03199_),
    .A2(_04084_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18810_ (.I0(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .I1(_11189_[0]),
    .S(_03154_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18811_ (.A1(net3370),
    .A2(_04086_),
    .B(_08982_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18812_ (.A1(_03091_),
    .A2(_03921_),
    .B(_04085_),
    .C(_04087_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18813_ (.I0(_04080_),
    .I1(_04088_),
    .S(_03218_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_391_clk_i_regs (.I(clknet_6_0__leaf_clk_i_regs),
    .Z(clknet_leaf_391_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18815_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .I1(_04089_),
    .S(_04030_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18816_ (.A1(net3470),
    .A2(_03609_),
    .A3(net37),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18817_ (.A1(_03076_),
    .A2(net3471),
    .A3(net29),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18818_ (.A1(_04091_),
    .A2(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18819_ (.A1(\load_store_unit_i.rdata_q[3] ),
    .A2(_03613_),
    .B1(_03614_),
    .B2(\load_store_unit_i.rdata_q[11] ),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18820_ (.I0(_04093_),
    .I1(_04094_),
    .S(_03079_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18821_ (.A1(_03076_),
    .A2(_03609_),
    .A3(net52),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18822_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net46),
    .B1(_03618_),
    .B2(\load_store_unit_i.rdata_q[19] ),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18823_ (.A1(_03620_),
    .A2(_04097_),
    .Z(_04098_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18824_ (.A1(_03228_),
    .A2(_04095_),
    .A3(_04096_),
    .A4(_04098_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18825_ (.A1(_03245_),
    .A2(_03893_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18826_ (.A1(_11419_[0]),
    .A2(_03181_),
    .B1(_03190_),
    .B2(net174),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18827_ (.A1(_11423_[0]),
    .A2(_03183_),
    .B(_04101_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18828_ (.A1(_11420_[0]),
    .A2(_03187_),
    .B1(_03347_),
    .B2(_03889_),
    .C(_04102_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18829_ (.A1(_03199_),
    .A2(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18830_ (.I0(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .I1(_11197_[0]),
    .S(_03154_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18831_ (.A1(net3370),
    .A2(_04105_),
    .B(_09490_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18832_ (.A1(_03218_),
    .A2(_04100_),
    .A3(_04104_),
    .A4(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18833_ (.A1(_04099_),
    .A2(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_398_clk_i_regs (.I(clknet_6_0__leaf_clk_i_regs),
    .Z(clknet_leaf_398_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18835_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .I1(_04108_),
    .S(net3183),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18836_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .I1(_03625_),
    .S(_04030_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18837_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .I1(_03878_),
    .S(_04030_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18838_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .I1(_04006_),
    .S(_04030_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18839_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .I1(_04023_),
    .S(_04030_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18840_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .I1(net3090),
    .S(_04030_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_396_clk_i_regs (.I(clknet_6_0__leaf_clk_i_regs),
    .Z(clknet_leaf_396_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18842_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .I1(_03315_),
    .S(_04030_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18843_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .I1(net3089),
    .S(_04030_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18844_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .I1(net3093),
    .S(_04030_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18845_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .I1(_03442_),
    .S(_04030_),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18846_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .I1(net3088),
    .S(_04030_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18847_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .I1(net3082),
    .S(_04030_),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18848_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .I1(net3081),
    .S(_04030_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18849_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .I1(net3056),
    .S(net3183),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18850_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .I1(_03588_),
    .S(_04030_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18851_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .I1(net3067),
    .S(_04030_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3088 (.I(_03471_),
    .Z(net3088));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18853_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .I1(net3066),
    .S(_04030_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18854_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .I1(net3065),
    .S(_04030_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18855_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .I1(net3080),
    .S(_04030_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18856_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .I1(net3076),
    .S(net3183),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18857_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .I1(net3064),
    .S(_04030_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18858_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .I1(net3063),
    .S(_04030_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18859_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .I1(net584),
    .S(_04030_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18860_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .I1(net467),
    .S(_04030_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18861_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .I1(net578),
    .S(_04030_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18862_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .I1(net3053),
    .S(_04030_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18863_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .I1(net409),
    .S(_04030_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18864_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .I1(net556),
    .S(_04030_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18865_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .I1(net547),
    .S(net3183),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_397_clk_i_regs (.I(clknet_6_0__leaf_clk_i_regs),
    .Z(clknet_leaf_397_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18867_ (.A1(_08291_),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18868_ (.A1(_03627_),
    .A2(_04113_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18869_ (.A1(_04028_),
    .A2(_04114_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3086 (.I(_03939_),
    .Z(net3086));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18871_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .A2(_04115_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18872_ (.A1(net3060),
    .A2(_04115_),
    .B(_04117_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18873_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .I1(_04071_),
    .S(_04115_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18874_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .I1(_04089_),
    .S(_04115_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18875_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .I1(_04108_),
    .S(_04115_),
    .Z(_00600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18876_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .I1(_03625_),
    .S(_04115_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18877_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .I1(_03878_),
    .S(_04115_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18878_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .I1(_04006_),
    .S(_04115_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18879_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .I1(_04023_),
    .S(_04115_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18880_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .I1(net3090),
    .S(_04115_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3085 (.I(_01980_),
    .Z(net3085));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18882_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .I1(_03315_),
    .S(_04115_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18883_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .I1(net3089),
    .S(_04115_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18884_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .I1(net3093),
    .S(_04115_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18885_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .I1(_03442_),
    .S(_04115_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18886_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .I1(net3088),
    .S(_04115_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18887_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .I1(net3082),
    .S(_04115_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18888_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .I1(net3081),
    .S(_04115_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18889_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .I1(net3056),
    .S(_04115_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18890_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .I1(net627),
    .S(_04115_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18891_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .I1(net3067),
    .S(net3182),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3084 (.I(_01987_),
    .Z(net3084));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18893_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .I1(net3066),
    .S(_04115_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18894_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .I1(net3065),
    .S(net3182),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18895_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .I1(net3080),
    .S(_04115_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18896_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .I1(net3076),
    .S(_04115_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18897_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .I1(net738),
    .S(_04115_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18898_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .I1(net3063),
    .S(_04115_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18899_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .I1(net584),
    .S(_04115_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18900_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .I1(net466),
    .S(_04115_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18901_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .I1(net578),
    .S(net3182),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18902_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .I1(net3053),
    .S(net3182),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18903_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .I1(net434),
    .S(net3182),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18904_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .I1(net555),
    .S(net3182),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18905_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .I1(net3050),
    .S(_04115_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18906_ (.A1(_08291_),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18907_ (.A1(_03627_),
    .A2(_04120_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18908_ (.A1(_04028_),
    .A2(_04121_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3082 (.I(_03506_),
    .Z(net3082));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18910_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .A2(_04122_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18911_ (.A1(net3060),
    .A2(_04122_),
    .B(_04124_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18912_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .I1(_04071_),
    .S(_04122_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18913_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .I1(_04089_),
    .S(net3181),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18914_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .I1(_04108_),
    .S(_04122_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18915_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .I1(_03625_),
    .S(_04122_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18916_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .I1(_03878_),
    .S(_04122_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18917_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .I1(_04006_),
    .S(_04122_),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18918_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .I1(_04023_),
    .S(_04122_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18919_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .I1(net3090),
    .S(_04122_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_408_clk_i_regs (.I(clknet_6_1__leaf_clk_i_regs),
    .Z(clknet_leaf_408_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18921_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .I1(_03315_),
    .S(_04122_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18922_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .I1(net3089),
    .S(_04122_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18923_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .I1(net3093),
    .S(_04122_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18924_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .I1(_03442_),
    .S(net3181),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18925_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .I1(net3088),
    .S(net3181),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18926_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .I1(net3082),
    .S(_04122_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18927_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .I1(net3081),
    .S(_04122_),
    .Z(_00644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18928_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .I1(net3056),
    .S(_04122_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18929_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .I1(net627),
    .S(_04122_),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18930_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .I1(net3067),
    .S(net3181),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_407_clk_i_regs (.I(clknet_6_1__leaf_clk_i_regs),
    .Z(clknet_leaf_407_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18932_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .I1(net3066),
    .S(net3181),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18933_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .I1(net3065),
    .S(net3181),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18934_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .I1(net3080),
    .S(net3181),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18935_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .I1(net3076),
    .S(_04122_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18936_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .I1(net3064),
    .S(_04122_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18937_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .I1(net3063),
    .S(_04122_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18938_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .I1(net580),
    .S(_04122_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18939_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .I1(net3055),
    .S(_04122_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18940_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .I1(net578),
    .S(_04122_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18941_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .I1(net3053),
    .S(_04122_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18942_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .I1(net434),
    .S(_04122_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18943_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .I1(net555),
    .S(_04122_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18944_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .I1(net385),
    .S(_04122_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18945_ (.A1(_03628_),
    .A2(_04028_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_405_clk_i_regs (.I(clknet_6_1__leaf_clk_i_regs),
    .Z(clknet_leaf_405_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18947_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .A2(_04127_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18948_ (.A1(net3060),
    .A2(_04127_),
    .B(_04129_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18949_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .I1(_04071_),
    .S(_04127_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18950_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .I1(_04089_),
    .S(_04127_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18951_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .I1(_04108_),
    .S(_04127_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18952_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .I1(_03625_),
    .S(_04127_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18953_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .I1(_03878_),
    .S(_04127_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18954_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .I1(_04006_),
    .S(_04127_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18955_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .I1(_04023_),
    .S(_04127_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18956_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .I1(net3090),
    .S(_04127_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_404_clk_i_regs (.I(clknet_6_24__leaf_clk_i_regs),
    .Z(clknet_leaf_404_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18958_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .I1(_03315_),
    .S(_04127_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18959_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .I1(net3089),
    .S(_04127_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18960_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .I1(net3093),
    .S(_04127_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18961_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .I1(_03442_),
    .S(_04127_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18962_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .I1(net3088),
    .S(_04127_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18963_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .I1(net3082),
    .S(_04127_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18964_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .I1(net3081),
    .S(_04127_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18965_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .I1(net3056),
    .S(_04127_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18966_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .I1(net627),
    .S(_04127_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18967_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .I1(net3067),
    .S(_04127_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_403_clk_i_regs (.I(clknet_6_24__leaf_clk_i_regs),
    .Z(clknet_leaf_403_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18969_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .I1(net3066),
    .S(_04127_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18970_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .I1(net3065),
    .S(_04127_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18971_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .I1(net3080),
    .S(_04127_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18972_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .I1(net3076),
    .S(_04127_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18973_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .I1(net3064),
    .S(_04127_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18974_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .I1(net3063),
    .S(_04127_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18975_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .I1(net580),
    .S(_04127_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18976_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .I1(net466),
    .S(_04127_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18977_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .I1(net578),
    .S(_04127_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18978_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .I1(net3053),
    .S(_04127_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18979_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .I1(net409),
    .S(_04127_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18980_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .I1(net556),
    .S(_04127_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18981_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .I1(net385),
    .S(_04127_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18982_ (.A1(_04027_),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18983_ (.A1(_04029_),
    .A2(_04132_),
    .Z(_04133_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_402_clk_i_regs (.I(clknet_6_24__leaf_clk_i_regs),
    .Z(clknet_leaf_402_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18985_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .A2(_04133_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18986_ (.A1(net3060),
    .A2(_04133_),
    .B(_04135_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18987_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .I1(_04071_),
    .S(net3180),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18988_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .I1(_04089_),
    .S(_04133_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18989_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .I1(_04108_),
    .S(_04133_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18990_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .I1(_03625_),
    .S(_04133_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18991_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .I1(_03878_),
    .S(_04133_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18992_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .I1(_04006_),
    .S(_04133_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18993_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .I1(_04023_),
    .S(net3180),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18994_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .I1(net3090),
    .S(net3180),
    .Z(_00701_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_400_clk_i_regs (.I(clknet_6_24__leaf_clk_i_regs),
    .Z(clknet_leaf_400_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18996_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .I1(_03315_),
    .S(net3180),
    .Z(_00702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18997_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .I1(net3089),
    .S(net3180),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18998_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .I1(net3093),
    .S(net3180),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18999_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .I1(_03442_),
    .S(_04133_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19000_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .I1(net3088),
    .S(_04133_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19001_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .I1(net3082),
    .S(_04133_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19002_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .I1(net3081),
    .S(_04133_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19003_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .I1(net3056),
    .S(_04133_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19004_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .I1(_03588_),
    .S(_04133_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19005_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .I1(net3067),
    .S(_04133_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_399_clk_i_regs (.I(clknet_6_24__leaf_clk_i_regs),
    .Z(clknet_leaf_399_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19007_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .I1(net3066),
    .S(_04133_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19008_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .I1(net3065),
    .S(_04133_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19009_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .I1(net3080),
    .S(_04133_),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19010_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .I1(net3076),
    .S(_04133_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19011_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .I1(net738),
    .S(net3180),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19012_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .I1(net3063),
    .S(_04133_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19013_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .I1(net584),
    .S(_04133_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19014_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .I1(net3055),
    .S(_04133_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19015_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .I1(net3054),
    .S(_04133_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19016_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .I1(net3053),
    .S(_04133_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19017_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .I1(net434),
    .S(_04133_),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19018_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .I1(net3052),
    .S(_04133_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19019_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .I1(net385),
    .S(_04133_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19020_ (.A1(_04114_),
    .A2(_04132_),
    .Z(_04138_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3081 (.I(_03540_),
    .Z(net3081));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19022_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .A2(_04138_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19023_ (.A1(net3060),
    .A2(_04138_),
    .B(_04140_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19024_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .I1(_04071_),
    .S(_04138_),
    .Z(_00726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19025_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .I1(_04089_),
    .S(_04138_),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19026_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .I1(_04108_),
    .S(_04138_),
    .Z(_00728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19027_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .I1(_03625_),
    .S(_04138_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19028_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .I1(_03878_),
    .S(_04138_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19029_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .I1(_04006_),
    .S(_04138_),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19030_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .I1(_04023_),
    .S(_04138_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19031_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .I1(net3090),
    .S(_04138_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_412_clk_i_regs (.I(clknet_6_25__leaf_clk_i_regs),
    .Z(clknet_leaf_412_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19033_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .I1(_03315_),
    .S(_04138_),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19034_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .I1(net3089),
    .S(_04138_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19035_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .I1(net3093),
    .S(_04138_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19036_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .I1(_03442_),
    .S(_04138_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19037_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .I1(net3088),
    .S(_04138_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19038_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .I1(net3082),
    .S(_04138_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19039_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .I1(net3081),
    .S(_04138_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19040_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .I1(net3056),
    .S(_04138_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19041_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .I1(net627),
    .S(_04138_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19042_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .I1(net3067),
    .S(_04138_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_409_clk_i_regs (.I(clknet_6_1__leaf_clk_i_regs),
    .Z(clknet_leaf_409_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19044_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .I1(net3066),
    .S(_04138_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19045_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .I1(net3065),
    .S(_04138_),
    .Z(_00745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19046_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .I1(net3080),
    .S(_04138_),
    .Z(_00746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19047_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .I1(net3076),
    .S(_04138_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19048_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .I1(net737),
    .S(_04138_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19049_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .I1(net3063),
    .S(_04138_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19050_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .I1(net3051),
    .S(_04138_),
    .Z(_00750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19051_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .I1(net467),
    .S(_04138_),
    .Z(_00751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19052_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .I1(net3054),
    .S(_04138_),
    .Z(_00752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19053_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .I1(net3053),
    .S(_04138_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19054_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .I1(net291),
    .S(_04138_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19055_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .I1(net556),
    .S(_04138_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19056_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .I1(net3050),
    .S(_04138_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19057_ (.A1(_04121_),
    .A2(_04132_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_417_clk_i_regs (.I(clknet_6_26__leaf_clk_i_regs),
    .Z(clknet_leaf_417_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19059_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .A2(_04143_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19060_ (.A1(net3060),
    .A2(_04143_),
    .B(_04145_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19061_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .I1(_04071_),
    .S(_04143_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19062_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .I1(_04089_),
    .S(_04143_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19063_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .I1(_04108_),
    .S(_04143_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19064_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .I1(_03625_),
    .S(_04143_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19065_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .I1(_03878_),
    .S(_04143_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19066_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .I1(_04006_),
    .S(_04143_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19067_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .I1(_04023_),
    .S(_04143_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19068_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .I1(net3090),
    .S(_04143_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_416_clk_i_regs (.I(clknet_6_26__leaf_clk_i_regs),
    .Z(clknet_leaf_416_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19070_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .I1(_03315_),
    .S(_04143_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19071_ (.A1(_06740_),
    .A2(_04114_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_418_clk_i_regs (.I(clknet_6_26__leaf_clk_i_regs),
    .Z(clknet_leaf_418_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19073_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .A2(_04147_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19074_ (.A1(net3060),
    .A2(_04147_),
    .B(_04149_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19075_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .I1(net3089),
    .S(_04143_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19076_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .I1(net3093),
    .S(_04143_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19077_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .I1(_03442_),
    .S(_04143_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19078_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .I1(net3088),
    .S(_04143_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19079_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .I1(net3082),
    .S(_04143_),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19080_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .I1(net3081),
    .S(_04143_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19081_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .I1(net3056),
    .S(_04143_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19082_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .I1(net627),
    .S(_04143_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19083_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .I1(net3067),
    .S(_04143_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3637 (.I(net480),
    .Z(net3637));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19085_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .I1(net3066),
    .S(_04143_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19086_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .I1(_04071_),
    .S(_04147_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19087_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .I1(net3065),
    .S(_04143_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19088_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .I1(net3080),
    .S(_04143_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19089_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .I1(net3076),
    .S(_04143_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19090_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .I1(net737),
    .S(_04143_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19091_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .I1(net3063),
    .S(_04143_),
    .Z(_00783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19092_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .I1(net584),
    .S(_04143_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19093_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .I1(net3055),
    .S(_04143_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19094_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .I1(net3054),
    .S(_04143_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19095_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .I1(net3053),
    .S(_04143_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19096_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .I1(net291),
    .S(_04143_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19097_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .I1(_04089_),
    .S(_04147_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19098_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .I1(net555),
    .S(_04143_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19099_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .I1(net385),
    .S(_04143_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19100_ (.A1(_03628_),
    .A2(_04132_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3080 (.I(_03717_),
    .Z(net3080));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19102_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .A2(_04151_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19103_ (.A1(net3060),
    .A2(_04151_),
    .B(_04153_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19104_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .I1(_04071_),
    .S(net3179),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19105_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .I1(_04089_),
    .S(_04151_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19106_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .I1(_04108_),
    .S(_04151_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19107_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .I1(_03625_),
    .S(_04151_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19108_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .I1(_03878_),
    .S(_04151_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19109_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .I1(_04006_),
    .S(net3179),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19110_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .I1(_04023_),
    .S(net3179),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19111_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .I1(_04108_),
    .S(_04147_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19112_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .I1(net3090),
    .S(net3179),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3079 (.I(_03851_),
    .Z(net3079));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19114_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .I1(_03315_),
    .S(net3179),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19115_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .I1(net3089),
    .S(net3179),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19116_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .I1(net3093),
    .S(net3179),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19117_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .I1(_03442_),
    .S(_04151_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19118_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .I1(net3088),
    .S(_04151_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19119_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .I1(net3082),
    .S(_04151_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19120_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .I1(net3081),
    .S(_04151_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19121_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .I1(net3056),
    .S(_04151_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19122_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .I1(net627),
    .S(_04151_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19123_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .I1(_03625_),
    .S(_04147_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19124_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .I1(net3067),
    .S(_04151_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_419_clk_i_regs (.I(clknet_6_27__leaf_clk_i_regs),
    .Z(clknet_leaf_419_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19126_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .I1(net3066),
    .S(_04151_),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19127_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .I1(net3065),
    .S(_04151_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19128_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .I1(net3080),
    .S(_04151_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19129_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .I1(net3076),
    .S(_04151_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19130_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .I1(net738),
    .S(net3179),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19131_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .I1(net3063),
    .S(_04151_),
    .Z(_00818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19132_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .I1(net580),
    .S(_04151_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19133_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .I1(net466),
    .S(_04151_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19134_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .I1(net579),
    .S(_04151_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19135_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .I1(_03878_),
    .S(_04147_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19136_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .I1(net3053),
    .S(_04151_),
    .Z(_00823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19137_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .I1(net291),
    .S(_04151_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19138_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .I1(net555),
    .S(_04151_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19139_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .I1(net385),
    .S(_04151_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19140_ (.A1(_03230_),
    .A2(_04029_),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_428_clk_i_regs (.I(clknet_6_3__leaf_clk_i_regs),
    .Z(clknet_leaf_428_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19142_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .A2(_04156_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19143_ (.A1(net3060),
    .A2(_04156_),
    .B(_04158_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19144_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .I1(_04071_),
    .S(net3178),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19145_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .I1(_04089_),
    .S(_04156_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19146_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .I1(_04108_),
    .S(_04156_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_427_clk_i_regs (.I(clknet_6_3__leaf_clk_i_regs),
    .Z(clknet_leaf_427_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19148_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .I1(_03625_),
    .S(_04156_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_426_clk_i_regs (.I(clknet_6_3__leaf_clk_i_regs),
    .Z(clknet_leaf_426_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19150_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .I1(_03878_),
    .S(_04156_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19151_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .I1(_04006_),
    .S(_04147_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_424_clk_i_regs (.I(clknet_6_4__leaf_clk_i_regs),
    .Z(clknet_leaf_424_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19153_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .I1(_04006_),
    .S(_04156_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19154_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .I1(_04023_),
    .S(_04156_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_423_clk_i_regs (.I(clknet_6_4__leaf_clk_i_regs),
    .Z(clknet_leaf_423_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19156_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .I1(net3090),
    .S(_04156_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_422_clk_i_regs (.I(clknet_6_4__leaf_clk_i_regs),
    .Z(clknet_leaf_422_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_420_clk_i_regs (.I(clknet_6_4__leaf_clk_i_regs),
    .Z(clknet_leaf_420_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19159_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .I1(_03315_),
    .S(net3178),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3074 (.I(_03910_),
    .Z(net3074));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19161_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .I1(net3089),
    .S(net3178),
    .Z(_00838_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_430_clk_i_regs (.I(clknet_6_6__leaf_clk_i_regs),
    .Z(clknet_leaf_430_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19163_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .I1(net3093),
    .S(_04156_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_433_clk_i_regs (.I(clknet_6_6__leaf_clk_i_regs),
    .Z(clknet_leaf_433_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19165_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .I1(_03442_),
    .S(_04156_),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_431_clk_i_regs (.I(clknet_6_6__leaf_clk_i_regs),
    .Z(clknet_leaf_431_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19167_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .I1(net3088),
    .S(_04156_),
    .Z(_00841_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3076 (.I(_03739_),
    .Z(net3076));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19169_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .I1(net3082),
    .S(net3178),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_453_clk_i_regs (.I(clknet_6_27__leaf_clk_i_regs),
    .Z(clknet_leaf_453_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19171_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .I1(net3081),
    .S(net3178),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_450_clk_i_regs (.I(clknet_6_4__leaf_clk_i_regs),
    .Z(clknet_leaf_450_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19173_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .I1(_04023_),
    .S(_04147_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_449_clk_i_regs (.I(clknet_6_4__leaf_clk_i_regs),
    .Z(clknet_leaf_449_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19175_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .I1(net3056),
    .S(_04156_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_447_clk_i_regs (.I(clknet_6_4__leaf_clk_i_regs),
    .Z(clknet_leaf_447_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19177_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .I1(_03588_),
    .S(_04156_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_446_clk_i_regs (.I(clknet_6_5__leaf_clk_i_regs),
    .Z(clknet_leaf_446_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19179_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .I1(net3067),
    .S(_04156_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_443_clk_i_regs (.I(clknet_6_7__leaf_clk_i_regs),
    .Z(clknet_leaf_443_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_442_clk_i_regs (.I(clknet_6_7__leaf_clk_i_regs),
    .Z(clknet_leaf_442_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19182_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .I1(net3066),
    .S(_04156_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_440_clk_i_regs (.I(clknet_6_7__leaf_clk_i_regs),
    .Z(clknet_leaf_440_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19184_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .I1(net3065),
    .S(_04156_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_436_clk_i_regs (.I(clknet_6_12__leaf_clk_i_regs),
    .Z(clknet_leaf_436_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19186_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .I1(net3080),
    .S(_04156_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_435_clk_i_regs (.I(clknet_6_6__leaf_clk_i_regs),
    .Z(clknet_leaf_435_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19188_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .I1(net3076),
    .S(_04156_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3101 (.I(_03686_),
    .Z(net3101));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19190_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .I1(net738),
    .S(net3178),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_456_clk_i_regs (.I(clknet_6_27__leaf_clk_i_regs),
    .Z(clknet_leaf_456_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19192_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .I1(net3063),
    .S(net3178),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3102 (.I(_03661_),
    .Z(net3102));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19194_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .I1(net584),
    .S(_04156_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19195_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .I1(net3090),
    .S(_04147_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3077 (.I(_02146_),
    .Z(net3077));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19197_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .I1(net467),
    .S(_04156_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3071 (.I(_05085_),
    .Z(net3071));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19199_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .I1(net579),
    .S(_04156_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_462_clk_i_regs (.I(clknet_6_30__leaf_clk_i_regs),
    .Z(clknet_leaf_462_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19201_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .I1(net3053),
    .S(_04156_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3067 (.I(_03647_),
    .Z(net3067));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19203_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .I1(net434),
    .S(_04156_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3066 (.I(_03670_),
    .Z(net3066));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19205_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .I1(net3052),
    .S(_04156_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_465_clk_i_regs (.I(clknet_6_5__leaf_clk_i_regs),
    .Z(clknet_leaf_465_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19207_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .I1(net3050),
    .S(_04156_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19208_ (.A1(_03230_),
    .A2(_04114_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3065 (.I(_03694_),
    .Z(net3065));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19210_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .A2(_04189_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19211_ (.A1(net3060),
    .A2(_04189_),
    .B(_04191_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3062 (.I(_03886_),
    .Z(net3062));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19213_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .I1(_04071_),
    .S(_04189_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_466_clk_i_regs (.I(clknet_6_5__leaf_clk_i_regs),
    .Z(clknet_leaf_466_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19215_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .I1(_04089_),
    .S(_04189_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3060 (.I(_04051_),
    .Z(net3060));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19217_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .I1(_04108_),
    .S(_04189_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3058 (.I(_05101_),
    .Z(net3058));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19219_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .I1(_03315_),
    .S(_04147_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19220_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .I1(_03625_),
    .S(_04189_),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19221_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .I1(_03878_),
    .S(_04189_),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19222_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .I1(_04006_),
    .S(_04189_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19223_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .I1(_04023_),
    .S(_04189_),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19224_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .I1(net3090),
    .S(_04189_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3057 (.I(_05256_),
    .Z(net3057));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19226_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .I1(_03315_),
    .S(_04189_),
    .Z(_00872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19227_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .I1(net3089),
    .S(_04189_),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19228_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .I1(net3093),
    .S(_04189_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19229_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .I1(_03442_),
    .S(_04189_),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19230_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .I1(net3088),
    .S(_04189_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19231_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .I1(net3089),
    .S(_04147_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19232_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .I1(net3082),
    .S(_04189_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19233_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .I1(net3081),
    .S(_04189_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19234_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .I1(net3056),
    .S(_04189_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19235_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .I1(_03588_),
    .S(_04189_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19236_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .I1(net3067),
    .S(_04189_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3056 (.I(_03567_),
    .Z(net3056));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19238_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .I1(net3066),
    .S(_04189_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19239_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .I1(net3065),
    .S(_04189_),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19240_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .I1(net3080),
    .S(_04189_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19241_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .I1(net3076),
    .S(_04189_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19242_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .I1(net737),
    .S(_04189_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19243_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .I1(net3093),
    .S(_04147_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19244_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .I1(net3063),
    .S(_04189_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19245_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .I1(net580),
    .S(_04189_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19246_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .I1(net467),
    .S(_04189_),
    .Z(_00891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19247_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .I1(net579),
    .S(_04189_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19248_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .I1(net3053),
    .S(_04189_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19249_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .I1(net434),
    .S(_04189_),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19250_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .I1(net555),
    .S(_04189_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19251_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .I1(net3050),
    .S(_04189_),
    .Z(_00896_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place3055 (.I(_03838_),
    .Z(net3055));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19253_ (.A1(_03230_),
    .A2(_04121_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3054 (.I(net487),
    .Z(net3054));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19255_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .A2(_04199_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19256_ (.A1(net3060),
    .A2(_04199_),
    .B(_04201_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19257_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .I1(_04071_),
    .S(_04199_),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19258_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .I1(_03442_),
    .S(_04147_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19259_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .I1(_04089_),
    .S(_04199_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19260_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .I1(_04108_),
    .S(_04199_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19261_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .I1(_03625_),
    .S(_04199_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19262_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .I1(_03878_),
    .S(_04199_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19263_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .I1(_04006_),
    .S(_04199_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19264_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .I1(_04023_),
    .S(_04199_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19265_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .I1(net3090),
    .S(_04199_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3053 (.I(_03903_),
    .Z(net3053));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19267_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .I1(_03315_),
    .S(_04199_),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19268_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .I1(net3089),
    .S(_04199_),
    .Z(_00908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19269_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .I1(net3093),
    .S(_04199_),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19270_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .I1(net3088),
    .S(_04147_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19271_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .I1(_03442_),
    .S(_04199_),
    .Z(_00911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19272_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .I1(net3088),
    .S(_04199_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19273_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .I1(net3082),
    .S(_04199_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19274_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .I1(net3081),
    .S(_04199_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19275_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .I1(net3056),
    .S(_04199_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19276_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .I1(net627),
    .S(_04199_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19277_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .I1(net3067),
    .S(_04199_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_467_clk_i_regs (.I(clknet_6_30__leaf_clk_i_regs),
    .Z(clknet_leaf_467_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19279_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .I1(net3066),
    .S(_04199_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19280_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .I1(net3065),
    .S(_04199_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19281_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .I1(net3080),
    .S(_04199_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19282_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .I1(net3082),
    .S(_04147_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19283_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .I1(net3076),
    .S(_04199_),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19284_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .I1(net738),
    .S(_04199_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19285_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .I1(net3063),
    .S(_04199_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19286_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .I1(net580),
    .S(_04199_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19287_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .I1(net467),
    .S(_04199_),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19288_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .I1(net579),
    .S(_04199_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19289_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .I1(net3053),
    .S(_04199_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19290_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .I1(net464),
    .S(_04199_),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19291_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .I1(net556),
    .S(_04199_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19292_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .I1(net459),
    .S(_04199_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19293_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .I1(net3081),
    .S(_04147_),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19294_ (.A1(_03230_),
    .A2(_03628_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place3052 (.I(_03956_),
    .Z(net3052));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19296_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .A2(_04204_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19297_ (.A1(net3060),
    .A2(_04204_),
    .B(_04206_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19298_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .I1(_04071_),
    .S(_04204_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19299_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .I1(_04089_),
    .S(_04204_),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19300_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .I1(_04108_),
    .S(_04204_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19301_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .I1(_03625_),
    .S(_04204_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19302_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .I1(_03878_),
    .S(_04204_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19303_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .I1(_04006_),
    .S(_04204_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19304_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .I1(_04023_),
    .S(_04204_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19305_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .I1(net3090),
    .S(_04204_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3670 (.I(net139),
    .Z(net3670));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19307_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .I1(_03315_),
    .S(_04204_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19308_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .I1(net3056),
    .S(_04147_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19309_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .I1(net3089),
    .S(_04204_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19310_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .I1(net3093),
    .S(_04204_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19311_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .I1(_03442_),
    .S(_04204_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19312_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .I1(net3088),
    .S(_04204_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19313_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .I1(net3082),
    .S(_04204_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19314_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .I1(net3081),
    .S(_04204_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19315_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .I1(net3056),
    .S(_04204_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19316_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .I1(net627),
    .S(_04204_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19317_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .I1(net3067),
    .S(_04204_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3653 (.I(\cs_registers_i.pc_if_i[1] ),
    .Z(net3653));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19319_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .I1(net3066),
    .S(_04204_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19320_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .I1(net627),
    .S(_04147_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19321_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .I1(net3065),
    .S(_04204_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19322_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .I1(net3080),
    .S(_04204_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19323_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .I1(net3076),
    .S(_04204_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19324_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .I1(net3064),
    .S(_04204_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19325_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .I1(net3063),
    .S(_04204_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19326_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .I1(net3051),
    .S(_04204_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19327_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .I1(net3055),
    .S(_04204_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19328_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .I1(net578),
    .S(_04204_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19329_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .I1(net3053),
    .S(_04204_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19330_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .I1(net464),
    .S(_04204_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19331_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .I1(net3067),
    .S(_04147_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19332_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .I1(net3052),
    .S(_04204_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19333_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .I1(net459),
    .S(_04204_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19334_ (.A1(_06740_),
    .A2(_03229_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19335_ (.A1(_06737_),
    .A2(_04209_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22914__3 (.ZN(net252));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19337_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .A2(_04210_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19338_ (.A1(net3060),
    .A2(_04210_),
    .B(_04212_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19339_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .I1(_04071_),
    .S(net3177),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19340_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .I1(_04089_),
    .S(_04210_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19341_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .I1(_04108_),
    .S(_04210_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19342_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .I1(_03625_),
    .S(_04210_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19343_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .I1(_03878_),
    .S(_04210_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19344_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .I1(_04006_),
    .S(_04210_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19345_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .I1(_04023_),
    .S(_04210_),
    .Z(_00975_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3652 (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(net3652));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19347_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .I1(net3066),
    .S(_04147_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19348_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .I1(net3090),
    .S(net3177),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3651 (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(net3651));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19350_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .I1(_03315_),
    .S(net3177),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19351_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .I1(net3089),
    .S(_04210_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19352_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .I1(net3093),
    .S(_04210_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19353_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .I1(_03442_),
    .S(_04210_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19354_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .I1(net3088),
    .S(_04210_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19355_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .I1(net3082),
    .S(net3177),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19356_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .I1(net3081),
    .S(net3177),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19357_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .I1(net3056),
    .S(_04210_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19358_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .I1(net627),
    .S(_04210_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19359_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .I1(net3065),
    .S(_04147_),
    .Z(_00987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19360_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .I1(net3067),
    .S(_04210_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3089 (.I(_03368_),
    .Z(net3089));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19362_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .I1(net3066),
    .S(_04210_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19363_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .I1(net3065),
    .S(_04210_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19364_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .I1(net3080),
    .S(_04210_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19365_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .I1(net3076),
    .S(_04210_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19366_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .I1(net737),
    .S(net3177),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19367_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .I1(net3063),
    .S(_04210_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19368_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .I1(net580),
    .S(_04210_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19369_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .I1(net3055),
    .S(_04210_),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19370_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .I1(net578),
    .S(_04210_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19371_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .I1(net3080),
    .S(_04147_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19372_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .I1(net3053),
    .S(_04210_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19373_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .I1(net464),
    .S(_04210_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19374_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .I1(net3052),
    .S(_04210_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19375_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .I1(net547),
    .S(_04210_),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19376_ (.A1(_04113_),
    .A2(_04209_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3636 (.I(net3634),
    .Z(net3636));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19378_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .A2(_04216_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19379_ (.A1(net3060),
    .A2(_04216_),
    .B(_04218_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19380_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .I1(_04071_),
    .S(_04216_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19381_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .I1(_04089_),
    .S(net3176),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19382_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .I1(_04108_),
    .S(_04216_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19383_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .I1(_03625_),
    .S(_04216_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19384_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .I1(_03878_),
    .S(_04216_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19385_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .I1(net3076),
    .S(_04147_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19386_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .I1(_04006_),
    .S(_04216_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19387_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .I1(_04023_),
    .S(_04216_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19388_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .I1(net3090),
    .S(_04216_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3444 (.I(net3443),
    .Z(net3444));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19390_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .I1(_03315_),
    .S(_04216_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19391_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .I1(net3089),
    .S(_04216_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19392_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .I1(net3093),
    .S(_04216_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19393_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .I1(_03442_),
    .S(net3176),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19394_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .I1(net3088),
    .S(net3176),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19395_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .I1(net3082),
    .S(_04216_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19396_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .I1(net3081),
    .S(_04216_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19397_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .I1(net3064),
    .S(_04147_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19398_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .I1(net3056),
    .S(_04216_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19399_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .I1(net627),
    .S(_04216_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19400_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .I1(net3067),
    .S(net3176),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk_i_regs (.I(clknet_6_51__leaf_clk_i_regs),
    .Z(clknet_leaf_15_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19402_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .I1(net3066),
    .S(net3176),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19403_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .I1(net3065),
    .S(net3176),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19404_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .I1(net3080),
    .S(_04216_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19405_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .I1(net3076),
    .S(_04216_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19406_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .I1(net737),
    .S(_04216_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19407_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .I1(net3063),
    .S(_04216_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19408_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .I1(net580),
    .S(_04216_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19409_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .I1(net3063),
    .S(_04147_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19410_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .I1(net3055),
    .S(_04216_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19411_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .I1(net578),
    .S(_04216_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19412_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .I1(net3053),
    .S(_04216_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19413_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .I1(net409),
    .S(_04216_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19414_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .I1(net3052),
    .S(_04216_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19415_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .I1(net547),
    .S(_04216_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19416_ (.A1(_04120_),
    .A2(_04209_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk_i_regs (.I(clknet_6_51__leaf_clk_i_regs),
    .Z(clknet_leaf_13_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19418_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .A2(_04221_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19419_ (.A1(net3060),
    .A2(_04221_),
    .B(_04223_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19420_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .I1(_04071_),
    .S(_04221_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19421_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .I1(_04089_),
    .S(net3175),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19422_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .I1(_04108_),
    .S(_04221_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19423_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .I1(net3051),
    .S(_04147_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19424_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .I1(_03625_),
    .S(_04221_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19425_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .I1(_03878_),
    .S(_04221_),
    .Z(_01044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19426_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .I1(_04006_),
    .S(_04221_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19427_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .I1(_04023_),
    .S(_04221_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19428_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .I1(net3090),
    .S(_04221_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_39_clk_i_regs (.I(clknet_6_54__leaf_clk_i_regs),
    .Z(clknet_leaf_39_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19430_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .I1(_03315_),
    .S(_04221_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19431_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .I1(net3089),
    .S(_04221_),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19432_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .I1(net3093),
    .S(_04221_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19433_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .I1(_03442_),
    .S(net3175),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19434_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .I1(net3088),
    .S(net3175),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19435_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .I1(net466),
    .S(_04147_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19436_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .I1(net3082),
    .S(_04221_),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19437_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .I1(net3081),
    .S(_04221_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19438_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .I1(net3056),
    .S(_04221_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19439_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .I1(_03588_),
    .S(_04221_),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19440_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .I1(net3067),
    .S(net3175),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3443 (.I(_06367_),
    .Z(net3443));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19442_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .I1(net3066),
    .S(net3175),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19443_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .I1(net3065),
    .S(net3175),
    .Z(_01060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19444_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .I1(net3080),
    .S(_04221_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19445_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .I1(net3076),
    .S(_04221_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19446_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .I1(net737),
    .S(_04221_),
    .Z(_01063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19447_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .I1(net3054),
    .S(_04147_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19448_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .I1(net3063),
    .S(_04221_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19449_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .I1(net584),
    .S(_04221_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19450_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .I1(net466),
    .S(_04221_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19451_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .I1(net578),
    .S(_04221_),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19452_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .I1(net3053),
    .S(_04221_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19453_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .I1(net409),
    .S(_04221_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19454_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .I1(net556),
    .S(_04221_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19455_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .I1(net3050),
    .S(_04221_),
    .Z(_01072_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19456_ (.A1(_03223_),
    .A2(_04209_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3665 (.I(net144),
    .Z(net3665));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19458_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .A2(net3174),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19459_ (.A1(net3060),
    .A2(net3174),
    .B(_04228_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19460_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .I1(_04071_),
    .S(_04226_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19461_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .I1(net3053),
    .S(_04147_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19462_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .I1(_04089_),
    .S(net3174),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19463_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .I1(_04108_),
    .S(net3174),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19464_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .I1(_03625_),
    .S(_04226_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19465_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .I1(_03878_),
    .S(_04226_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19466_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .I1(_04006_),
    .S(_04226_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19467_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .I1(_04023_),
    .S(_04226_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19468_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .I1(net3090),
    .S(_04226_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3584 (.I(net3583),
    .Z(net3584));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19470_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .I1(_03315_),
    .S(_04226_),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19471_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .I1(net3089),
    .S(_04226_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19472_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .I1(net3093),
    .S(_04226_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19473_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .I1(net291),
    .S(_04147_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19474_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .I1(_03442_),
    .S(net3174),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19475_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .I1(net3088),
    .S(net3174),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19476_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .I1(net3082),
    .S(_04226_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19477_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .I1(net3081),
    .S(_04226_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19478_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .I1(net3056),
    .S(net3174),
    .Z(_01091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19479_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .I1(net627),
    .S(_04226_),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19480_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .I1(net3067),
    .S(net3174),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3442 (.I(_06367_),
    .Z(net3442));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19482_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .I1(net3066),
    .S(net3174),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19483_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .I1(net3065),
    .S(_04226_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19484_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .I1(net3080),
    .S(_04226_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19485_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .I1(net3052),
    .S(_04147_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19486_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .I1(net3076),
    .S(net3174),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19487_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .I1(net737),
    .S(_04226_),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19488_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .I1(net3063),
    .S(net3174),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19489_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .I1(net3051),
    .S(_04226_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19490_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .I1(net466),
    .S(_04226_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19491_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .I1(net3054),
    .S(_04226_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19492_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .I1(net3053),
    .S(_04226_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19493_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .I1(net464),
    .S(_04226_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19494_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .I1(net556),
    .S(_04226_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19495_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .I1(net547),
    .S(net3174),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19496_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .I1(net459),
    .S(_04147_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19497_ (.A1(_03229_),
    .A2(_04028_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19498_ (.A1(_06737_),
    .A2(_04231_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_90_clk_i_regs (.I(clknet_6_62__leaf_clk_i_regs),
    .Z(clknet_leaf_90_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19500_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .A2(_04232_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19501_ (.A1(net3060),
    .A2(_04232_),
    .B(_04234_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19502_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .I1(_04071_),
    .S(net3173),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19503_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .I1(_04089_),
    .S(_04232_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19504_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .I1(_04108_),
    .S(_04232_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19505_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .I1(_03625_),
    .S(_04232_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19506_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .I1(_03878_),
    .S(_04232_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19507_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .I1(_04006_),
    .S(net3173),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19508_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .I1(_04023_),
    .S(net3173),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19509_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .I1(net3090),
    .S(net3173),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3235 (.I(_08567_),
    .Z(net3235));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19511_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .I1(_03315_),
    .S(net3173),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19512_ (.A1(_06740_),
    .A2(_04121_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_38_clk_i_regs (.I(clknet_6_54__leaf_clk_i_regs),
    .Z(clknet_leaf_38_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19514_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .A2(_04236_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19515_ (.A1(net3060),
    .A2(net3172),
    .B(_04238_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19516_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .I1(net3089),
    .S(net3173),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19517_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .I1(net3093),
    .S(net3173),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19518_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .I1(_03442_),
    .S(_04232_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19519_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .I1(net3088),
    .S(_04232_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19520_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .I1(net3082),
    .S(_04232_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19521_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .I1(net3081),
    .S(_04232_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19522_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .I1(net3056),
    .S(_04232_),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19523_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .I1(net627),
    .S(_04232_),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19524_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .I1(net3067),
    .S(_04232_),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3215 (.I(net298),
    .Z(net3215));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19526_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .I1(net3066),
    .S(_04232_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19527_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .I1(_04071_),
    .S(_04236_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19528_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .I1(net3065),
    .S(_04232_),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19529_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .I1(net3080),
    .S(_04232_),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19530_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .I1(net3076),
    .S(_04232_),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19531_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .I1(net737),
    .S(_04232_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19532_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .I1(net3063),
    .S(_04232_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19533_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .I1(net580),
    .S(_04232_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19534_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .I1(net467),
    .S(_04232_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19535_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .I1(net579),
    .S(_04232_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19536_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .I1(net3053),
    .S(_04232_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19537_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .I1(net434),
    .S(_04232_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19538_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .I1(_04089_),
    .S(_04236_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19539_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .I1(net3052),
    .S(_04232_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19540_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .I1(net3050),
    .S(_04232_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19541_ (.A1(_04113_),
    .A2(_04231_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3612 (.I(net333),
    .Z(net3612));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19543_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .A2(_04240_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19544_ (.A1(net3060),
    .A2(_04240_),
    .B(_04242_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19545_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .I1(_04071_),
    .S(_04240_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19546_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .I1(_04089_),
    .S(_04240_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19547_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .I1(_04108_),
    .S(_04240_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19548_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .I1(_03625_),
    .S(_04240_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19549_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .I1(_03878_),
    .S(_04240_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19550_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .I1(_04006_),
    .S(_04240_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19551_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .I1(_04023_),
    .S(_04240_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19552_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .I1(_04108_),
    .S(_04236_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output249 (.I(net249),
    .Z(instr_req_o));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19554_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .I1(net3090),
    .S(_04240_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output248 (.I(net248),
    .Z(instr_addr_o[9]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output247 (.I(net247),
    .Z(instr_addr_o[8]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19557_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .I1(_03315_),
    .S(_04240_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output246 (.I(net246),
    .Z(instr_addr_o[7]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19559_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .I1(net3089),
    .S(_04240_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output245 (.I(net245),
    .Z(instr_addr_o[6]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19561_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .I1(net3093),
    .S(_04240_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output244 (.I(net244),
    .Z(instr_addr_o[5]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19563_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .I1(_03442_),
    .S(_04240_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output243 (.I(net243),
    .Z(instr_addr_o[4]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19565_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .I1(net3088),
    .S(_04240_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output242 (.I(net242),
    .Z(instr_addr_o[3]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19567_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .I1(net3082),
    .S(_04240_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 output241 (.I(net241),
    .Z(instr_addr_o[31]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19569_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .I1(net3081),
    .S(_04240_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 output240 (.I(net240),
    .Z(instr_addr_o[30]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19571_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .I1(net3056),
    .S(_04240_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output239 (.I(net239),
    .Z(instr_addr_o[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19573_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .I1(_03588_),
    .S(_04240_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 output238 (.I(net238),
    .Z(instr_addr_o[29]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19575_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .I1(_03625_),
    .S(_04236_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output237 (.I(net237),
    .Z(instr_addr_o[28]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19577_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .I1(net3067),
    .S(_04240_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 output236 (.I(net236),
    .Z(instr_addr_o[27]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 output235 (.I(net235),
    .Z(instr_addr_o[26]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19580_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .I1(net3066),
    .S(_04240_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output234 (.I(net234),
    .Z(instr_addr_o[25]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19582_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .I1(net3065),
    .S(_04240_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output233 (.I(net233),
    .Z(instr_addr_o[24]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19584_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .I1(net3080),
    .S(net3171),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 output232 (.I(net232),
    .Z(instr_addr_o[23]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19586_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .I1(net3076),
    .S(_04240_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output231 (.I(net231),
    .Z(instr_addr_o[22]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19588_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .I1(net737),
    .S(_04240_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output230 (.I(net230),
    .Z(instr_addr_o[21]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19590_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .I1(net3063),
    .S(_04240_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output229 (.I(net229),
    .Z(instr_addr_o[20]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19592_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .I1(net580),
    .S(net3171),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output228 (.I(net228),
    .Z(instr_addr_o[19]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19594_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .I1(net466),
    .S(net3171),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output227 (.I(net227),
    .Z(instr_addr_o[18]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19596_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .I1(net3054),
    .S(net3171),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output226 (.I(net226),
    .Z(instr_addr_o[17]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19598_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .I1(_03878_),
    .S(net3172),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output225 (.I(net225),
    .Z(instr_addr_o[16]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19600_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .I1(net3053),
    .S(net3171),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output224 (.I(net224),
    .Z(instr_addr_o[15]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19602_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .I1(net464),
    .S(net3171),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output223 (.I(net223),
    .Z(instr_addr_o[14]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19604_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .I1(net555),
    .S(net3171),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output222 (.I(net222),
    .Z(instr_addr_o[13]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19606_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .I1(net547),
    .S(_04240_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19607_ (.A1(_04120_),
    .A2(_04231_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output221 (.I(net221),
    .Z(instr_addr_o[12]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19609_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .A2(_04271_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19610_ (.A1(net3060),
    .A2(_04271_),
    .B(_04273_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output220 (.I(net220),
    .Z(instr_addr_o[11]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19612_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .I1(_04071_),
    .S(_04271_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output219 (.I(net219),
    .Z(instr_addr_o[10]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19614_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .I1(_04089_),
    .S(_04271_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output218 (.I(net218),
    .Z(data_we_o));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19616_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .I1(_04108_),
    .S(_04271_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19617_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .I1(_03625_),
    .S(_04271_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19618_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .I1(_03878_),
    .S(net3170),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output217 (.I(net217),
    .Z(data_wdata_o[9]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19620_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .I1(_04006_),
    .S(_04236_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19621_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .I1(_04006_),
    .S(_04271_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output216 (.I(net216),
    .Z(data_wdata_o[8]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19623_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .I1(_04023_),
    .S(_04271_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19624_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .I1(net3090),
    .S(_04271_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output215 (.I(net215),
    .Z(data_wdata_o[7]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19626_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .I1(_03315_),
    .S(_04271_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19627_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .I1(net3089),
    .S(_04271_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19628_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .I1(net3093),
    .S(_04271_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19629_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .I1(_03442_),
    .S(_04271_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19630_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .I1(net3088),
    .S(_04271_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19631_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .I1(net3082),
    .S(net3170),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19632_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .I1(net3081),
    .S(net3170),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19633_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .I1(_04023_),
    .S(_04236_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19634_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .I1(net3056),
    .S(_04271_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19635_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .I1(_03588_),
    .S(_04271_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19636_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .I1(net3067),
    .S(_04271_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output214 (.I(net214),
    .Z(data_wdata_o[6]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19638_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .I1(net3066),
    .S(_04271_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19639_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .I1(net3065),
    .S(_04271_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19640_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .I1(net3080),
    .S(_04271_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19641_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .I1(net3076),
    .S(_04271_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19642_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .I1(net3064),
    .S(net3170),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19643_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .I1(net3063),
    .S(net3170),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19644_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .I1(net580),
    .S(_04271_),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19645_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .I1(net3090),
    .S(_04236_),
    .Z(_01207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19646_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .I1(net3055),
    .S(_04271_),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19647_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .I1(net578),
    .S(_04271_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19648_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .I1(net3053),
    .S(_04271_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19649_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .I1(net409),
    .S(_04271_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19650_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .I1(net555),
    .S(_04271_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19651_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .I1(net547),
    .S(_04271_),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19652_ (.A1(_03223_),
    .A2(_04231_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output213 (.I(net213),
    .Z(data_wdata_o[5]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19654_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .A2(_04281_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19655_ (.A1(net3060),
    .A2(_04281_),
    .B(_04283_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19656_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .I1(_04071_),
    .S(_04281_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19657_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .I1(_04089_),
    .S(_04281_),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19658_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .I1(_04108_),
    .S(_04281_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output212 (.I(net212),
    .Z(data_wdata_o[4]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19660_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .I1(_03315_),
    .S(_04236_),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19661_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .I1(_03625_),
    .S(_04281_),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19662_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .I1(_03878_),
    .S(net3169),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19663_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .I1(_04006_),
    .S(_04281_),
    .Z(_01221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19664_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .I1(_04023_),
    .S(_04281_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19665_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .I1(net3090),
    .S(_04281_),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output211 (.I(net211),
    .Z(data_wdata_o[3]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19667_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .I1(_03315_),
    .S(_04281_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19668_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .I1(net3089),
    .S(_04281_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19669_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .I1(net3093),
    .S(_04281_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19670_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .I1(_03442_),
    .S(_04281_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19671_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .I1(net3088),
    .S(_04281_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19672_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .I1(net3089),
    .S(_04236_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19673_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .I1(net3082),
    .S(net3169),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19674_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .I1(net3081),
    .S(net3169),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19675_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .I1(net3056),
    .S(_04281_),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19676_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .I1(_03588_),
    .S(_04281_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19677_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .I1(net3067),
    .S(_04281_),
    .Z(_01234_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output210 (.I(net210),
    .Z(data_wdata_o[31]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19679_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .I1(net3066),
    .S(_04281_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19680_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .I1(net3065),
    .S(_04281_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19681_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .I1(net3080),
    .S(_04281_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19682_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .I1(net3076),
    .S(_04281_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19683_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .I1(net737),
    .S(net3169),
    .Z(_01239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19684_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .I1(net3093),
    .S(_04236_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19685_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .I1(net3063),
    .S(net3169),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19686_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .I1(net580),
    .S(_04281_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19687_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .I1(net466),
    .S(_04281_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19688_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .I1(net578),
    .S(_04281_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19689_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .I1(net3053),
    .S(_04281_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19690_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .I1(net409),
    .S(_04281_),
    .Z(_01246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19691_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .I1(net555),
    .S(_04281_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19692_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .I1(net459),
    .S(_04281_),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19693_ (.A1(_03229_),
    .A2(_04132_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19694_ (.A1(_06737_),
    .A2(_04287_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output209 (.I(net209),
    .Z(data_wdata_o[30]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19696_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .A2(_04288_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19697_ (.A1(net3060),
    .A2(_04288_),
    .B(_04290_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19698_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .I1(_04071_),
    .S(_04288_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19699_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .I1(_03442_),
    .S(_04236_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19700_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .I1(_04089_),
    .S(net3168),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19701_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .I1(_04108_),
    .S(_04288_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19702_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .I1(_03625_),
    .S(_04288_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19703_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .I1(_03878_),
    .S(_04288_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19704_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .I1(_04006_),
    .S(_04288_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19705_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .I1(_04023_),
    .S(_04288_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19706_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .I1(net3090),
    .S(_04288_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output208 (.I(net208),
    .Z(data_wdata_o[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19708_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .I1(_03315_),
    .S(_04288_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19709_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .I1(net3089),
    .S(_04288_),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19710_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .I1(net3093),
    .S(_04288_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19711_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .I1(net3088),
    .S(_04236_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19712_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .I1(_03442_),
    .S(net3168),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19713_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .I1(net3088),
    .S(net3168),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19714_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .I1(net3082),
    .S(_04288_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19715_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .I1(net3081),
    .S(_04288_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19716_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .I1(net3056),
    .S(_04288_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19717_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .I1(_03588_),
    .S(_04288_),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19718_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .I1(net3067),
    .S(net3168),
    .Z(_01269_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output207 (.I(net207),
    .Z(data_wdata_o[29]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19720_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .I1(net3066),
    .S(net3168),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19721_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .I1(net3065),
    .S(_04288_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19722_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .I1(net3080),
    .S(_04288_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19723_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .I1(net3082),
    .S(net3172),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19724_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .I1(net3076),
    .S(_04288_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19725_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .I1(net3064),
    .S(_04288_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19726_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .I1(net3063),
    .S(_04288_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19727_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .I1(net580),
    .S(net3168),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19728_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .I1(net466),
    .S(_04288_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19729_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .I1(net579),
    .S(_04288_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19730_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .I1(net3053),
    .S(_04288_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19731_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .I1(net409),
    .S(_04288_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19732_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .I1(net556),
    .S(_04288_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19733_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .I1(net3050),
    .S(_04288_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19734_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .I1(net3081),
    .S(net3172),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19735_ (.A1(_04113_),
    .A2(_04287_),
    .Z(_04293_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output206 (.I(net206),
    .Z(data_wdata_o[28]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19737_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .A2(_04293_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19738_ (.A1(net3060),
    .A2(_04293_),
    .B(_04295_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19739_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .I1(_04071_),
    .S(_04293_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19740_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .I1(_04089_),
    .S(net3167),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19741_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .I1(_04108_),
    .S(_04293_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19742_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .I1(_03625_),
    .S(_04293_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19743_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .I1(_03878_),
    .S(_04293_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19744_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .I1(_04006_),
    .S(_04293_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19745_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .I1(_04023_),
    .S(_04293_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19746_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .I1(net3090),
    .S(_04293_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output205 (.I(net205),
    .Z(data_wdata_o[27]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19748_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .I1(_03315_),
    .S(_04293_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19749_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .I1(net3056),
    .S(_04236_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19750_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .I1(net3089),
    .S(_04293_),
    .Z(_01296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19751_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .I1(net3093),
    .S(_04293_),
    .Z(_01297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19752_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .I1(_03442_),
    .S(net3167),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19753_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .I1(net3088),
    .S(net3167),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19754_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .I1(net3082),
    .S(_04293_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19755_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .I1(net3081),
    .S(_04293_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19756_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .I1(net3056),
    .S(_04293_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19757_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .I1(_03588_),
    .S(_04293_),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19758_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .I1(net3067),
    .S(net3167),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output204 (.I(net204),
    .Z(data_wdata_o[26]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19760_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .I1(net3066),
    .S(net3167),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19761_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .I1(_03588_),
    .S(_04236_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19762_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .I1(net3065),
    .S(_04293_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19763_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .I1(net3080),
    .S(_04293_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19764_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .I1(net3076),
    .S(_04293_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19765_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .I1(net738),
    .S(_04293_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19766_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .I1(net3063),
    .S(_04293_),
    .Z(_01311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19767_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .I1(net3051),
    .S(net3167),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19768_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .I1(net466),
    .S(_04293_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19769_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .I1(net578),
    .S(_04293_),
    .Z(_01314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19770_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .I1(net3053),
    .S(_04293_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19771_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .I1(net291),
    .S(_04293_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19772_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .I1(net3067),
    .S(_04236_),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19773_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .I1(net3052),
    .S(_04293_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19774_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .I1(net459),
    .S(_04293_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19775_ (.A1(_04120_),
    .A2(_04287_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output203 (.I(net203),
    .Z(data_wdata_o[25]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19777_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .A2(_04298_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19778_ (.A1(net3060),
    .A2(_04298_),
    .B(_04300_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19779_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .I1(_04071_),
    .S(_04298_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19780_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .I1(_04089_),
    .S(net3166),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19781_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .I1(_04108_),
    .S(_04298_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19782_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .I1(_03625_),
    .S(_04298_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19783_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .I1(_03878_),
    .S(_04298_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19784_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .I1(_04006_),
    .S(_04298_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19785_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .I1(_04023_),
    .S(_04298_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output202 (.I(net202),
    .Z(data_wdata_o[24]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19787_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .I1(net3066),
    .S(_04236_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19788_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .I1(net3090),
    .S(_04298_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output201 (.I(net201),
    .Z(data_wdata_o[23]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19790_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .I1(_03315_),
    .S(_04298_),
    .Z(_01330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19791_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .I1(net3089),
    .S(_04298_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19792_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .I1(net3093),
    .S(_04298_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19793_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .I1(_03442_),
    .S(net3166),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19794_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .I1(net3088),
    .S(net3166),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19795_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .I1(net3082),
    .S(_04298_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19796_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .I1(net3081),
    .S(_04298_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19797_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .I1(net3056),
    .S(_04298_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19798_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .I1(net627),
    .S(_04298_),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19799_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .I1(net3065),
    .S(_04236_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19800_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .I1(net3067),
    .S(net3166),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output200 (.I(net200),
    .Z(data_wdata_o[22]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19802_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .I1(net3066),
    .S(net3166),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19803_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .I1(net3065),
    .S(_04298_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19804_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .I1(net3080),
    .S(_04298_),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19805_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .I1(net3076),
    .S(_04298_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19806_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .I1(net737),
    .S(_04298_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19807_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .I1(net3063),
    .S(_04298_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19808_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .I1(net3051),
    .S(net3166),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19809_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .I1(net466),
    .S(_04298_),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19810_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .I1(net3054),
    .S(_04298_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19811_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .I1(net3080),
    .S(_04236_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19812_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .I1(net3053),
    .S(_04298_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19813_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .I1(net464),
    .S(_04298_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19814_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .I1(net555),
    .S(_04298_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19815_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .I1(net459),
    .S(_04298_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19816_ (.A1(_03223_),
    .A2(_04287_),
    .Z(_04304_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output199 (.I(net199),
    .Z(data_wdata_o[21]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19818_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .A2(_04304_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19819_ (.A1(net3060),
    .A2(_04304_),
    .B(_04306_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19820_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .I1(_04071_),
    .S(_04304_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19821_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .I1(_04089_),
    .S(net3165),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19822_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .I1(_04108_),
    .S(_04304_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19823_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .I1(_03625_),
    .S(_04304_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19824_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .I1(_03878_),
    .S(_04304_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19825_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .I1(net3076),
    .S(_04236_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19826_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .I1(_04006_),
    .S(_04304_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19827_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .I1(_04023_),
    .S(_04304_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19828_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .I1(net3090),
    .S(_04304_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output198 (.I(net198),
    .Z(data_wdata_o[20]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19830_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .I1(_03315_),
    .S(_04304_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19831_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .I1(net3089),
    .S(_04304_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19832_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .I1(net3093),
    .S(_04304_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19833_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .I1(_03442_),
    .S(net3165),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19834_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .I1(net3088),
    .S(net3165),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19835_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .I1(net3082),
    .S(_04304_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19836_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .I1(net3081),
    .S(_04304_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19837_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .I1(net737),
    .S(net3172),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19838_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .I1(net3056),
    .S(_04304_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19839_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .I1(_03588_),
    .S(_04304_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19840_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .I1(net3067),
    .S(net3165),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output197 (.I(net197),
    .Z(data_wdata_o[1]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19842_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .I1(net3066),
    .S(net3165),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19843_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .I1(net3065),
    .S(_04304_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19844_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .I1(net3080),
    .S(_04304_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19845_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .I1(net3076),
    .S(_04304_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19846_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .I1(net737),
    .S(_04304_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19847_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .I1(net3063),
    .S(_04304_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19848_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .I1(net580),
    .S(net3165),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19849_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .I1(net3063),
    .S(net3172),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19850_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .I1(net466),
    .S(_04304_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19851_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .I1(net3054),
    .S(_04304_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19852_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .I1(net3053),
    .S(_04304_),
    .Z(_01386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19853_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .I1(net291),
    .S(_04304_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19854_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .I1(net555),
    .S(_04304_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19855_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .I1(net459),
    .S(_04304_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19856_ (.A1(_06737_),
    .A2(_03231_),
    .Z(_04309_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output196 (.I(net196),
    .Z(data_wdata_o[19]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19858_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .A2(_04309_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19859_ (.A1(net3060),
    .A2(_04309_),
    .B(_04311_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19860_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .I1(_04071_),
    .S(_04309_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19861_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .I1(_04089_),
    .S(_04309_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19862_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .I1(_04108_),
    .S(_04309_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19863_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .I1(net584),
    .S(_04236_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19864_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .I1(_03625_),
    .S(net3164),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19865_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .I1(_03878_),
    .S(net3164),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19866_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .I1(_04006_),
    .S(_04309_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19867_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .I1(_04023_),
    .S(_04309_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19868_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .I1(net3090),
    .S(_04309_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output195 (.I(net195),
    .Z(data_wdata_o[18]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19870_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .I1(_03315_),
    .S(_04309_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19871_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .I1(net3089),
    .S(_04309_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19872_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .I1(net3093),
    .S(_04309_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19873_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .I1(_03442_),
    .S(_04309_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19874_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .I1(net3088),
    .S(_04309_),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19875_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .I1(net467),
    .S(_04236_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19876_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .I1(net3082),
    .S(net3164),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19877_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .I1(net3081),
    .S(net3164),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19878_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .I1(net3056),
    .S(_04309_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19879_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .I1(_03588_),
    .S(net3164),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19880_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .I1(net3067),
    .S(_04309_),
    .Z(_01410_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output194 (.I(net194),
    .Z(data_wdata_o[17]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19882_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .I1(net3066),
    .S(_04309_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19883_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .I1(net3065),
    .S(_04309_),
    .Z(_01412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19884_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .I1(net3080),
    .S(_04309_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19885_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .I1(net3076),
    .S(_04309_),
    .Z(_01414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19886_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .I1(net738),
    .S(net3164),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19887_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .I1(net578),
    .S(_04236_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19888_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .I1(net3063),
    .S(_04309_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19889_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .I1(net3051),
    .S(_04309_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19890_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .I1(net467),
    .S(_04309_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19891_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .I1(net579),
    .S(_04309_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19892_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .I1(net3053),
    .S(_04309_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19893_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .I1(net464),
    .S(_04309_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19894_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .I1(net555),
    .S(_04309_),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19895_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .I1(net385),
    .S(_04309_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19896_ (.A1(_03231_),
    .A2(_04113_),
    .Z(_04314_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output193 (.I(net193),
    .Z(data_wdata_o[16]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19898_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .A2(_04314_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19899_ (.A1(net3060),
    .A2(net3163),
    .B(_04316_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19900_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .I1(_04071_),
    .S(_04314_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19901_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .I1(net3053),
    .S(_04236_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19902_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .I1(_04089_),
    .S(net3163),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19903_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .I1(_04108_),
    .S(net3163),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19904_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .I1(_03625_),
    .S(_04314_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19905_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .I1(_03878_),
    .S(_04314_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19906_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .I1(_04006_),
    .S(_04314_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19907_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .I1(_04023_),
    .S(_04314_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19908_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .I1(net3090),
    .S(_04314_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output192 (.I(net192),
    .Z(data_wdata_o[15]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19910_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .I1(_03315_),
    .S(_04314_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19911_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .I1(net3089),
    .S(_04314_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19912_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .I1(net3093),
    .S(_04314_),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19913_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .I1(net434),
    .S(_04236_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19914_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .I1(_03442_),
    .S(_04314_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19915_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .I1(net3088),
    .S(_04314_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19916_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .I1(net3082),
    .S(_04314_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19917_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .I1(net3081),
    .S(_04314_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19918_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .I1(net3056),
    .S(_04314_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19919_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .I1(net627),
    .S(net3163),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19920_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .I1(net3067),
    .S(_04314_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output191 (.I(net191),
    .Z(data_wdata_o[14]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19922_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .I1(net3066),
    .S(net3163),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19923_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .I1(net3065),
    .S(_04314_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19924_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .I1(net3080),
    .S(_04314_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19925_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .I1(net555),
    .S(_04236_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19926_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .I1(net3076),
    .S(_04314_),
    .Z(_01450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19927_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .I1(net737),
    .S(_04314_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19928_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .I1(net3063),
    .S(_04314_),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19929_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .I1(net580),
    .S(_04314_),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19930_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .I1(net3055),
    .S(_04314_),
    .Z(_01454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19931_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .I1(net579),
    .S(_04314_),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19932_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .I1(net3053),
    .S(_04314_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19933_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .I1(net409),
    .S(_04314_),
    .Z(_01457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19934_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .I1(net555),
    .S(_04314_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19935_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .I1(net547),
    .S(net3163),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19936_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .I1(net385),
    .S(_04236_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _19937_ (.A1(_03231_),
    .A2(_04120_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output190 (.I(net190),
    .Z(data_wdata_o[13]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19939_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .A2(_04319_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19940_ (.A1(net3060),
    .A2(_04319_),
    .B(_04321_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19941_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .I1(_04071_),
    .S(_04319_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19942_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .I1(_04089_),
    .S(net3162),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19943_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .I1(_04108_),
    .S(net3162),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19944_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .I1(_03625_),
    .S(_04319_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19945_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .I1(_03878_),
    .S(_04319_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19946_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .I1(_04006_),
    .S(_04319_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19947_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .I1(_04023_),
    .S(_04319_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19948_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .I1(net3090),
    .S(_04319_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output189 (.I(net189),
    .Z(data_wdata_o[12]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19950_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .I1(_03315_),
    .S(_04319_),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19951_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .A2(_03629_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19952_ (.A1(_03629_),
    .A2(net3060),
    .B(_04323_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19953_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .I1(net3089),
    .S(_04319_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19954_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .I1(net3093),
    .S(_04319_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19955_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .I1(_03442_),
    .S(net3162),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19956_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .I1(net3088),
    .S(net3162),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19957_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .I1(net3082),
    .S(_04319_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19958_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .I1(net3081),
    .S(_04319_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19959_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .I1(net3056),
    .S(_04319_),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19960_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .I1(_03588_),
    .S(_04319_),
    .Z(_01479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19961_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .I1(net3067),
    .S(net3162),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output188 (.I(net188),
    .Z(data_wdata_o[11]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19963_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .I1(net3066),
    .S(net3162),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19964_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .I1(_04071_),
    .S(net3184),
    .Z(_01482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19965_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .I1(net3065),
    .S(_04319_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19966_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .I1(net3080),
    .S(_04319_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19967_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .I1(net3076),
    .S(_04319_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19968_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .I1(net3064),
    .S(_04319_),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19969_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .I1(net3063),
    .S(_04319_),
    .Z(_01487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19970_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .I1(net580),
    .S(_04319_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19971_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .I1(net466),
    .S(_04319_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19972_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .I1(net578),
    .S(_04319_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19973_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .I1(net3053),
    .S(_04319_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19974_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .I1(net291),
    .S(_04319_),
    .Z(_01492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19975_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .I1(_04089_),
    .S(_03629_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19976_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .I1(net555),
    .S(_04319_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19977_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .I1(net3050),
    .S(net3162),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _19978_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .A2(_03232_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19979_ (.A1(_03232_),
    .A2(net3060),
    .B(_04325_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19980_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .I1(_04071_),
    .S(_03232_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19981_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .I1(_04089_),
    .S(_03232_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19982_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .I1(_04108_),
    .S(_03232_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19983_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .I1(_03625_),
    .S(net3185),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19984_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .I1(_03878_),
    .S(net3185),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19985_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .I1(_04006_),
    .S(_03232_),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19986_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .I1(_04023_),
    .S(_03232_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19987_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .I1(_04108_),
    .S(_03629_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _19988_ (.A1(net3473),
    .A2(\cs_registers_i.dcsr_q[2] ),
    .B(net60),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19989_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_04326_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _19990_ (.A1(_02019_),
    .A2(_04327_),
    .Z(_04328_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output187 (.I(net187),
    .Z(data_wdata_o[10]));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19992_ (.I(_08384_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _19993_ (.A1(net3440),
    .A2(_08948_),
    .A3(_11149_[0]),
    .A4(_08378_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _19994_ (.A1(_11149_[0]),
    .A2(net3412),
    .A3(_04330_),
    .B(_04331_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _19995_ (.A1(net3473),
    .A2(net3425),
    .A3(_08308_),
    .Z(_04333_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _19996_ (.A1(_08949_),
    .A2(_04332_),
    .A3(_04333_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _19997_ (.A1(_08383_),
    .A2(_08400_),
    .A3(_02386_),
    .A4(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19998_ (.I(_04335_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _19999_ (.A1(\id_stage_i.controller_i.instr_fetch_err_i ),
    .A2(_08393_),
    .A3(_04336_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20000_ (.A1(_08265_),
    .A2(_08374_),
    .B(_04337_),
    .C(_06782_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20001_ (.A1(_06345_),
    .A2(_08391_),
    .B(_04335_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20002_ (.A1(_04338_),
    .A2(_04339_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20003_ (.A1(_08363_),
    .A2(_04340_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20004_ (.A1(_04328_),
    .A2(_04341_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20005_ (.A1(_08389_),
    .A2(_08390_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20006_ (.A1(_08632_),
    .A2(_08636_),
    .B(_04327_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20007_ (.A1(_04343_),
    .A2(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20008_ (.A1(_08628_),
    .A2(_08666_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20009_ (.A1(_08383_),
    .A2(_04346_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20010_ (.A1(_04345_),
    .A2(_04347_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20011_ (.A1(net3382),
    .A2(_08654_),
    .A3(_08655_),
    .Z(_04349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20012_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_08361_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20013_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .A2(_04350_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20014_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(net60),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20015_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_04352_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20016_ (.A1(_08370_),
    .A2(_04349_),
    .A3(_04351_),
    .A4(_04353_),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20017_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20018_ (.A1(_08360_),
    .A2(_04327_),
    .Z(_04356_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _20019_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_08658_),
    .A3(_04356_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20020_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_04355_),
    .B(_04357_),
    .C(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _20021_ (.A1(_08660_),
    .A2(_04348_),
    .A3(_04354_),
    .A4(_04358_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20022_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_08871_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20023_ (.A1(_08640_),
    .A2(net3354),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20024_ (.A1(_08389_),
    .A2(_08362_),
    .Z(_04362_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20025_ (.A1(_02019_),
    .A2(_04361_),
    .A3(_04362_),
    .A4(_04356_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20026_ (.A1(_04342_),
    .A2(_04359_),
    .B(_04360_),
    .C(_04363_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20027_ (.A1(_08624_),
    .A2(_04338_),
    .A3(_04339_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20028_ (.A1(_04362_),
    .A2(_04356_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20029_ (.A1(_08370_),
    .A2(_04349_),
    .A3(_04352_),
    .Z(_04366_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20030_ (.A1(_08389_),
    .A2(_04366_),
    .B(_04351_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20031_ (.A1(_04361_),
    .A2(_04365_),
    .B(_04367_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20032_ (.A1(_08383_),
    .A2(_04345_),
    .A3(_04346_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20033_ (.A1(_02019_),
    .A2(_04361_),
    .B(_08360_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20034_ (.A1(_08624_),
    .A2(_04328_),
    .A3(_04370_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _20035_ (.A1(_04364_),
    .A2(_04368_),
    .A3(_04369_),
    .A4(_04371_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20036_ (.A1(_08628_),
    .A2(_08637_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20037_ (.A1(_08871_),
    .A2(_04350_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20038_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_08658_),
    .B1(_04362_),
    .B2(_04327_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20039_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_04374_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20040_ (.A1(_04348_),
    .A2(_04372_),
    .B1(_04373_),
    .B2(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .C(_04375_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20041_ (.A1(_04328_),
    .A2(_04340_),
    .B(_08624_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20042_ (.A1(_04376_),
    .A2(_04377_),
    .B(_04360_),
    .C(_04354_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20043_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_08632_),
    .A3(_08636_),
    .Z(_04378_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20044_ (.A1(_08360_),
    .A2(_04372_),
    .B1(_04378_),
    .B2(_04327_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20045_ (.A1(_04362_),
    .A2(_04379_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20046_ (.A1(_08363_),
    .A2(_04328_),
    .A3(_04340_),
    .B(_04380_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20047_ (.A1(_08389_),
    .A2(_04352_),
    .B(_08681_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _20048_ (.A1(_08385_),
    .A2(_02380_),
    .A3(_04346_),
    .B1(_04381_),
    .B2(\cs_registers_i.debug_mode_i ),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20049_ (.I(_04382_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20050_ (.A1(net145),
    .A2(_08642_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20051_ (.A1(net3473),
    .A2(_06411_),
    .A3(_06205_),
    .A4(_06244_),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20052_ (.A1(_06720_),
    .A2(_04384_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20053_ (.A1(_08384_),
    .A2(_04385_),
    .A3(_08665_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output186 (.I(net186),
    .Z(data_wdata_o[0]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output185 (.I(net185),
    .Z(data_req_o));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output184 (.I(net184),
    .Z(data_be_o[3]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20057_ (.A1(_08638_),
    .A2(_04383_),
    .B(_04386_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20058_ (.A1(_08880_),
    .A2(_06782_),
    .A3(_08396_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20059_ (.A1(_08404_),
    .A2(_01967_),
    .A3(_04390_),
    .Z(_04391_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _20060_ (.A1(_06994_),
    .A2(net3091),
    .A3(_01958_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20061_ (.A1(_08880_),
    .A2(_01968_),
    .A3(_04392_),
    .B(_01960_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20062_ (.A1(_06246_),
    .A2(_04391_),
    .B(_04393_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20063_ (.I0(net334),
    .I1(\alu_adder_result_ex[0] ),
    .S(net3292),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20064_ (.I0(\ex_block_i.alu_i.imd_val_q_i[0] ),
    .I1(_04394_),
    .S(_08411_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output183 (.I(net183),
    .Z(data_be_o[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20066_ (.I0(net151),
    .I1(net425),
    .S(_08462_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20067_ (.I0(\ex_block_i.alu_i.imd_val_q_i[10] ),
    .I1(_04396_),
    .S(_08411_),
    .Z(_01513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20068_ (.I0(net152),
    .I1(net422),
    .S(_08462_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20069_ (.I0(\ex_block_i.alu_i.imd_val_q_i[11] ),
    .I1(_04397_),
    .S(_08411_),
    .Z(_01514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20070_ (.I0(net153),
    .I1(net420),
    .S(_08462_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20071_ (.I0(\ex_block_i.alu_i.imd_val_q_i[12] ),
    .I1(_04398_),
    .S(_08411_),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20072_ (.I0(net154),
    .I1(net424),
    .S(_08462_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20073_ (.I0(\ex_block_i.alu_i.imd_val_q_i[13] ),
    .I1(_04399_),
    .S(_08411_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20074_ (.I0(net364),
    .I1(_07449_),
    .S(_08462_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20075_ (.I0(\ex_block_i.alu_i.imd_val_q_i[14] ),
    .I1(_04400_),
    .S(_08411_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20076_ (.I0(net156),
    .I1(_07486_),
    .S(_08462_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20077_ (.I0(\ex_block_i.alu_i.imd_val_q_i[15] ),
    .I1(_04401_),
    .S(_08411_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20078_ (.I0(net402),
    .I1(_07544_),
    .S(_08462_),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20079_ (.I0(\ex_block_i.alu_i.imd_val_q_i[16] ),
    .I1(_04402_),
    .S(_08411_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20080_ (.I0(net158),
    .I1(_07582_),
    .S(_08462_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20081_ (.I0(\ex_block_i.alu_i.imd_val_q_i[17] ),
    .I1(_04403_),
    .S(_08411_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20082_ (.I0(net361),
    .I1(net414),
    .S(_08462_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output182 (.I(net182),
    .Z(data_be_o[1]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20084_ (.I0(\ex_block_i.alu_i.imd_val_q_i[18] ),
    .I1(_04404_),
    .S(_08411_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20085_ (.I0(net160),
    .I1(net441),
    .S(_08462_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20086_ (.I0(\ex_block_i.alu_i.imd_val_q_i[19] ),
    .I1(_04406_),
    .S(_08411_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20087_ (.I0(net276),
    .I1(\alu_adder_result_ex[1] ),
    .S(net3292),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20088_ (.I0(\ex_block_i.alu_i.imd_val_q_i[1] ),
    .I1(_04407_),
    .S(_08411_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 output181 (.I(net181),
    .Z(data_be_o[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20090_ (.I0(net161),
    .I1(net410),
    .S(_08462_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20091_ (.I0(\ex_block_i.alu_i.imd_val_q_i[20] ),
    .I1(_04409_),
    .S(_08411_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20092_ (.I0(net162),
    .I1(net442),
    .S(_08462_),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20093_ (.I0(\ex_block_i.alu_i.imd_val_q_i[21] ),
    .I1(_04410_),
    .S(_08411_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20094_ (.I0(net163),
    .I1(_07838_),
    .S(_08462_),
    .Z(_04411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20095_ (.I0(\ex_block_i.alu_i.imd_val_q_i[22] ),
    .I1(_04411_),
    .S(_08411_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20096_ (.I0(net372),
    .I1(_07875_),
    .S(_08462_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20097_ (.I0(\ex_block_i.alu_i.imd_val_q_i[23] ),
    .I1(_04412_),
    .S(_08411_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20098_ (.I0(net376),
    .I1(_07936_),
    .S(_08462_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20099_ (.I0(\ex_block_i.alu_i.imd_val_q_i[24] ),
    .I1(_04413_),
    .S(_08411_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20100_ (.I0(net289),
    .I1(_07973_),
    .S(_08462_),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20101_ (.I0(\ex_block_i.alu_i.imd_val_q_i[25] ),
    .I1(_04414_),
    .S(_08411_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20102_ (.I0(net167),
    .I1(_08017_),
    .S(_08462_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20103_ (.I0(\ex_block_i.alu_i.imd_val_q_i[26] ),
    .I1(_04415_),
    .S(_08411_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20104_ (.I0(net366),
    .I1(_08055_),
    .S(_08462_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output180 (.I(net180),
    .Z(data_addr_o[9]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20106_ (.I0(\ex_block_i.alu_i.imd_val_q_i[27] ),
    .I1(_04416_),
    .S(_08411_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20107_ (.I0(net169),
    .I1(net530),
    .S(_08462_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20108_ (.I0(\ex_block_i.alu_i.imd_val_q_i[28] ),
    .I1(_04418_),
    .S(_08411_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20109_ (.I0(net337),
    .I1(_08145_),
    .S(_08462_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20110_ (.I0(\ex_block_i.alu_i.imd_val_q_i[29] ),
    .I1(_04419_),
    .S(_08411_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20111_ (.I0(net171),
    .I1(net557),
    .S(_08462_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20112_ (.I0(\ex_block_i.alu_i.imd_val_q_i[2] ),
    .I1(_04420_),
    .S(_08411_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20113_ (.I0(net258),
    .I1(_08193_),
    .S(_08462_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20114_ (.I0(\ex_block_i.alu_i.imd_val_q_i[30] ),
    .I1(_04421_),
    .S(_08411_),
    .Z(_01535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20115_ (.A1(net279),
    .A2(_08461_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20116_ (.A1(net432),
    .A2(_04422_),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20117_ (.I0(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .I1(_04423_),
    .S(_08411_),
    .Z(_01536_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20118_ (.A1(_11171_[0]),
    .A2(_02984_),
    .B(_08459_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output179 (.I(net179),
    .Z(data_addr_o[8]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20120_ (.I0(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .I1(\alu_adder_result_ex[0] ),
    .S(_02981_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20121_ (.A1(_08456_),
    .A2(_04426_),
    .B(net3656),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output178 (.I(net178),
    .Z(data_addr_o[7]));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20123_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_11172_[0]),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20124_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_11172_[0]),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20125_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_11172_[0]),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20126_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_11172_[0]),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20127_ (.I0(_04429_),
    .I1(_04430_),
    .I2(_04431_),
    .I3(_04432_),
    .S0(_02912_),
    .S1(_02915_),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20128_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_11172_[0]),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20129_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_11172_[0]),
    .Z(_04435_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20130_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_11172_[0]),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20131_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_11172_[0]),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20132_ (.I0(_04434_),
    .I1(_04435_),
    .I2(_04436_),
    .I3(_04437_),
    .S0(_02912_),
    .S1(_02915_),
    .Z(_04438_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20133_ (.A1(_08401_),
    .A2(_02917_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20134_ (.I0(_04433_),
    .I1(_04438_),
    .S(_04439_),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20135_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .A2(_04440_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output177 (.I(net177),
    .Z(data_addr_o[6]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20137_ (.A1(_02906_),
    .A2(_08452_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20138_ (.A1(net3658),
    .A2(\alu_adder_result_ex[0] ),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .C(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20139_ (.A1(_04424_),
    .A2(_04427_),
    .B(_04441_),
    .C(_04444_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _20140_ (.A1(net3658),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A3(_07017_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20141_ (.A1(_06744_),
    .A2(_02906_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20142_ (.A1(_04446_),
    .A2(_04447_),
    .Z(_04448_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20143_ (.A1(net3647),
    .A2(_04448_),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20144_ (.A1(_07025_),
    .A2(_04449_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20145_ (.I0(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .I1(_11184_[0]),
    .S(_03152_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20146_ (.A1(net3647),
    .A2(_04451_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20147_ (.A1(net3371),
    .A2(_04445_),
    .A3(_04450_),
    .A4(_04452_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20148_ (.A1(net3371),
    .A2(_08405_),
    .A3(_08468_),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output176 (.I(net176),
    .Z(data_addr_o[5]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output175 (.I(net175),
    .Z(data_addr_o[4]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20151_ (.I0(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .I1(_04453_),
    .S(_04454_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20152_ (.A1(_06744_),
    .A2(_02906_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 output174 (.I(net174),
    .Z(data_addr_o[3]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20154_ (.I0(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .I1(\alu_adder_result_ex[1] ),
    .S(_02981_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20155_ (.A1(_04457_),
    .A2(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output173 (.I(net295),
    .Z(data_addr_o[31]));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20157_ (.A1(_08403_),
    .A2(_03022_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output172 (.I(net257),
    .Z(data_addr_o[30]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20159_ (.A1(net3647),
    .A2(_08452_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20160_ (.A1(net3658),
    .A2(\alu_adder_result_ex[1] ),
    .B1(_04426_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04464_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20161_ (.A1(_07016_),
    .A2(_04460_),
    .A3(_04462_),
    .B(_04465_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20162_ (.A1(_06935_),
    .A2(_04449_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20163_ (.I0(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .I1(_11187_[0]),
    .S(_03152_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20164_ (.A1(net3647),
    .A2(_04468_),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20165_ (.A1(net3371),
    .A2(_04466_),
    .A3(_04467_),
    .A4(_04469_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20166_ (.I0(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .I1(_04470_),
    .S(_04454_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20167_ (.A1(_11175_[0]),
    .A2(_02984_),
    .B(_08459_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20168_ (.I0(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .I1(net171),
    .S(_02981_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20169_ (.A1(_08456_),
    .A2(_04472_),
    .B(net3656),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output171 (.I(net171),
    .Z(data_addr_o[2]));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20171_ (.A1(net3658),
    .A2(net171),
    .B1(_04459_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04443_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20172_ (.A1(_04471_),
    .A2(_04473_),
    .B(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20173_ (.I0(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .I1(_11189_[0]),
    .S(_03152_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20174_ (.A1(_02906_),
    .A2(_04477_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20175_ (.A1(_04446_),
    .A2(_04447_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20176_ (.A1(net3372),
    .A2(_03512_),
    .A3(_04479_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20177_ (.A1(net3371),
    .A2(_04476_),
    .A3(_04478_),
    .A4(_04480_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20178_ (.I0(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .I1(_04481_),
    .S(_04454_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _20179_ (.A1(_08469_),
    .A2(_03545_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20180_ (.A1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A2(_03545_),
    .B1(_04482_),
    .B2(_11197_[0]),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20181_ (.A1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A2(_08469_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output170 (.I(net170),
    .Z(data_addr_o[29]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output169 (.I(net169),
    .Z(data_addr_o[28]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20184_ (.I0(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .I1(net174),
    .S(_02981_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20185_ (.A1(_04457_),
    .A2(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output168 (.I(net168),
    .Z(data_addr_o[27]));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20187_ (.A1(_11179_[0]),
    .A2(_02984_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output167 (.I(net167),
    .Z(data_addr_o[26]));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20189_ (.A1(net3658),
    .A2(net174),
    .B1(_04472_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04446_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20190_ (.A1(_07016_),
    .A2(_04488_),
    .A3(_04490_),
    .B(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20191_ (.A1(net3647),
    .A2(_04454_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20192_ (.I(_04494_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20193_ (.A1(net3369),
    .A2(_04479_),
    .B(_04493_),
    .C(_04495_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20194_ (.A1(net3647),
    .A2(_04483_),
    .B(_04484_),
    .C(_04496_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20195_ (.I0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .I1(net175),
    .S(_02981_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20196_ (.A1(_04457_),
    .A2(_04497_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20197_ (.A1(_11171_[0]),
    .A2(_03060_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20198_ (.A1(net3658),
    .A2(net175),
    .B1(_04487_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04464_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20199_ (.A1(_07016_),
    .A2(_04498_),
    .A3(_04499_),
    .B(_04500_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20200_ (.A1(_07106_),
    .A2(_04449_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20201_ (.I0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .I1(_11201_[0]),
    .S(_03152_),
    .Z(_04503_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20202_ (.A1(net3647),
    .A2(_04503_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20203_ (.A1(net3371),
    .A2(_04501_),
    .A3(_04502_),
    .A4(_04504_),
    .Z(_04505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20204_ (.I0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .I1(_04505_),
    .S(_04454_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20205_ (.I0(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .I1(net176),
    .S(_02981_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20206_ (.A1(_04457_),
    .A2(_04506_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20207_ (.A1(_11177_[0]),
    .A2(_03060_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20208_ (.A1(net3658),
    .A2(net176),
    .B1(_04497_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04464_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20209_ (.A1(_07016_),
    .A2(_04507_),
    .A3(_04508_),
    .B(_04509_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20210_ (.A1(net3367),
    .A2(_04449_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20211_ (.I0(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .I1(_11210_[0]),
    .S(_03152_),
    .Z(_04512_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20212_ (.A1(net3647),
    .A2(_04512_),
    .Z(_04513_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20213_ (.A1(net3371),
    .A2(_04510_),
    .A3(_04511_),
    .A4(_04513_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20214_ (.I0(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .I1(_04514_),
    .S(_04454_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20215_ (.I0(net436),
    .I1(net174),
    .S(net3292),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20216_ (.I0(\ex_block_i.alu_i.imd_val_q_i[3] ),
    .I1(_04515_),
    .S(_08411_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20217_ (.A1(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A2(_03545_),
    .B1(_04482_),
    .B2(_11221_[0]),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20218_ (.A1(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A2(_08469_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20219_ (.I0(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .I1(net177),
    .S(_02981_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20220_ (.A1(_04457_),
    .A2(_04518_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20221_ (.A1(_11175_[0]),
    .A2(_03060_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20222_ (.A1(net3658),
    .A2(net177),
    .B1(_04506_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04446_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20223_ (.A1(_07016_),
    .A2(_04519_),
    .A3(_04520_),
    .B(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output166 (.I(net166),
    .Z(data_addr_o[25]));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20225_ (.A1(net3366),
    .A2(_04448_),
    .B(_04494_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20226_ (.A1(_04522_),
    .A2(_04524_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20227_ (.A1(net3647),
    .A2(_04516_),
    .B(_04517_),
    .C(_04525_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20228_ (.I0(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .I1(net178),
    .S(_02981_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20229_ (.A1(_11179_[0]),
    .A2(_03060_),
    .Z(_04527_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20230_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .A2(_08459_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20231_ (.A1(_08456_),
    .A2(_04526_),
    .B1(_04527_),
    .B2(_04528_),
    .C(net3656),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20232_ (.A1(net3658),
    .A2(net178),
    .B1(_04518_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04446_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20233_ (.A1(net3365),
    .A2(_04448_),
    .B1(_04529_),
    .B2(_04530_),
    .C(_04494_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20234_ (.A1(_09860_[0]),
    .A2(_02906_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20235_ (.I0(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .I1(_04532_),
    .S(_04482_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20236_ (.A1(_04531_),
    .A2(_04533_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20237_ (.A1(_11171_[0]),
    .A2(_02990_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20238_ (.I0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .I1(net179),
    .S(_02981_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20239_ (.A1(_08456_),
    .A2(_04535_),
    .B(net3656),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20240_ (.A1(net3658),
    .A2(net179),
    .B1(_04526_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04464_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20241_ (.A1(_04534_),
    .A2(_04536_),
    .B(_04537_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20242_ (.A1(net3364),
    .A2(_04449_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20243_ (.I0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .I1(_03151_),
    .S(_03152_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20244_ (.A1(net3647),
    .A2(_04540_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20245_ (.A1(net3371),
    .A2(_04538_),
    .A3(_04539_),
    .A4(_04541_),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20246_ (.I0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .I1(_04542_),
    .S(_04454_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20247_ (.I0(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .I1(net180),
    .S(_02981_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20248_ (.A1(_04457_),
    .A2(_04543_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20249_ (.A1(_11177_[0]),
    .A2(_02990_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20250_ (.A1(net3658),
    .A2(net180),
    .B1(_04535_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04464_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20251_ (.A1(_07016_),
    .A2(_04544_),
    .A3(_04545_),
    .B(_04546_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20252_ (.A1(net3363),
    .A2(_04449_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20253_ (.I0(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .I1(_03310_),
    .S(_03152_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20254_ (.A1(net3647),
    .A2(_04549_),
    .Z(_04550_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20255_ (.A1(net3371),
    .A2(_04547_),
    .A3(_04548_),
    .A4(_04550_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output165 (.I(net165),
    .Z(data_addr_o[24]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20257_ (.I0(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .I1(_04551_),
    .S(_04454_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20258_ (.I0(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .I1(net151),
    .S(_02981_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20259_ (.A1(_04457_),
    .A2(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20260_ (.A1(_11175_[0]),
    .A2(_02990_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20261_ (.A1(_07016_),
    .A2(_04554_),
    .A3(_04555_),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20262_ (.A1(net3658),
    .A2(net151),
    .B1(_04543_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04446_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20263_ (.A1(net3362),
    .A2(_04448_),
    .B1(_04556_),
    .B2(_04557_),
    .C(_04494_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output164 (.I(net164),
    .Z(data_addr_o[23]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20265_ (.A1(_03512_),
    .A2(_03339_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20266_ (.I0(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .I1(_04560_),
    .S(_04482_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20267_ (.A1(_04558_),
    .A2(_04561_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20268_ (.A1(_11179_[0]),
    .A2(_02990_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20269_ (.I0(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .I1(net152),
    .S(_02981_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20270_ (.A1(_04457_),
    .A2(_04563_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20271_ (.A1(_04457_),
    .A2(_04562_),
    .B(_04564_),
    .C(_07016_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20272_ (.A1(net3658),
    .A2(net152),
    .B1(_04553_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C(_04446_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20273_ (.A1(net3377),
    .A2(_04448_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20274_ (.A1(_04566_),
    .A2(_04567_),
    .B(_02906_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20275_ (.A1(_04565_),
    .A2(_04568_),
    .B(_03398_),
    .C(_04454_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20276_ (.A1(_07282_),
    .A2(_04454_),
    .B(_04569_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20277_ (.A1(net3381),
    .A2(_04448_),
    .B(net3417),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20278_ (.I0(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .I1(net153),
    .S(_02981_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20279_ (.A1(_04457_),
    .A2(_04571_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20280_ (.A1(_11171_[0]),
    .A2(_02998_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20281_ (.A1(net3658),
    .A2(net153),
    .B1(_04563_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20282_ (.A1(_07016_),
    .A2(_04572_),
    .A3(_04573_),
    .B(_04574_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20283_ (.A1(_04570_),
    .A2(_04575_),
    .B(_03418_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20284_ (.A1(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .A2(_04454_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20285_ (.A1(_04454_),
    .A2(_04576_),
    .B(_04577_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20286_ (.A1(_08469_),
    .A2(_03545_),
    .A3(_03459_),
    .Z(_04578_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20287_ (.A1(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .A2(_03152_),
    .B(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20288_ (.I0(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .I1(net154),
    .S(_02981_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20289_ (.A1(_04457_),
    .A2(_04580_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20290_ (.A1(_11177_[0]),
    .A2(_02998_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20291_ (.A1(net3658),
    .A2(net154),
    .B1(_04571_),
    .B2(net3654),
    .C(_04464_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20292_ (.A1(_07016_),
    .A2(_04581_),
    .A3(_04582_),
    .B(_04583_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20293_ (.A1(_08469_),
    .A2(_04584_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20294_ (.A1(net3647),
    .A2(_04448_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20295_ (.A1(net3361),
    .A2(_04586_),
    .B(net3373),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20296_ (.I0(_04587_),
    .I1(_07372_),
    .S(_08469_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20297_ (.A1(net3417),
    .A2(_04579_),
    .B(_04585_),
    .C(_04588_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20298_ (.I0(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .I1(net365),
    .S(_02981_),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20299_ (.A1(_04457_),
    .A2(_04589_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20300_ (.A1(_11175_[0]),
    .A2(_02998_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20301_ (.A1(net3658),
    .A2(net365),
    .B1(_04580_),
    .B2(net3654),
    .C(_04443_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20302_ (.A1(_07016_),
    .A2(_04590_),
    .A3(_04591_),
    .B(_04592_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20303_ (.A1(_02906_),
    .A2(_04448_),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20304_ (.A1(net3351),
    .A2(_04594_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20305_ (.A1(net3371),
    .A2(_03498_),
    .A3(_04593_),
    .A4(_04595_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20306_ (.I0(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .I1(_04596_),
    .S(_04454_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20307_ (.I0(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .I1(net156),
    .S(_02981_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20308_ (.A1(_04457_),
    .A2(_04597_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20309_ (.A1(_11179_[0]),
    .A2(_02998_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20310_ (.A1(net3658),
    .A2(net156),
    .B1(_04589_),
    .B2(net3654),
    .C(_04443_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20311_ (.A1(_07016_),
    .A2(_04598_),
    .A3(_04599_),
    .B(_04600_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20312_ (.A1(_08812_),
    .A2(_04594_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20313_ (.A1(_03526_),
    .A2(_04601_),
    .A3(_04602_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20314_ (.I0(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .I1(_04603_),
    .S(_04454_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20315_ (.I0(net175),
    .I1(net331),
    .S(_08462_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20316_ (.I0(\ex_block_i.alu_i.imd_val_q_i[4] ),
    .I1(_04604_),
    .S(_08411_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20317_ (.I0(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .I1(net404),
    .S(_02981_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20318_ (.A1(_04457_),
    .A2(_04605_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20319_ (.A1(_11171_[0]),
    .A2(_03010_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20320_ (.A1(net3658),
    .A2(net404),
    .B1(_04597_),
    .B2(net3654),
    .C(_04443_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20321_ (.A1(_07016_),
    .A2(_04606_),
    .A3(_04607_),
    .B(_04608_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20322_ (.A1(_07526_),
    .A2(_04594_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20323_ (.A1(_03556_),
    .A2(_04609_),
    .A3(_04610_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20324_ (.I0(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .I1(_04611_),
    .S(_04454_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20325_ (.I0(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .I1(net158),
    .S(_02981_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20326_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(_08403_),
    .A3(_02981_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _20327_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .A2(_04447_),
    .A3(_04613_),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20328_ (.A1(_08456_),
    .A2(_04612_),
    .B(_04614_),
    .C(net3656),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20329_ (.A1(net3658),
    .A2(net158),
    .B1(_04605_),
    .B2(net3654),
    .C(_04443_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20330_ (.I(_03580_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20331_ (.A1(net3349),
    .A2(_04594_),
    .B1(_04615_),
    .B2(_04616_),
    .C(_04617_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20332_ (.I0(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .I1(_04618_),
    .S(_04454_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20333_ (.I0(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .I1(net361),
    .S(_02981_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20334_ (.A1(_04457_),
    .A2(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20335_ (.A1(_11175_[0]),
    .A2(_03010_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20336_ (.A1(net3658),
    .A2(net361),
    .B1(_04612_),
    .B2(net3654),
    .C(_04443_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20337_ (.A1(_07016_),
    .A2(_04620_),
    .A3(_04621_),
    .B(_04622_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20338_ (.A1(_08823_),
    .A2(_04594_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20339_ (.A1(net3371),
    .A2(_03642_),
    .A3(_04623_),
    .A4(_04624_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20340_ (.I0(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .I1(_04625_),
    .S(_04454_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20341_ (.A1(_11179_[0]),
    .A2(_03010_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20342_ (.I0(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .I1(net160),
    .S(_02981_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20343_ (.A1(_04457_),
    .A2(_04627_),
    .B(net3656),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20344_ (.A1(net3658),
    .A2(net160),
    .B1(_04619_),
    .B2(net3654),
    .C(_04443_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20345_ (.A1(_04626_),
    .A2(_04628_),
    .B(_04629_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20346_ (.A1(net3348),
    .A2(_04594_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20347_ (.A1(net3371),
    .A2(_03666_),
    .A3(_04630_),
    .A4(_04631_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20348_ (.I0(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .I1(_04632_),
    .S(_04454_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20349_ (.I0(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .I1(net161),
    .S(_02981_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20350_ (.A1(_11171_[0]),
    .A2(_03026_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _20351_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .A2(_04447_),
    .A3(_04634_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20352_ (.A1(_08456_),
    .A2(_04633_),
    .B(_04635_),
    .C(net3656),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20353_ (.A1(net3658),
    .A2(net161),
    .B1(_04627_),
    .B2(net3654),
    .C(_04443_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20354_ (.A1(net3371),
    .A2(_03691_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20355_ (.A1(_07712_),
    .A2(_04594_),
    .B1(_04636_),
    .B2(_04637_),
    .C(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20356_ (.I0(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .I1(_04639_),
    .S(_04454_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20357_ (.I0(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .I1(net162),
    .S(_02981_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20358_ (.A1(_04457_),
    .A2(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20359_ (.A1(_11177_[0]),
    .A2(_03026_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20360_ (.A1(net3658),
    .A2(net162),
    .B1(_04633_),
    .B2(net3654),
    .C(_04443_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20361_ (.A1(_07016_),
    .A2(_04641_),
    .A3(_04642_),
    .B(_04643_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20362_ (.A1(net3347),
    .A2(_04594_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20363_ (.A1(_03705_),
    .A2(_04644_),
    .A3(_04645_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20364_ (.I0(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .I1(_04646_),
    .S(_04454_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20365_ (.A1(_11175_[0]),
    .A2(_03026_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20366_ (.I0(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .I1(net163),
    .S(_02981_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20367_ (.A1(_04457_),
    .A2(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20368_ (.A1(_04457_),
    .A2(_04647_),
    .B(_04649_),
    .C(_07016_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20369_ (.A1(net3658),
    .A2(net163),
    .B1(_04640_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20370_ (.A1(net3346),
    .A2(_04448_),
    .B(_04651_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20371_ (.A1(_04494_),
    .A2(_04650_),
    .A3(_04652_),
    .Z(_04653_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20372_ (.A1(net3373),
    .A2(_03735_),
    .Z(_04654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20373_ (.I0(_04654_),
    .I1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .S(_08469_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20374_ (.A1(_04653_),
    .A2(_04655_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20375_ (.I0(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .I1(net372),
    .S(_02981_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20376_ (.A1(_11179_[0]),
    .A2(_03026_),
    .Z(_04657_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _20377_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .A2(_04447_),
    .A3(_04657_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20378_ (.A1(_08456_),
    .A2(_04656_),
    .B(_04658_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20379_ (.A1(net3656),
    .A2(_02906_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20380_ (.A1(net3345),
    .A2(_04448_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20381_ (.A1(net3658),
    .A2(net372),
    .B1(_04648_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20382_ (.A1(_03512_),
    .A2(_04661_),
    .A3(_04662_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20383_ (.A1(_02906_),
    .A2(net3092),
    .B1(_04659_),
    .B2(_04660_),
    .C(_04663_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20384_ (.I0(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .I1(_04664_),
    .S(_04454_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20385_ (.A1(net3658),
    .A2(net377),
    .B1(_04656_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20386_ (.I0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .I1(net377),
    .S(_02981_),
    .Z(_04666_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20387_ (.A1(_11171_[0]),
    .A2(_03036_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20388_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .A2(_08459_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20389_ (.A1(_08456_),
    .A2(_04666_),
    .B1(_04667_),
    .B2(_04668_),
    .C(net3656),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20390_ (.A1(net3344),
    .A2(_04448_),
    .B1(_04665_),
    .B2(_04669_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20391_ (.I0(_03769_),
    .I1(_04670_),
    .S(_02906_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20392_ (.I0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .I1(_04671_),
    .S(_04454_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20393_ (.A1(net3343),
    .A2(_04448_),
    .Z(_04672_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20394_ (.A1(net3658),
    .A2(net289),
    .B1(_04666_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20395_ (.I0(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .I1(net289),
    .S(_02981_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20396_ (.A1(_11177_[0]),
    .A2(_03036_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20397_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .A2(_08459_),
    .Z(_04676_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20398_ (.A1(_08456_),
    .A2(_04674_),
    .B1(_04675_),
    .B2(_04676_),
    .C(net3656),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20399_ (.A1(_04673_),
    .A2(_04677_),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20400_ (.A1(_02906_),
    .A2(net3075),
    .Z(_04679_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20401_ (.A1(_03512_),
    .A2(_04672_),
    .A3(_04678_),
    .B(_04679_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20402_ (.I0(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .I1(_04680_),
    .S(_04454_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20403_ (.I0(net341),
    .I1(net176),
    .S(net3292),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20404_ (.I0(\ex_block_i.alu_i.imd_val_q_i[5] ),
    .I1(_04681_),
    .S(_08411_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20405_ (.A1(_11175_[0]),
    .A2(_03036_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20406_ (.I0(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .I1(net167),
    .S(_02981_),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20407_ (.A1(_04457_),
    .A2(_04683_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20408_ (.A1(_04457_),
    .A2(_04682_),
    .B(_04684_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20409_ (.A1(net3658),
    .A2(net167),
    .B1(_04674_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20410_ (.A1(net3342),
    .A2(_04448_),
    .B(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20411_ (.A1(net3656),
    .A2(_04685_),
    .B(_04687_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20412_ (.I(_08470_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20413_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(_08469_),
    .B1(_04689_),
    .B2(net3087),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20414_ (.A1(_04494_),
    .A2(_04688_),
    .B(_04690_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20415_ (.A1(_11179_[0]),
    .A2(_03036_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20416_ (.I0(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .I1(net368),
    .S(_02981_),
    .Z(_04692_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20417_ (.A1(_08456_),
    .A2(_04692_),
    .B(net3656),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20418_ (.A1(net3658),
    .A2(net368),
    .B1(_04683_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20419_ (.A1(_04691_),
    .A2(_04693_),
    .B(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20420_ (.A1(net3357),
    .A2(_04448_),
    .B(_03512_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20421_ (.I(_04454_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20422_ (.A1(_03512_),
    .A2(net3079),
    .B1(_04695_),
    .B2(_04696_),
    .C(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20423_ (.A1(_08041_),
    .A2(_08469_),
    .B(_04698_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20424_ (.A1(_03512_),
    .A2(net3062),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20425_ (.A1(net3341),
    .A2(_04448_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20426_ (.A1(net3658),
    .A2(net169),
    .B1(_04692_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20427_ (.I0(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .I1(net169),
    .S(_02981_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20428_ (.A1(_04457_),
    .A2(_04702_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20429_ (.A1(_11171_[0]),
    .A2(_03046_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _20430_ (.A1(_03512_),
    .A2(_04700_),
    .A3(_04701_),
    .B1(_04703_),
    .B2(_04704_),
    .B3(_04660_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20431_ (.A1(_04699_),
    .A2(_04705_),
    .Z(_04706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20432_ (.I0(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .I1(_04706_),
    .S(_04454_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20433_ (.I0(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .I1(net339),
    .S(_02981_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20434_ (.A1(_04457_),
    .A2(_04707_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20435_ (.A1(_11177_[0]),
    .A2(_03046_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20436_ (.A1(net3658),
    .A2(net339),
    .B1(_04702_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20437_ (.A1(net3340),
    .A2(_04448_),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _20438_ (.A1(_07016_),
    .A2(_04708_),
    .A3(_04709_),
    .B1(_04710_),
    .B2(_04711_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20439_ (.I0(net3074),
    .I1(_04712_),
    .S(_02906_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20440_ (.I0(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .I1(_04713_),
    .S(_04454_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20441_ (.I0(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .I1(net257),
    .S(_02981_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20442_ (.A1(_04457_),
    .A2(_04714_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20443_ (.A1(_11175_[0]),
    .A2(_03046_),
    .B(_04447_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20444_ (.A1(net3658),
    .A2(net257),
    .B1(_04707_),
    .B2(net3654),
    .C(_04446_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20445_ (.A1(net3339),
    .A2(_04448_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _20446_ (.A1(_07016_),
    .A2(_04715_),
    .A3(_04716_),
    .B1(_04717_),
    .B2(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20447_ (.I0(net3073),
    .I1(_04719_),
    .S(_02906_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20448_ (.I0(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .I1(_04720_),
    .S(_04454_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20449_ (.A1(net3656),
    .A2(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A3(_04447_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20450_ (.A1(net3658),
    .A2(_04721_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20451_ (.A1(net3656),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .A3(_04457_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20452_ (.A1(net3094),
    .A2(_04722_),
    .B(_04723_),
    .C(_08452_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20453_ (.A1(net3656),
    .A2(_11179_[0]),
    .A3(_04457_),
    .A4(_03046_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20454_ (.A1(net3654),
    .A2(_04714_),
    .B(_04724_),
    .C(_04725_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20455_ (.A1(_08235_),
    .A2(_04448_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20456_ (.A1(_03512_),
    .A2(net3061),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20457_ (.A1(_03512_),
    .A2(_04726_),
    .A3(_04727_),
    .B(_04728_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20458_ (.I0(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .I1(_04729_),
    .S(_04454_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20459_ (.A1(_11373_[0]),
    .A2(net3086),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20460_ (.A1(_03980_),
    .A2(_04730_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20461_ (.A1(_11379_[0]),
    .A2(_04731_),
    .B(_11378_[0]),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20462_ (.A1(_11387_[0]),
    .A2(_04732_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20463_ (.A1(_03512_),
    .A2(_03152_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20464_ (.A1(net3654),
    .A2(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A3(net173),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20465_ (.A1(_04446_),
    .A2(_04457_),
    .B(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20466_ (.A1(_04733_),
    .A2(_04734_),
    .B1(_04736_),
    .B2(_03512_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20467_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .I1(_04737_),
    .S(_04454_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20468_ (.A1(net3204),
    .A2(_10978_[0]),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20469_ (.A1(_10980_[0]),
    .A2(_10972_[0]),
    .A3(_04738_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20470_ (.A1(_10913_[0]),
    .A2(_11383_[0]),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20471_ (.A1(_10992_[0]),
    .A2(_10995_[0]),
    .A3(_04740_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20472_ (.A1(_10983_[0]),
    .A2(_10985_[0]),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20473_ (.A1(_10976_[0]),
    .A2(net3217),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20474_ (.A1(_10989_[0]),
    .A2(_10914_[0]),
    .A3(_11381_[0]),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20475_ (.A1(_04742_),
    .A2(_04743_),
    .A3(_04744_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20476_ (.A1(_04739_),
    .A2(_04741_),
    .A3(_04745_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20477_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .A2(net3303),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20478_ (.A1(_08589_),
    .A2(_04747_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20479_ (.A1(_04746_),
    .A2(_04748_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20480_ (.A1(net3233),
    .A2(net3229),
    .A3(_04749_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20481_ (.A1(_03932_),
    .A2(net3078),
    .B(_03980_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20482_ (.A1(_11379_[0]),
    .A2(_11387_[0]),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20483_ (.A1(_11387_[0]),
    .A2(_11378_[0]),
    .B1(_04751_),
    .B2(_04752_),
    .C(_11386_[0]),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20484_ (.A1(_04750_),
    .A2(_04753_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20485_ (.A1(_08452_),
    .A2(_04447_),
    .B1(_04734_),
    .B2(_04754_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20486_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .I1(_04755_),
    .S(_04454_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20487_ (.I0(net177),
    .I1(_08275_),
    .S(_08462_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20488_ (.I0(\ex_block_i.alu_i.imd_val_q_i[6] ),
    .I1(_04756_),
    .S(_08411_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20489_ (.I0(net178),
    .I1(net426),
    .S(_08462_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20490_ (.I0(\ex_block_i.alu_i.imd_val_q_i[7] ),
    .I1(_04757_),
    .S(_08411_),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20491_ (.I0(net179),
    .I1(net412),
    .S(_08462_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20492_ (.I0(\ex_block_i.alu_i.imd_val_q_i[8] ),
    .I1(_04758_),
    .S(_08411_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20493_ (.I0(net180),
    .I1(net408),
    .S(_08462_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20494_ (.I0(\ex_block_i.alu_i.imd_val_q_i[9] ),
    .I1(_04759_),
    .S(_08411_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20495_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .A2(net3221),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20496_ (.A1(_08370_),
    .A2(_08629_),
    .B(_08681_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20497_ (.A1(_08681_),
    .A2(_08682_),
    .B(_04761_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20498_ (.A1(\cs_registers_i.csr_mepc_o[9] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[9] ),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20499_ (.A1(\cs_registers_i.csr_depc_o[9] ),
    .A2(_08684_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20500_ (.A1(_07254_),
    .A2(_08363_),
    .B(_04763_),
    .C(_04764_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _20501_ (.I(net3254),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20502_ (.I0(net24),
    .I1(_04765_),
    .S(_04766_),
    .Z(_04767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20503_ (.A1(net3224),
    .A2(_04767_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20504_ (.A1(_04760_),
    .A2(_04768_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20505_ (.I(net3104),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20506_ (.A1(_07788_),
    .A2(_07789_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20507_ (.A1(_04770_),
    .A2(_04771_),
    .B(net319),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20508_ (.A1(net319),
    .A2(_04770_),
    .A3(_04771_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20509_ (.A1(\cs_registers_i.csr_mepc_o[8] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[8] ),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20510_ (.I(_04774_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20511_ (.A1(\cs_registers_i.csr_depc_o[8] ),
    .A2(_08684_),
    .B1(net3254),
    .B2(net23),
    .C(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _20512_ (.A1(_04772_),
    .A2(_04773_),
    .A3(_08363_),
    .B(_04776_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20513_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .I1(_04777_),
    .S(net3224),
    .Z(_04778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20514_ (.A1(\cs_registers_i.csr_depc_o[4] ),
    .A2(_08684_),
    .B1(_08709_),
    .B2(\cs_registers_i.csr_mepc_o[4] ),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _20515_ (.A1(_08669_),
    .A2(_02568_),
    .A3(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20516_ (.A1(_08624_),
    .A2(net175),
    .B(_04780_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20517_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .A2(net3224),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20518_ (.A1(_08378_),
    .A2(_04385_),
    .A3(_08665_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output163 (.I(net163),
    .Z(data_addr_o[22]));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20520_ (.A1(\cs_registers_i.csr_depc_o[5] ),
    .A2(_04783_),
    .B1(_04386_),
    .B2(\cs_registers_i.csr_mepc_o[5] ),
    .C(_02579_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20521_ (.A1(_08624_),
    .A2(net176),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _20522_ (.A1(_04785_),
    .A2(_04786_),
    .B(_08676_),
    .C(net3254),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20523_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .A2(net3222),
    .B(_04787_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20524_ (.A1(\cs_registers_i.csr_mepc_o[6] ),
    .A2(_04386_),
    .B(_02586_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20525_ (.A1(\cs_registers_i.csr_depc_o[6] ),
    .A2(_04783_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20526_ (.A1(_08669_),
    .A2(_04789_),
    .A3(_04790_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _20527_ (.A1(_07202_),
    .A2(_07203_),
    .A3(_08363_),
    .B(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20528_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .A2(net3224),
    .B(_04792_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _20529_ (.A1(_04781_),
    .A2(_04782_),
    .A3(_04788_),
    .A4(_04793_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20530_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20531_ (.A1(net178),
    .A2(_08624_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _20532_ (.A1(\cs_registers_i.csr_depc_o[7] ),
    .A2(_08684_),
    .B1(_08709_),
    .B2(\cs_registers_i.csr_mepc_o[7] ),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20533_ (.A1(net3223),
    .A2(_04766_),
    .A3(_04796_),
    .A4(_04797_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20534_ (.A1(_04795_),
    .A2(_08676_),
    .B(_04798_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20535_ (.A1(_11664_[0]),
    .A2(_04778_),
    .A3(_04794_),
    .A4(_04799_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20536_ (.A1(_04769_),
    .A2(_04800_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output162 (.I(net162),
    .Z(data_addr_o[21]));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20538_ (.A1(_11661_[0]),
    .A2(_04801_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .C(net3224),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output161 (.I(net161),
    .Z(data_addr_o[20]));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20540_ (.A1(net281),
    .A2(net286),
    .A3(_07306_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20541_ (.A1(net286),
    .A2(_07306_),
    .B(net281),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20542_ (.A1(\cs_registers_i.csr_mepc_o[10] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[10] ),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20543_ (.I(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20544_ (.A1(\cs_registers_i.csr_depc_o[10] ),
    .A2(_08684_),
    .B1(net3254),
    .B2(net1),
    .C(_04808_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _20545_ (.A1(_04805_),
    .A2(_04806_),
    .A3(_08363_),
    .B(_04809_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20546_ (.A1(net3221),
    .A2(_04810_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20547_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .A2(_11661_[0]),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20548_ (.I0(_04810_),
    .I1(_04812_),
    .S(net3221),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20549_ (.I0(_04811_),
    .I1(_04813_),
    .S(_04801_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20550_ (.A1(_04803_),
    .A2(_04814_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20551_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .A2(net3221),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20552_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(_04761_),
    .B(_08683_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20553_ (.A1(\cs_registers_i.csr_mepc_o[11] ),
    .A2(_08709_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20554_ (.A1(\cs_registers_i.csr_depc_o[11] ),
    .A2(_04783_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20555_ (.A1(_04816_),
    .A2(_04817_),
    .A3(_04818_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20556_ (.A1(_02927_),
    .A2(_08363_),
    .B(_04766_),
    .C(_04819_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _20557_ (.A1(net2),
    .A2(_04766_),
    .B(_04820_),
    .C(net3223),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20558_ (.A1(_04815_),
    .A2(_04821_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20559_ (.A1(_04794_),
    .A2(_04799_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20560_ (.A1(_11662_[0]),
    .A2(_11663_[0]),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20561_ (.A1(_04778_),
    .A2(_04823_),
    .A3(_04824_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20562_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .I1(_04810_),
    .S(net3224),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20563_ (.A1(_04769_),
    .A2(_04826_),
    .Z(_04827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20564_ (.A1(_04825_),
    .A2(_04827_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20565_ (.A1(_04822_),
    .A2(_04828_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20566_ (.A1(net3221),
    .A2(_08878_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output160 (.I(net160),
    .Z(data_addr_o[19]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20568_ (.I0(_04829_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .S(_04830_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _20569_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .A2(net3224),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20570_ (.A1(_04822_),
    .A2(_04827_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20571_ (.A1(_04800_),
    .A2(_04833_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20572_ (.A1(\cs_registers_i.csr_mepc_o[12] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[12] ),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20573_ (.A1(\cs_registers_i.csr_depc_o[12] ),
    .A2(_04783_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20574_ (.A1(net3),
    .A2(net3254),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _20575_ (.A1(net3223),
    .A2(_04835_),
    .A3(_04836_),
    .A4(_04837_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20576_ (.A1(net153),
    .A2(_08624_),
    .B(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20577_ (.I(_04839_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20578_ (.A1(_04834_),
    .A2(_04840_),
    .B(_04830_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20579_ (.A1(_11661_[0]),
    .A2(_04832_),
    .B(_04839_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20580_ (.A1(_04832_),
    .A2(_04841_),
    .B1(_04842_),
    .B2(_04834_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20581_ (.A1(\cs_registers_i.csr_mepc_o[13] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[13] ),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20582_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(_04783_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20583_ (.A1(_04843_),
    .A2(_04844_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20584_ (.A1(net154),
    .A2(_08624_),
    .B1(net3254),
    .B2(net4),
    .C(_04845_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20585_ (.A1(net3224),
    .A2(_04846_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20586_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .A2(net3224),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20587_ (.A1(_04847_),
    .A2(_04848_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20588_ (.A1(_04832_),
    .A2(_04839_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20589_ (.A1(_04825_),
    .A2(_04833_),
    .A3(_04850_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20590_ (.A1(_04849_),
    .A2(_04851_),
    .Z(_04852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20591_ (.I0(_04852_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .S(_04830_),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20592_ (.A1(_04760_),
    .A2(_04768_),
    .B(_04832_),
    .C(_04839_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20593_ (.A1(_04822_),
    .A2(_04826_),
    .A3(_04849_),
    .A4(_04853_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20594_ (.A1(_04800_),
    .A2(_04854_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20595_ (.A1(_08878_),
    .A2(_04855_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20596_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .A2(_04856_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output159 (.I(net159),
    .Z(data_addr_o[18]));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20598_ (.A1(\cs_registers_i.csr_mepc_o[14] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[14] ),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20599_ (.A1(\cs_registers_i.csr_depc_o[14] ),
    .A2(_04783_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20600_ (.A1(_04859_),
    .A2(_04860_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20601_ (.A1(_08624_),
    .A2(net3097),
    .B1(net3254),
    .B2(net5),
    .C(_04861_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20602_ (.A1(_04855_),
    .A2(net363),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20603_ (.I0(_04857_),
    .I1(_04863_),
    .S(net3224),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20604_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20605_ (.A1(net156),
    .A2(_08624_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20606_ (.A1(\cs_registers_i.csr_mepc_o[15] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[15] ),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output158 (.I(net158),
    .Z(data_addr_o[17]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20608_ (.A1(\cs_registers_i.csr_depc_o[15] ),
    .A2(_04783_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20609_ (.A1(net6),
    .A2(net3254),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20610_ (.A1(net3223),
    .A2(_04866_),
    .A3(_04868_),
    .A4(_04869_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20611_ (.A1(_04864_),
    .A2(net3221),
    .B1(_04865_),
    .B2(_04870_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20612_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .A2(net3224),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20613_ (.A1(net3224),
    .A2(_04862_),
    .B(_04872_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20614_ (.A1(_04825_),
    .A2(_04854_),
    .A3(_04873_),
    .Z(_04874_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20615_ (.A1(_04871_),
    .A2(_04874_),
    .Z(_04875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20616_ (.I0(_04875_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .S(_04830_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20617_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20618_ (.A1(net7),
    .A2(net3254),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20619_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(_04761_),
    .B(_08683_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20620_ (.A1(\cs_registers_i.csr_depc_o[16] ),
    .A2(_04783_),
    .B1(_04386_),
    .B2(\cs_registers_i.csr_mepc_o[16] ),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20621_ (.A1(net3224),
    .A2(_04877_),
    .A3(_04878_),
    .A4(_04879_),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20622_ (.A1(net157),
    .A2(_08624_),
    .B(_04880_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20623_ (.A1(_04876_),
    .A2(net3221),
    .B(_04881_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20624_ (.A1(_04800_),
    .A2(_04854_),
    .A3(_04871_),
    .A4(_04873_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20625_ (.A1(net405),
    .A2(_04883_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20626_ (.I0(_04884_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .S(_04830_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20627_ (.A1(\cs_registers_i.csr_mepc_o[17] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[17] ),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20628_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(_04783_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20629_ (.A1(_04885_),
    .A2(_04886_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20630_ (.A1(net158),
    .A2(_08624_),
    .B1(net3254),
    .B2(net8),
    .C(_04887_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20631_ (.A1(net3221),
    .A2(_04888_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20632_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .A2(net3221),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20633_ (.A1(_04889_),
    .A2(_04890_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20634_ (.A1(_04854_),
    .A2(_04871_),
    .A3(_04873_),
    .A4(net406),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20635_ (.A1(_04825_),
    .A2(_04892_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20636_ (.A1(_04891_),
    .A2(_04893_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20637_ (.I0(_04894_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .S(_04830_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20638_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20639_ (.A1(net159),
    .A2(_08624_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20640_ (.A1(\cs_registers_i.csr_mepc_o[18] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[18] ),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20641_ (.A1(\cs_registers_i.csr_depc_o[18] ),
    .A2(_04783_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20642_ (.A1(net9),
    .A2(net3254),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20643_ (.A1(net3224),
    .A2(_04897_),
    .A3(_04898_),
    .A4(_04899_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _20644_ (.A1(_04895_),
    .A2(net3221),
    .B1(_04896_),
    .B2(_04900_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20645_ (.A1(_04800_),
    .A2(_04891_),
    .A3(_04892_),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20646_ (.A1(_04901_),
    .A2(_04902_),
    .Z(_04903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20647_ (.I0(_04903_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .S(_04830_),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20648_ (.A1(\cs_registers_i.csr_mepc_o[19] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[19] ),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20649_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(_04783_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20650_ (.A1(_04904_),
    .A2(_04905_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20651_ (.A1(net160),
    .A2(_08624_),
    .B1(net3254),
    .B2(net10),
    .C(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20652_ (.A1(net3221),
    .A2(_04907_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20653_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .A2(net3221),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20654_ (.A1(_04908_),
    .A2(_04909_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20655_ (.A1(_04891_),
    .A2(_04901_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20656_ (.A1(_04825_),
    .A2(_04892_),
    .A3(_04911_),
    .Z(_04912_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20657_ (.A1(_04910_),
    .A2(_04912_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20658_ (.I0(_04913_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .S(_04830_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20659_ (.A1(_07788_),
    .A2(_07789_),
    .A3(_07794_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20660_ (.I(net386),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20661_ (.A1(net343),
    .A2(_04914_),
    .A3(_04915_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20662_ (.A1(_04914_),
    .A2(_04915_),
    .B(net343),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20663_ (.A1(net11),
    .A2(net3254),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20664_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_04761_),
    .B(_08683_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20665_ (.A1(\cs_registers_i.csr_depc_o[20] ),
    .A2(_04783_),
    .B1(_04386_),
    .B2(\cs_registers_i.csr_mepc_o[20] ),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20666_ (.A1(net3223),
    .A2(_04918_),
    .A3(_04919_),
    .A4(_04920_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20667_ (.A1(_04916_),
    .A2(_04917_),
    .A3(_08363_),
    .B(_04921_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20668_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .A2(net3224),
    .Z(_04923_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20669_ (.A1(_04922_),
    .A2(_04923_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20670_ (.A1(_04901_),
    .A2(_04910_),
    .Z(_04925_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20671_ (.A1(_04800_),
    .A2(_04891_),
    .A3(_04892_),
    .A4(_04925_),
    .Z(_04926_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20672_ (.A1(_04924_),
    .A2(_04926_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20673_ (.I0(_04927_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .S(_04830_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20674_ (.A1(\cs_registers_i.csr_mepc_o[21] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[21] ),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20675_ (.I(_04928_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20676_ (.A1(\cs_registers_i.csr_depc_o[21] ),
    .A2(_08684_),
    .B1(net3254),
    .B2(net12),
    .C(_04929_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20677_ (.A1(_08363_),
    .A2(_07787_),
    .B(_04930_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20678_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .I1(_04931_),
    .S(net3224),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20679_ (.A1(_04825_),
    .A2(_04891_),
    .A3(_04892_),
    .A4(_04925_),
    .Z(_04933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20680_ (.A1(_04933_),
    .A2(_04924_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20681_ (.A1(net391),
    .A2(_04934_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20682_ (.I0(_04935_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .S(_04830_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20683_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _20684_ (.A1(_07894_),
    .A2(_07897_),
    .A3(_07902_),
    .A4(_08363_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20685_ (.A1(\cs_registers_i.csr_mepc_o[22] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[22] ),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20686_ (.A1(\cs_registers_i.csr_depc_o[22] ),
    .A2(_04783_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20687_ (.A1(net13),
    .A2(net3254),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20688_ (.A1(net3224),
    .A2(_04938_),
    .A3(_04939_),
    .A4(_04940_),
    .Z(_04941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _20689_ (.A1(_04936_),
    .A2(net3222),
    .B1(_04937_),
    .B2(_04941_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20690_ (.A1(_04924_),
    .A2(_04932_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20691_ (.A1(_04926_),
    .A2(_04943_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20692_ (.A1(net633),
    .A2(_04944_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output157 (.I(net157),
    .Z(data_addr_o[16]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20694_ (.I0(_04945_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .S(_04830_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20695_ (.A1(\cs_registers_i.csr_mepc_o[23] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[23] ),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20696_ (.A1(\cs_registers_i.csr_depc_o[23] ),
    .A2(_04783_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20697_ (.A1(_04947_),
    .A2(_04948_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20698_ (.A1(_08624_),
    .A2(net164),
    .B1(net3254),
    .B2(net14),
    .C(_04949_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20699_ (.A1(_04950_),
    .A2(net3221),
    .Z(_04951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20700_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .A2(_08676_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20701_ (.A1(_04952_),
    .A2(_04951_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20702_ (.A1(_04933_),
    .A2(_04942_),
    .A3(_04943_),
    .Z(_04954_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20703_ (.A1(net375),
    .A2(_04954_),
    .Z(_04955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20704_ (.I0(_04955_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .S(_04830_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20705_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20706_ (.A1(_04956_),
    .A2(net3221),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20707_ (.A1(\cs_registers_i.csr_mepc_o[24] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[24] ),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20708_ (.A1(\cs_registers_i.csr_depc_o[24] ),
    .A2(_04783_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20709_ (.A1(net15),
    .A2(net3254),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20710_ (.A1(net3224),
    .A2(_04958_),
    .A3(_04959_),
    .A4(_04960_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20711_ (.A1(_08624_),
    .A2(net165),
    .B(_04961_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20712_ (.A1(_04924_),
    .A2(net391),
    .A3(_04942_),
    .A4(_04953_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20713_ (.A1(_04926_),
    .A2(_04963_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20714_ (.A1(net380),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20715_ (.A1(_04956_),
    .A2(_11661_[0]),
    .A3(_04926_),
    .A4(_04963_),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20716_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .A2(_08878_),
    .B(_04966_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output156 (.I(net156),
    .Z(data_addr_o[15]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output155 (.I(net3097),
    .Z(data_addr_o[14]));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20719_ (.A1(_04957_),
    .A2(_04965_),
    .B1(_04967_),
    .B2(net3224),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20720_ (.A1(net16),
    .A2(net3254),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20721_ (.A1(\cs_registers_i.csr_mtvec_o[25] ),
    .A2(_04761_),
    .B(_08683_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20722_ (.A1(\cs_registers_i.csr_depc_o[25] ),
    .A2(_04783_),
    .B1(_04386_),
    .B2(\cs_registers_i.csr_mepc_o[25] ),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20723_ (.A1(_08624_),
    .A2(net166),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _20724_ (.A1(_04971_),
    .A2(_04973_),
    .A3(_04972_),
    .A4(_04970_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20725_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .I1(_04974_),
    .S(net3224),
    .Z(_04975_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _20726_ (.A1(_04957_),
    .A2(_04962_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20727_ (.A1(_04933_),
    .A2(_04963_),
    .A3(_04976_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20728_ (.A1(_04975_),
    .A2(_04977_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20729_ (.I0(_04978_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .S(_04830_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20730_ (.A1(_04800_),
    .A2(_04910_),
    .Z(_04979_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20731_ (.A1(_04963_),
    .A2(_04975_),
    .A3(_04976_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20732_ (.A1(_04892_),
    .A2(_04911_),
    .A3(_04979_),
    .A4(_04980_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20733_ (.A1(_11661_[0]),
    .A2(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20734_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .A2(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20735_ (.A1(\cs_registers_i.csr_mepc_o[26] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[26] ),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20736_ (.I(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20737_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(_08684_),
    .B1(net3254),
    .B2(net17),
    .C(_04985_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20738_ (.A1(_08363_),
    .A2(_08078_),
    .B(_04986_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20739_ (.A1(_04981_),
    .A2(net358),
    .Z(_04988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20740_ (.I0(_04983_),
    .I1(_04988_),
    .S(net3224),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20741_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_04761_),
    .B(_08683_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20742_ (.A1(\cs_registers_i.csr_depc_o[27] ),
    .A2(_04783_),
    .B1(_04386_),
    .B2(\cs_registers_i.csr_mepc_o[27] ),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20743_ (.A1(_04989_),
    .A2(_04990_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20744_ (.A1(net168),
    .A2(_08624_),
    .B1(net3254),
    .B2(net18),
    .C(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20745_ (.A1(net3221),
    .A2(_04992_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20746_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .A2(net3221),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20747_ (.A1(_04993_),
    .A2(_04994_),
    .Z(_04995_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20748_ (.A1(_04825_),
    .A2(_04892_),
    .A3(_04910_),
    .A4(_04911_),
    .Z(_04996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20749_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .I1(_04987_),
    .S(net3224),
    .Z(_04997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20750_ (.A1(_04980_),
    .A2(net346),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20751_ (.A1(_04996_),
    .A2(_04998_),
    .Z(_04999_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20752_ (.A1(_04995_),
    .A2(_04999_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20753_ (.I0(_05000_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .S(_04830_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20754_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _20755_ (.A1(_08154_),
    .A2(_08160_),
    .B(_08363_),
    .C(_08161_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20756_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(_04761_),
    .B(_08683_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20757_ (.A1(\cs_registers_i.csr_depc_o[28] ),
    .A2(_04783_),
    .B1(_04386_),
    .B2(\cs_registers_i.csr_mepc_o[28] ),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20758_ (.A1(_05003_),
    .A2(_05004_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20759_ (.A1(net19),
    .A2(_04766_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _20760_ (.A1(net3254),
    .A2(_05002_),
    .A3(_05005_),
    .B(_05006_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20761_ (.I0(_05001_),
    .I1(_05007_),
    .S(net3224),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20762_ (.A1(_04994_),
    .A2(_04993_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20763_ (.A1(_04981_),
    .A2(net346),
    .A3(_05009_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20764_ (.A1(_05008_),
    .A2(_05010_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20765_ (.I0(_05011_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .S(_04830_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20766_ (.A1(\cs_registers_i.csr_mepc_o[29] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[29] ),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20767_ (.A1(\cs_registers_i.csr_depc_o[29] ),
    .A2(_04783_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20768_ (.A1(_05012_),
    .A2(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20769_ (.A1(net170),
    .A2(_08624_),
    .B1(net3254),
    .B2(net20),
    .C(_05014_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20770_ (.A1(net3221),
    .A2(_05015_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20771_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .A2(net3221),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20772_ (.A1(_05016_),
    .A2(_05017_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20773_ (.A1(_04995_),
    .A2(net625),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20774_ (.A1(_04996_),
    .A2(_04998_),
    .A3(_05019_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20775_ (.A1(net461),
    .A2(_05020_),
    .Z(_05021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20776_ (.I0(_05021_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .S(_04830_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20777_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .S(_04830_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20778_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20779_ (.A1(\cs_registers_i.csr_mepc_o[30] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[30] ),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20780_ (.A1(\cs_registers_i.csr_depc_o[30] ),
    .A2(_04783_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20781_ (.A1(net21),
    .A2(net3254),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _20782_ (.A1(net3223),
    .A2(_05023_),
    .A3(_05024_),
    .A4(_05025_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20783_ (.A1(_08624_),
    .A2(net172),
    .B(_05026_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20784_ (.A1(_05022_),
    .A2(_08676_),
    .B(_05027_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20785_ (.A1(_05018_),
    .A2(_05019_),
    .Z(_05029_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20786_ (.A1(_04981_),
    .A2(_04997_),
    .A3(_05029_),
    .Z(_05030_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20787_ (.A1(net397),
    .A2(_05030_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20788_ (.I0(_05031_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .S(_04830_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20789_ (.A1(\cs_registers_i.csr_mepc_o[31] ),
    .A2(_04386_),
    .B1(_04762_),
    .B2(\cs_registers_i.csr_mtvec_o[31] ),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20790_ (.A1(\cs_registers_i.csr_depc_o[31] ),
    .A2(_04783_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20791_ (.A1(_05032_),
    .A2(_05033_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20792_ (.A1(net173),
    .A2(_08624_),
    .B1(net3254),
    .B2(net22),
    .C(_05034_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20793_ (.A1(net3222),
    .A2(_05035_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20794_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .A2(net3221),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20795_ (.A1(_05036_),
    .A2(_05037_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20796_ (.A1(_04996_),
    .A2(_04998_),
    .A3(net397),
    .A4(_05029_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20797_ (.A1(net336),
    .A2(_05039_),
    .Z(_05040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20798_ (.I0(_05040_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .S(_04830_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20799_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .S(_04830_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20800_ (.A1(_04781_),
    .A2(_04782_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20801_ (.A1(_11664_[0]),
    .A2(_05041_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20802_ (.I0(_05042_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .S(_04830_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20803_ (.A1(_05041_),
    .A2(_04824_),
    .Z(_05043_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20804_ (.A1(_04788_),
    .A2(_05043_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20805_ (.I0(_05044_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .S(_04830_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20806_ (.I(_04788_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20807_ (.A1(_11664_[0]),
    .A2(_05041_),
    .A3(_05045_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20808_ (.A1(_04793_),
    .A2(_05046_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20809_ (.I0(_05047_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .S(_04830_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20810_ (.A1(_04794_),
    .A2(_04824_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20811_ (.A1(_04799_),
    .A2(_05048_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20812_ (.I0(_05049_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .S(_04830_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20813_ (.A1(_11664_[0]),
    .A2(_04823_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20814_ (.A1(_08878_),
    .A2(_05050_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20815_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .A2(_05051_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20816_ (.A1(_04777_),
    .A2(_05050_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20817_ (.I0(_05052_),
    .I1(_05053_),
    .S(net3224),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20818_ (.A1(_04769_),
    .A2(_04825_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20819_ (.I0(_05054_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .S(_04830_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output154 (.I(net154),
    .Z(data_addr_o[13]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20821_ (.I0(net94),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20822_ (.I(_05056_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20823_ (.A1(_04361_),
    .A2(_04327_),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .C(_08658_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20824_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_08658_),
    .B(_05058_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20825_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net128),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20826_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_05060_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20827_ (.A1(_08736_),
    .A2(_05061_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output153 (.I(net153),
    .Z(data_addr_o[12]));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _20829_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_05060_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20830_ (.A1(net3652),
    .A2(_05064_),
    .Z(_05065_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20831_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(_05065_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20832_ (.A1(net3653),
    .A2(_08745_),
    .Z(_05067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20833_ (.I0(_05062_),
    .I1(_05066_),
    .S(_05067_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _20834_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_05059_),
    .B(_05068_),
    .C(_04343_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 _20835_ (.I(net3651),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _20836_ (.I(_08739_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20837_ (.A1(_06782_),
    .A2(_01973_),
    .Z(_05072_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20838_ (.A1(_05070_),
    .A2(_05071_),
    .A3(_05072_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _20839_ (.A1(_04364_),
    .A2(_05069_),
    .A3(_05073_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20840_ (.A1(_01987_),
    .A2(_05074_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output152 (.I(net152),
    .Z(data_addr_o[11]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output151 (.I(net151),
    .Z(data_addr_o[10]));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _20843_ (.A1(_05071_),
    .A2(_05072_),
    .A3(_04364_),
    .A4(_05069_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20844_ (.A1(_08736_),
    .A2(_05064_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20845_ (.A1(_01987_),
    .A2(_05078_),
    .B(_05079_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output150 (.I(net150),
    .Z(core_sleep_o));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20847_ (.A1(_05075_),
    .A2(net3072),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20848_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20849_ (.A1(_05057_),
    .A2(_05064_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20850_ (.A1(_01987_),
    .A2(_05078_),
    .Z(_05085_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input149 (.I(test_en_i),
    .Z(net149));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20852_ (.I0(_05083_),
    .I1(_05084_),
    .S(net3071),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input148 (.I(rst_ni),
    .Z(net148));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input147 (.I(irq_timer_i),
    .Z(net147));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input146 (.I(irq_software_i),
    .Z(net146));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input145 (.I(irq_nm_i),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20857_ (.A1(_08736_),
    .A2(_05070_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input144 (.I(irq_fast_i[9]),
    .Z(net144));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20859_ (.A1(_05083_),
    .A2(_05092_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20860_ (.A1(_01987_),
    .A2(_05078_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _20861_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .A2(_05064_),
    .A3(_05075_),
    .B1(_05094_),
    .B2(_05095_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20862_ (.A1(_05057_),
    .A2(_05082_),
    .B1(_05087_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .C(_05096_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input143 (.I(irq_fast_i[8]),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20864_ (.I0(net94),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20865_ (.A1(_01987_),
    .A2(_05078_),
    .B(net3651),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20866_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(_01987_),
    .A3(_05078_),
    .Z(_05100_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20867_ (.A1(_05064_),
    .A2(_05075_),
    .B1(_05099_),
    .B2(_05065_),
    .C(_05100_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input142 (.I(irq_fast_i[7]),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20869_ (.I0(_05098_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .S(net3058),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input141 (.I(irq_fast_i[6]),
    .Z(net141));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input140 (.I(irq_fast_i[5]),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _20872_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A3(_05061_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input139 (.I(irq_fast_i[4]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20874_ (.I0(net94),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .S(_05105_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20875_ (.A1(\alu_adder_result_ex[1] ),
    .A2(_08624_),
    .Z(_05107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20876_ (.A1(\cs_registers_i.csr_depc_o[1] ),
    .A2(_08684_),
    .B1(_08709_),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .C(_05107_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _20877_ (.A1(_05072_),
    .A2(_04364_),
    .A3(_05069_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input138 (.I(irq_fast_i[3]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input137 (.I(irq_fast_i[2]),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20880_ (.A1(_01987_),
    .A2(_05109_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input136 (.I(irq_fast_i[1]),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20882_ (.A1(_08745_),
    .A2(_05112_),
    .B(net3653),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20883_ (.A1(_01987_),
    .A2(_05109_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input135 (.I(irq_fast_i[14]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input134 (.I(irq_fast_i[13]),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20886_ (.A1(_05071_),
    .A2(net3070),
    .B(_08669_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20887_ (.A1(_08669_),
    .A2(_05108_),
    .B1(_05114_),
    .B2(_05118_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input133 (.I(irq_fast_i[12]),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20889_ (.A1(\cs_registers_i.pc_if_i[9] ),
    .A2(\cs_registers_i.pc_if_i[10] ),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _20890_ (.I(\cs_registers_i.pc_if_i[3] ),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _20891_ (.A1(_05121_),
    .A2(_11000_[0]),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20892_ (.A1(\cs_registers_i.pc_if_i[4] ),
    .A2(\cs_registers_i.pc_if_i[5] ),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20893_ (.A1(\cs_registers_i.pc_if_i[6] ),
    .A2(\cs_registers_i.pc_if_i[7] ),
    .A3(_05123_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20894_ (.A1(\cs_registers_i.pc_if_i[8] ),
    .A2(_05124_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20895_ (.A1(_05122_),
    .A2(_05125_),
    .Z(_05126_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20896_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05120_),
    .A4(_05126_),
    .Z(_05127_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20897_ (.A1(\cs_registers_i.pc_if_i[11] ),
    .A2(_05127_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20898_ (.A1(net3224),
    .A2(_05128_),
    .B(_04821_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input132 (.I(irq_fast_i[11]),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20900_ (.A1(net3653),
    .A2(_11390_[0]),
    .A3(_08746_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20901_ (.A1(_11389_[0]),
    .A2(_05130_),
    .Z(_05131_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20902_ (.A1(\cs_registers_i.pc_if_i[3] ),
    .A2(_05131_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input131 (.I(irq_fast_i[10]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20904_ (.A1(\cs_registers_i.pc_if_i[11] ),
    .A2(_05125_),
    .A3(_05120_),
    .A4(_05132_),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20905_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05134_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20906_ (.A1(\cs_registers_i.pc_if_i[12] ),
    .A2(_05135_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20907_ (.A1(net3221),
    .A2(_05136_),
    .B(_04839_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20908_ (.A1(\cs_registers_i.pc_if_i[11] ),
    .A2(\cs_registers_i.pc_if_i[12] ),
    .A3(_05120_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20909_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05126_),
    .A4(_05137_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20910_ (.A1(\cs_registers_i.pc_if_i[13] ),
    .A2(_05138_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20911_ (.I(_04847_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20912_ (.A1(net3221),
    .A2(_05139_),
    .B(_05140_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20913_ (.A1(\cs_registers_i.pc_if_i[13] ),
    .A2(_05137_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20914_ (.A1(_05125_),
    .A2(_05132_),
    .A3(_05141_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20915_ (.A1(net3070),
    .A2(_05142_),
    .B(\cs_registers_i.pc_if_i[14] ),
    .C(net3224),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20916_ (.A1(\cs_registers_i.pc_if_i[14] ),
    .A2(net3221),
    .A3(net3070),
    .A4(_05142_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20917_ (.A1(net3224),
    .A2(net362),
    .B(_05143_),
    .C(_05144_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20918_ (.A1(\cs_registers_i.pc_if_i[14] ),
    .A2(_05141_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20919_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05126_),
    .A4(_05145_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20920_ (.A1(\cs_registers_i.pc_if_i[15] ),
    .A2(_05146_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20921_ (.A1(_04865_),
    .A2(_04870_),
    .B1(_05147_),
    .B2(net3221),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20922_ (.A1(\cs_registers_i.pc_if_i[15] ),
    .A2(_05145_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20923_ (.A1(_05125_),
    .A2(_05132_),
    .A3(_05148_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20924_ (.A1(net3070),
    .A2(_05149_),
    .B(\cs_registers_i.pc_if_i[16] ),
    .C(net3224),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20925_ (.A1(\cs_registers_i.pc_if_i[16] ),
    .A2(net3221),
    .A3(net3070),
    .A4(_05149_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _20926_ (.A1(_04881_),
    .A2(_05150_),
    .A3(_05151_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20927_ (.I(\cs_registers_i.pc_if_i[17] ),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _20928_ (.A1(net3084),
    .A2(_05109_),
    .B(net3223),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20929_ (.A1(_05122_),
    .A2(_05125_),
    .A3(_05148_),
    .Z(_05154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20930_ (.A1(\cs_registers_i.pc_if_i[16] ),
    .A2(_05154_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20931_ (.A1(_04889_),
    .A2(_05155_),
    .Z(_05156_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20932_ (.A1(_05153_),
    .A2(_05156_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20933_ (.A1(\cs_registers_i.pc_if_i[16] ),
    .A2(\cs_registers_i.pc_if_i[17] ),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20934_ (.A1(_05154_),
    .A2(_05158_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input130 (.I(irq_fast_i[0]),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20936_ (.A1(_05112_),
    .A2(_05159_),
    .B(net3221),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20937_ (.A1(_05152_),
    .A2(_05157_),
    .B1(_05161_),
    .B2(_04889_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20938_ (.A1(_05125_),
    .A2(_05132_),
    .A3(_05148_),
    .A4(_05158_),
    .Z(_05162_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20939_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05162_),
    .Z(_05163_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20940_ (.A1(\cs_registers_i.pc_if_i[18] ),
    .A2(_05163_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20941_ (.A1(_04896_),
    .A2(_04900_),
    .B1(_05164_),
    .B2(net3221),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20942_ (.I(\cs_registers_i.pc_if_i[19] ),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20943_ (.A1(\cs_registers_i.pc_if_i[18] ),
    .A2(_05154_),
    .A3(_05158_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20944_ (.A1(_04908_),
    .A2(_05166_),
    .Z(_05167_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20945_ (.A1(_05153_),
    .A2(_05167_),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _20946_ (.A1(\cs_registers_i.pc_if_i[18] ),
    .A2(\cs_registers_i.pc_if_i[19] ),
    .A3(_05158_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20947_ (.A1(_05154_),
    .A2(_05169_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20948_ (.I(_05170_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20949_ (.A1(_05112_),
    .A2(_05171_),
    .B(net3221),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20950_ (.A1(_05165_),
    .A2(_05168_),
    .B1(_05172_),
    .B2(_04908_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20951_ (.A1(net161),
    .A2(_08624_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20952_ (.A1(_05125_),
    .A2(_05132_),
    .A3(_05148_),
    .A4(_05169_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20953_ (.A1(net3070),
    .A2(_05174_),
    .B(\cs_registers_i.pc_if_i[20] ),
    .C(net3223),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20954_ (.A1(\cs_registers_i.pc_if_i[20] ),
    .A2(net3222),
    .A3(net3070),
    .A4(_05174_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20955_ (.A1(_05173_),
    .A2(_04921_),
    .B(_05175_),
    .C(_05176_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20956_ (.I0(_10997_[0]),
    .I1(_11001_[0]),
    .S(net3070),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20957_ (.A1(_08669_),
    .A2(_05177_),
    .B(_08713_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20958_ (.I(\cs_registers_i.pc_if_i[21] ),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20959_ (.A1(net3223),
    .A2(net392),
    .B1(_05170_),
    .B2(\cs_registers_i.pc_if_i[20] ),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20960_ (.A1(_05153_),
    .A2(_05179_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20961_ (.A1(\cs_registers_i.pc_if_i[20] ),
    .A2(\cs_registers_i.pc_if_i[21] ),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20962_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05170_),
    .A4(_05181_),
    .Z(_05182_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20963_ (.A1(net3223),
    .A2(_05182_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20964_ (.A1(net3223),
    .A2(net392),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20965_ (.A1(_05178_),
    .A2(_05180_),
    .B1(_05183_),
    .B2(_05184_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20966_ (.A1(_05125_),
    .A2(_05132_),
    .A3(_05148_),
    .A4(_05169_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20967_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05185_),
    .A4(_05181_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20968_ (.A1(\cs_registers_i.pc_if_i[22] ),
    .A2(_05186_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20969_ (.A1(_04937_),
    .A2(_04941_),
    .B1(_05187_),
    .B2(net3222),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20970_ (.I(\cs_registers_i.pc_if_i[23] ),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20971_ (.A1(\cs_registers_i.pc_if_i[22] ),
    .A2(_05181_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20972_ (.A1(_05170_),
    .A2(_05189_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20973_ (.A1(_05188_),
    .A2(_05112_),
    .A3(_05190_),
    .B(net3221),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20974_ (.A1(_04951_),
    .A2(_05190_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20975_ (.A1(_05153_),
    .A2(_05192_),
    .Z(_05193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20976_ (.A1(_04951_),
    .A2(_05191_),
    .B1(_05193_),
    .B2(_05188_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20977_ (.A1(_05185_),
    .A2(_05189_),
    .Z(_05194_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20978_ (.A1(\cs_registers_i.pc_if_i[23] ),
    .A2(net3084),
    .A3(_05109_),
    .A4(_05194_),
    .Z(_05195_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20979_ (.A1(\cs_registers_i.pc_if_i[24] ),
    .A2(_05195_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20980_ (.A1(_08676_),
    .A2(_05196_),
    .B(net381),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20981_ (.I(\cs_registers_i.pc_if_i[25] ),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20982_ (.A1(\cs_registers_i.pc_if_i[23] ),
    .A2(\cs_registers_i.pc_if_i[24] ),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20983_ (.A1(net3224),
    .A2(_04974_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20984_ (.A1(_05190_),
    .A2(_05198_),
    .B(_05199_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20985_ (.A1(net3224),
    .A2(net3070),
    .B(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _20986_ (.A1(_05126_),
    .A2(_05148_),
    .A3(_05169_),
    .A4(_05189_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20987_ (.A1(_05197_),
    .A2(_05198_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20988_ (.A1(_05202_),
    .A2(_05203_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20989_ (.A1(_05112_),
    .A2(_05204_),
    .B(net3221),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20990_ (.A1(_05197_),
    .A2(_05201_),
    .B1(_05205_),
    .B2(_05199_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20991_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05194_),
    .A4(_05203_),
    .Z(_05206_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20992_ (.A1(\cs_registers_i.pc_if_i[26] ),
    .A2(_05206_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20993_ (.I0(_04987_),
    .I1(_05207_),
    .S(net3222),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20994_ (.I(\cs_registers_i.pc_if_i[27] ),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20995_ (.A1(\cs_registers_i.pc_if_i[26] ),
    .A2(_05203_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20996_ (.A1(_05202_),
    .A2(_05209_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20997_ (.A1(_04993_),
    .A2(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20998_ (.A1(net3224),
    .A2(net3070),
    .B(_05211_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20999_ (.A1(\cs_registers_i.pc_if_i[27] ),
    .A2(_05209_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21000_ (.A1(_05202_),
    .A2(_05213_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21001_ (.A1(_05112_),
    .A2(_05214_),
    .B(_08676_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21002_ (.A1(_05208_),
    .A2(_05212_),
    .B1(_05215_),
    .B2(_04993_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21003_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05194_),
    .A4(_05213_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21004_ (.A1(\cs_registers_i.pc_if_i[28] ),
    .A2(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21005_ (.A1(net3224),
    .A2(_05007_),
    .Z(_05218_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21006_ (.A1(_08676_),
    .A2(_05217_),
    .B(_05218_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21007_ (.I(\cs_registers_i.pc_if_i[29] ),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21008_ (.A1(\cs_registers_i.pc_if_i[28] ),
    .A2(_05213_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21009_ (.A1(_05190_),
    .A2(_05220_),
    .B(net340),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21010_ (.A1(net3224),
    .A2(net3070),
    .B(_05221_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21011_ (.A1(_05219_),
    .A2(_05220_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21012_ (.A1(_05202_),
    .A2(_05223_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21013_ (.A1(_05112_),
    .A2(_05224_),
    .B(_08676_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21014_ (.A1(_05219_),
    .A2(_05222_),
    .B1(_05225_),
    .B2(net340),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21015_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05194_),
    .A4(_05223_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21016_ (.A1(\cs_registers_i.pc_if_i[30] ),
    .A2(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21017_ (.A1(net3222),
    .A2(_05227_),
    .B(_05027_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21018_ (.A1(_11000_[0]),
    .A2(_08728_),
    .Z(_05228_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21019_ (.A1(_05153_),
    .A2(_05228_),
    .Z(_05229_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21020_ (.A1(_05121_),
    .A2(_11000_[0]),
    .A3(_05112_),
    .B(net3222),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21021_ (.A1(_05121_),
    .A2(_05229_),
    .B1(_05230_),
    .B2(_08728_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21022_ (.I(\cs_registers_i.pc_if_i[31] ),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21023_ (.A1(\cs_registers_i.pc_if_i[30] ),
    .A2(_05202_),
    .A3(_05223_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21024_ (.A1(_05231_),
    .A2(_05112_),
    .A3(_05232_),
    .B(net3222),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21025_ (.A1(_05036_),
    .A2(_05232_),
    .Z(_05234_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21026_ (.A1(_05153_),
    .A2(_05234_),
    .Z(_05235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21027_ (.A1(_05036_),
    .A2(_05233_),
    .B1(_05235_),
    .B2(_05231_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21028_ (.A1(net3070),
    .A2(_05132_),
    .B(\cs_registers_i.pc_if_i[4] ),
    .C(net3223),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21029_ (.A1(\cs_registers_i.pc_if_i[4] ),
    .A2(net3222),
    .A3(net3070),
    .A4(_05132_),
    .Z(_05237_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21030_ (.A1(_04781_),
    .A2(_05236_),
    .A3(_05237_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21031_ (.I(\cs_registers_i.pc_if_i[5] ),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21032_ (.A1(\cs_registers_i.pc_if_i[4] ),
    .A2(_05122_),
    .B(_04787_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21033_ (.A1(_05153_),
    .A2(_05239_),
    .Z(_05240_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _21034_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05122_),
    .A4(_05123_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21035_ (.A1(net3222),
    .A2(_05241_),
    .B(_04787_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21036_ (.A1(_05238_),
    .A2(_05240_),
    .B(_05242_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21037_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05123_),
    .A4(_05132_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21038_ (.A1(\cs_registers_i.pc_if_i[6] ),
    .A2(_05243_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21039_ (.I(_04792_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21040_ (.A1(net3222),
    .A2(_05244_),
    .B(_05245_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21041_ (.A1(\cs_registers_i.pc_if_i[6] ),
    .A2(_05122_),
    .A3(_05123_),
    .Z(_05246_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21042_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05246_),
    .Z(_05247_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21043_ (.A1(\cs_registers_i.pc_if_i[7] ),
    .A2(_05247_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21044_ (.A1(net3222),
    .A2(_05248_),
    .B(_04798_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21045_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05124_),
    .A4(_05132_),
    .Z(_05249_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21046_ (.A1(\cs_registers_i.pc_if_i[8] ),
    .A2(_05249_),
    .Z(_05250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21047_ (.I0(_04777_),
    .I1(_05250_),
    .S(net3222),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21048_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05126_),
    .Z(_05251_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21049_ (.A1(\cs_registers_i.pc_if_i[9] ),
    .A2(_05251_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21050_ (.A1(net3224),
    .A2(_05252_),
    .B(_04768_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21051_ (.A1(\cs_registers_i.pc_if_i[9] ),
    .A2(_05125_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21052_ (.A1(net3084),
    .A2(_05109_),
    .A3(_05132_),
    .A4(_05253_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21053_ (.A1(\cs_registers_i.pc_if_i[10] ),
    .A2(_05254_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21054_ (.A1(net3221),
    .A2(_05255_),
    .B(_04811_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21055_ (.A1(_05075_),
    .A2(_05080_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input129 (.I(irq_external_i),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21057_ (.I0(net96),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05258_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21058_ (.I(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21059_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21060_ (.A1(_05064_),
    .A2(_05258_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21061_ (.I0(_05260_),
    .I1(_05261_),
    .S(net3071),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input128 (.I(instr_rvalid_i),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input127 (.I(instr_rdata_i[9]),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input126 (.I(instr_rdata_i[8]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21065_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .A2(_05092_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input125 (.I(instr_rdata_i[7]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input124 (.I(instr_rdata_i[6]),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21068_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .A2(_05061_),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21069_ (.A1(_01987_),
    .A2(_05074_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input123 (.I(instr_rdata_i[5]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21071_ (.A1(net3071),
    .A2(_05266_),
    .B1(_05269_),
    .B2(_05270_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21072_ (.A1(net3057),
    .A2(_05259_),
    .B1(_05262_),
    .B2(_08736_),
    .C(_05272_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21073_ (.I0(net97),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21074_ (.I(_05273_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21075_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21076_ (.A1(_05064_),
    .A2(_05273_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21077_ (.I0(_05275_),
    .I1(_05276_),
    .S(net3071),
    .Z(_05277_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21078_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .A2(_05092_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21079_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .A2(_05061_),
    .Z(_05279_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21080_ (.A1(net3071),
    .A2(_05278_),
    .B1(_05279_),
    .B2(_05270_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21081_ (.A1(net3057),
    .A2(_05274_),
    .B1(_05277_),
    .B2(_08736_),
    .C(_05280_),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21082_ (.I0(net98),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21083_ (.I(_05281_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21084_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21085_ (.A1(_05064_),
    .A2(_05281_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input122 (.I(instr_rdata_i[4]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21087_ (.I0(_05283_),
    .I1(_05284_),
    .S(net3071),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21088_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .A2(_05092_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21089_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .A2(_05061_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21090_ (.A1(net3071),
    .A2(_05287_),
    .B1(_05288_),
    .B2(_05270_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21091_ (.A1(net3057),
    .A2(_05282_),
    .B1(_05286_),
    .B2(_08736_),
    .C(_05289_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21092_ (.I0(net99),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21093_ (.I(_05290_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21094_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21095_ (.A1(_05064_),
    .A2(_05290_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21096_ (.I0(_05292_),
    .I1(_05293_),
    .S(net3071),
    .Z(_05294_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21097_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .A2(_05092_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21098_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .A2(_05061_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21099_ (.A1(net3071),
    .A2(_05295_),
    .B1(_05296_),
    .B2(_05270_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21100_ (.A1(net3057),
    .A2(_05291_),
    .B1(_05294_),
    .B2(_08736_),
    .C(_05297_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21101_ (.I0(net100),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .S(net3651),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21102_ (.I(_05298_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21103_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21104_ (.A1(_05064_),
    .A2(_05298_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21105_ (.I0(_05300_),
    .I1(_05301_),
    .S(net3071),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21106_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .A2(_05092_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21107_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .A2(_05061_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21108_ (.A1(net3071),
    .A2(_05303_),
    .B1(_05304_),
    .B2(_05270_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21109_ (.A1(net3057),
    .A2(_05299_),
    .B1(_05302_),
    .B2(_08736_),
    .C(_05305_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21110_ (.I0(net101),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .S(net3651),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21111_ (.I(_05306_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21112_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21113_ (.A1(_05064_),
    .A2(_05306_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21114_ (.I0(_05308_),
    .I1(_05309_),
    .S(net3071),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21115_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .A2(_05092_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21116_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .A2(_05061_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21117_ (.A1(net3071),
    .A2(_05311_),
    .B1(_05312_),
    .B2(_05270_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21118_ (.A1(net3057),
    .A2(_05307_),
    .B1(_05310_),
    .B2(_08736_),
    .C(_05313_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21119_ (.I0(net102),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .S(net3651),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21120_ (.I(_05314_),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21121_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21122_ (.A1(_05064_),
    .A2(_05314_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21123_ (.I0(_05316_),
    .I1(_05317_),
    .S(net3071),
    .Z(_05318_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21124_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .A2(_05092_),
    .Z(_05319_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21125_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .A2(_05061_),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21126_ (.A1(net3071),
    .A2(_05319_),
    .B1(_05320_),
    .B2(_05270_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21127_ (.A1(net3057),
    .A2(_05315_),
    .B1(_05318_),
    .B2(_08736_),
    .C(_05321_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _21128_ (.A1(_01987_),
    .A2(_05065_),
    .A3(_05078_),
    .Z(_05322_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input121 (.I(instr_rdata_i[3]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21130_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05324_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input120 (.I(instr_rdata_i[31]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21132_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _21133_ (.A1(net3091),
    .A2(_01958_),
    .A3(_01961_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _21134_ (.A1(_05071_),
    .A2(_05072_),
    .A3(_04364_),
    .A4(_05069_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21135_ (.A1(_05327_),
    .A2(_05328_),
    .B(_05079_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21136_ (.A1(_05326_),
    .A2(net3068),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input119 (.I(instr_rdata_i[30]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input118 (.I(instr_rdata_i[2]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21139_ (.A1(net3652),
    .A2(net103),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input117 (.I(instr_rdata_i[29]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input116 (.I(instr_rdata_i[28]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21142_ (.A1(_08736_),
    .A2(net103),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05336_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input115 (.I(instr_rdata_i[27]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21144_ (.I0(_05333_),
    .I1(_05336_),
    .S(net3071),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21145_ (.A1(_05324_),
    .A2(_05330_),
    .A3(_05338_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21146_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05339_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input114 (.I(instr_rdata_i[26]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21148_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21149_ (.A1(net3068),
    .A2(_05341_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21150_ (.A1(net3652),
    .A2(net104),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21151_ (.A1(_08736_),
    .A2(net104),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21152_ (.I0(_05343_),
    .I1(_05344_),
    .S(net3071),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21153_ (.A1(_05339_),
    .A2(_05342_),
    .A3(_05345_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21154_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05346_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21155_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21156_ (.A1(net3068),
    .A2(_05347_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21157_ (.A1(net3652),
    .A2(net105),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input113 (.I(instr_rdata_i[25]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21159_ (.A1(_08736_),
    .A2(net105),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21160_ (.I0(_05349_),
    .I1(_05351_),
    .S(net3071),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21161_ (.A1(_05346_),
    .A2(_05348_),
    .A3(_05352_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21162_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21163_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21164_ (.A1(net3068),
    .A2(_05354_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input112 (.I(instr_rdata_i[24]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21166_ (.A1(net3652),
    .A2(net106),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21167_ (.A1(_08736_),
    .A2(net106),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21168_ (.I0(_05357_),
    .I1(_05358_),
    .S(net3071),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21169_ (.A1(_05353_),
    .A2(_05355_),
    .A3(_05359_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21170_ (.I0(net107),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05360_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21171_ (.I(_05360_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21172_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input111 (.I(instr_rdata_i[23]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21174_ (.A1(_05064_),
    .A2(_05360_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21175_ (.I0(_05362_),
    .I1(_05364_),
    .S(net3071),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21176_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .A2(_05092_),
    .Z(_05366_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21177_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .A2(_05061_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21178_ (.A1(net3071),
    .A2(_05366_),
    .B1(_05367_),
    .B2(_05270_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21179_ (.A1(net3057),
    .A2(_05361_),
    .B1(_05365_),
    .B2(_08736_),
    .C(_05368_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21180_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21181_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21182_ (.A1(net3068),
    .A2(_05370_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21183_ (.A1(net3652),
    .A2(net108),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05372_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21184_ (.A1(_08736_),
    .A2(net108),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21185_ (.I0(_05372_),
    .I1(_05373_),
    .S(net3071),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21186_ (.A1(_05369_),
    .A2(_05371_),
    .A3(_05374_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21187_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05375_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21188_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21189_ (.A1(net3068),
    .A2(_05376_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input110 (.I(instr_rdata_i[22]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21191_ (.A1(net3652),
    .A2(net109),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A4(_05061_),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21192_ (.A1(_08736_),
    .A2(net109),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A4(_05061_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21193_ (.I0(_05379_),
    .I1(_05380_),
    .S(net3071),
    .Z(_05381_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21194_ (.A1(_05375_),
    .A2(_05377_),
    .A3(_05381_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21195_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21196_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21197_ (.A1(net3068),
    .A2(_05383_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21198_ (.A1(net3652),
    .A2(net110),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A4(_05061_),
    .Z(_05385_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21199_ (.A1(_08736_),
    .A2(net110),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A4(_05061_),
    .Z(_05386_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input109 (.I(instr_rdata_i[21]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21201_ (.I0(_05385_),
    .I1(_05386_),
    .S(net3071),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21202_ (.A1(_05382_),
    .A2(_05384_),
    .A3(_05388_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21203_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05389_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21204_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21205_ (.A1(net3068),
    .A2(_05390_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21206_ (.A1(net3652),
    .A2(net111),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05392_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21207_ (.A1(_08736_),
    .A2(net111),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21208_ (.I0(_05392_),
    .I1(_05393_),
    .S(net3071),
    .Z(_05394_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21209_ (.A1(_05389_),
    .A2(_05391_),
    .A3(_05394_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21210_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21211_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21212_ (.A1(net3068),
    .A2(_05396_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21213_ (.A1(net3652),
    .A2(net112),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21214_ (.A1(_08736_),
    .A2(net112),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21215_ (.I0(_05398_),
    .I1(_05399_),
    .S(net3071),
    .Z(_05400_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21216_ (.A1(_05395_),
    .A2(_05397_),
    .A3(_05400_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21217_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21218_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21219_ (.A1(net3068),
    .A2(_05402_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21220_ (.A1(net3652),
    .A2(net113),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21221_ (.A1(_08736_),
    .A2(net113),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21222_ (.I0(_05404_),
    .I1(_05405_),
    .S(net3071),
    .Z(_05406_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21223_ (.A1(_05401_),
    .A2(_05403_),
    .A3(_05406_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21224_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05407_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21225_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21226_ (.A1(net3068),
    .A2(_05408_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21227_ (.A1(net3652),
    .A2(net114),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21228_ (.A1(_08736_),
    .A2(net114),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21229_ (.I0(_05410_),
    .I1(_05411_),
    .S(net3071),
    .Z(_05412_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21230_ (.A1(_05407_),
    .A2(_05409_),
    .A3(_05412_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21231_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21232_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21233_ (.A1(net3068),
    .A2(_05414_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21234_ (.A1(net3652),
    .A2(net115),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A4(_05061_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21235_ (.A1(_08736_),
    .A2(net115),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A4(_05061_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21236_ (.I0(_05416_),
    .I1(_05417_),
    .S(net3071),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21237_ (.A1(_05413_),
    .A2(_05415_),
    .A3(_05418_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21238_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05419_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21239_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21240_ (.A1(net3068),
    .A2(_05420_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21241_ (.A1(net3652),
    .A2(net116),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A4(_05061_),
    .Z(_05422_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21242_ (.A1(_08736_),
    .A2(net116),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A4(_05061_),
    .Z(_05423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21243_ (.I0(_05422_),
    .I1(_05423_),
    .S(net3071),
    .Z(_05424_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21244_ (.A1(_05419_),
    .A2(_05421_),
    .A3(_05424_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21245_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21246_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21247_ (.A1(net3068),
    .A2(_05426_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21248_ (.A1(net3652),
    .A2(net117),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05428_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21249_ (.A1(_08736_),
    .A2(net117),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21250_ (.I0(_05428_),
    .I1(_05429_),
    .S(net3071),
    .Z(_05430_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21251_ (.A1(_05425_),
    .A2(_05427_),
    .A3(_05430_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21252_ (.I0(net118),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21253_ (.I(_05431_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21254_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21255_ (.A1(_05064_),
    .A2(_05431_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21256_ (.I0(_05433_),
    .I1(_05434_),
    .S(net3071),
    .Z(_05435_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21257_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .A2(_05092_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21258_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .A2(_05061_),
    .Z(_05437_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21259_ (.A1(net3071),
    .A2(_05436_),
    .B1(_05437_),
    .B2(_05270_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21260_ (.A1(net3057),
    .A2(_05432_),
    .B1(_05435_),
    .B2(_08736_),
    .C(_05438_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21261_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21262_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21263_ (.A1(net3068),
    .A2(_05440_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21264_ (.A1(net3652),
    .A2(net119),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05442_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21265_ (.A1(_08736_),
    .A2(net119),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21266_ (.I0(_05442_),
    .I1(_05443_),
    .S(net3071),
    .Z(_05444_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21267_ (.A1(_05439_),
    .A2(_05441_),
    .A3(_05444_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21268_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .A2(_05075_),
    .A3(net3072),
    .A4(_05322_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21269_ (.A1(_05070_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21270_ (.A1(net3068),
    .A2(_05446_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21271_ (.A1(net3652),
    .A2(net120),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21272_ (.A1(_08736_),
    .A2(net120),
    .A3(net3651),
    .A4(_05061_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21273_ (.I0(_05448_),
    .I1(_05449_),
    .S(net3071),
    .Z(_05450_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21274_ (.A1(_05445_),
    .A2(_05447_),
    .A3(_05450_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21275_ (.I0(net96),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21276_ (.I0(_05451_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .S(net3058),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21277_ (.I0(net107),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21278_ (.I0(_05452_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .S(net3058),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21279_ (.I0(net118),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(net3650),
    .Z(_05453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21280_ (.I0(_05453_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .S(net3058),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21281_ (.I0(net121),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(net3650),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21282_ (.I0(_05454_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .S(net3058),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21283_ (.I0(net122),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(net3650),
    .Z(_05455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21284_ (.I0(_05455_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .S(net3058),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21285_ (.I0(net123),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(net3650),
    .Z(_05456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21286_ (.I0(_05456_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .S(net3058),
    .Z(_01672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21287_ (.I0(net124),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(net3650),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21288_ (.I0(_05457_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .S(net3058),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21289_ (.I0(net125),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(net3650),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21290_ (.I0(_05458_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .S(net3058),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21291_ (.I0(net121),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05459_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21292_ (.I(_05459_),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21293_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21294_ (.A1(_05064_),
    .A2(_05459_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21295_ (.I0(_05461_),
    .I1(_05462_),
    .S(net3071),
    .Z(_05463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21296_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .A2(_05092_),
    .Z(_05464_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21297_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .A2(_05061_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21298_ (.A1(net3071),
    .A2(_05464_),
    .B1(_05465_),
    .B2(_05270_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21299_ (.A1(net3057),
    .A2(_05460_),
    .B1(_05463_),
    .B2(_08736_),
    .C(_05466_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input108 (.I(instr_rdata_i[20]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21301_ (.I0(net126),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(net3650),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21302_ (.I0(_05468_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .S(net3058),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21303_ (.I0(net127),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(net3650),
    .Z(_05469_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input107 (.I(instr_rdata_i[1]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21305_ (.I0(_05469_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .S(net3058),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21306_ (.I0(net97),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(net3650),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21307_ (.I0(_05471_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .S(net3058),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21308_ (.I0(net98),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(net3650),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21309_ (.I0(_05472_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .S(net3058),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21310_ (.I0(net99),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(net3650),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21311_ (.I0(_05473_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .S(net3058),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21312_ (.I0(net100),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(net3650),
    .Z(_05474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21313_ (.I0(_05474_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .S(net3058),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21314_ (.I0(net101),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(net3650),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21315_ (.I0(_05475_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .S(net3058),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21316_ (.I0(net102),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(net3650),
    .Z(_05476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21317_ (.I0(_05476_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .S(net3058),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21318_ (.I0(net103),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21319_ (.I0(_05477_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .S(net3059),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21320_ (.I0(net104),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21321_ (.I0(_05478_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .S(net3059),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21322_ (.I0(net122),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05479_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21323_ (.I(_05479_),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21324_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21325_ (.A1(_05064_),
    .A2(_05479_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21326_ (.I0(_05481_),
    .I1(_05482_),
    .S(net3071),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21327_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .A2(_05092_),
    .Z(_05484_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21328_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .A2(_05061_),
    .Z(_05485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21329_ (.A1(net3071),
    .A2(_05484_),
    .B1(_05485_),
    .B2(_05270_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21330_ (.A1(net3057),
    .A2(_05480_),
    .B1(_05483_),
    .B2(_08736_),
    .C(_05486_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input106 (.I(instr_rdata_i[19]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21332_ (.I0(net105),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21333_ (.I0(_05488_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .S(net3059),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21334_ (.I0(net106),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(net3650),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input105 (.I(instr_rdata_i[18]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21336_ (.I0(_05489_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .S(net3059),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21337_ (.I0(net108),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(net3650),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21338_ (.I0(_05491_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .S(net3059),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21339_ (.I0(net109),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(net3650),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21340_ (.I0(_05492_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .S(net3058),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21341_ (.I0(net110),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(net3650),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21342_ (.I0(_05493_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .S(net3058),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21343_ (.I0(net111),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21344_ (.I0(_05494_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .S(net3059),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21345_ (.I0(net112),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21346_ (.I0(_05495_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .S(net3059),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21347_ (.I0(net113),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21348_ (.I0(_05496_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .S(net3059),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21349_ (.I0(net114),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(net3650),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21350_ (.I0(_05497_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .S(net3059),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21351_ (.I0(net115),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(net3650),
    .Z(_05498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21352_ (.I0(_05498_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .S(net3058),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21353_ (.I0(net123),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21354_ (.I(_05499_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21355_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .ZN(_05501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21356_ (.A1(_05064_),
    .A2(_05499_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21357_ (.I0(_05501_),
    .I1(_05502_),
    .S(net3071),
    .Z(_05503_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21358_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .A2(_05092_),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21359_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .A2(_05061_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21360_ (.A1(net3071),
    .A2(_05504_),
    .B1(_05505_),
    .B2(_05270_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21361_ (.A1(net3057),
    .A2(_05500_),
    .B1(_05503_),
    .B2(_08736_),
    .C(_05506_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21362_ (.I0(net116),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(net3650),
    .Z(_05507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21363_ (.I0(_05507_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .S(net3058),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21364_ (.I0(net117),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21365_ (.I0(_05508_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .S(net3059),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21366_ (.I0(net119),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21367_ (.I0(_05509_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .S(net3059),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21368_ (.I0(net120),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(_05510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21369_ (.I0(_05510_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .S(net3059),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21370_ (.I0(net96),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(_05105_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21371_ (.I0(net107),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(_05105_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21372_ (.I0(net118),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(_05105_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21373_ (.I0(net121),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(_05105_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21374_ (.I0(net122),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(_05105_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21375_ (.I0(net123),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(_05105_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21376_ (.I0(net124),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21377_ (.I(_05511_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21378_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21379_ (.A1(_05064_),
    .A2(_05511_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21380_ (.I0(_05513_),
    .I1(_05514_),
    .S(net3071),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21381_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .A2(_05092_),
    .Z(_05516_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21382_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .A2(_05061_),
    .Z(_05517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21383_ (.A1(net3071),
    .A2(_05516_),
    .B1(_05517_),
    .B2(_05270_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21384_ (.A1(net3057),
    .A2(_05512_),
    .B1(_05515_),
    .B2(_08736_),
    .C(_05518_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21385_ (.I0(net124),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(_05105_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21386_ (.I0(net125),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(_05105_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21387_ (.I0(net126),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(_05105_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input104 (.I(instr_rdata_i[17]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21389_ (.I0(net127),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(_05105_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21390_ (.I0(net97),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(_05105_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21391_ (.I0(net98),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(_05105_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21392_ (.I0(net99),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(_05105_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21393_ (.I0(net100),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(_05105_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21394_ (.I0(net101),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(_05105_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21395_ (.I0(net102),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(_05105_),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21396_ (.I0(net125),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .S(net3651),
    .Z(_05520_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21397_ (.I(_05520_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21398_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21399_ (.A1(_05064_),
    .A2(_05520_),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21400_ (.I0(_05522_),
    .I1(_05523_),
    .S(net3071),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21401_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .A2(_05092_),
    .Z(_05525_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21402_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .A2(_05061_),
    .Z(_05526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21403_ (.A1(net3071),
    .A2(_05525_),
    .B1(_05526_),
    .B2(_05270_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21404_ (.A1(net3057),
    .A2(_05521_),
    .B1(_05524_),
    .B2(_08736_),
    .C(_05527_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21405_ (.I0(net103),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(_05105_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21406_ (.I0(net104),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(_05105_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21407_ (.I0(net105),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(_05105_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input103 (.I(instr_rdata_i[16]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21409_ (.I0(net106),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(_05105_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21410_ (.I0(net108),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(_05105_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21411_ (.I0(net109),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(_05105_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21412_ (.I0(net110),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(_05105_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21413_ (.I0(net111),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(_05105_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21414_ (.I0(net112),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(_05105_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21415_ (.I0(net113),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(_05105_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21416_ (.I0(net126),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05529_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21417_ (.I(_05529_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21418_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21419_ (.A1(_05064_),
    .A2(_05529_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21420_ (.I0(_05531_),
    .I1(_05532_),
    .S(net3071),
    .Z(_05533_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21421_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .A2(_05092_),
    .Z(_05534_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21422_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .A2(_05061_),
    .Z(_05535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21423_ (.A1(net3071),
    .A2(_05534_),
    .B1(_05535_),
    .B2(_05270_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21424_ (.A1(net3057),
    .A2(_05530_),
    .B1(_05533_),
    .B2(_08736_),
    .C(_05536_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21425_ (.I0(net114),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(_05105_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21426_ (.I0(net115),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(_05105_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21427_ (.I0(net116),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(_05105_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21428_ (.I0(net117),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(_05105_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21429_ (.I0(net119),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(_05105_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21430_ (.I0(net120),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(_05105_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21431_ (.I0(net127),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21432_ (.I(_05537_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21433_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21434_ (.A1(_05064_),
    .A2(_05537_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21435_ (.I0(_05539_),
    .I1(_05540_),
    .S(net3071),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21436_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .A2(_05092_),
    .Z(_05542_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21437_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .A2(_05061_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21438_ (.A1(net3071),
    .A2(_05542_),
    .B1(_05543_),
    .B2(_05270_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21439_ (.A1(net3057),
    .A2(_05538_),
    .B1(_05541_),
    .B2(_08736_),
    .C(_05544_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input102 (.I(instr_rdata_i[15]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21441_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .I1(_04826_),
    .S(_08869_),
    .Z(net219));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _21442_ (.I(net95),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21443_ (.A1(_05546_),
    .A2(_11661_[0]),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input101 (.I(instr_rdata_i[14]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21445_ (.I0(net219),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .S(_05547_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21446_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .I1(_04822_),
    .S(_08869_),
    .Z(net220));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21447_ (.I0(net220),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .S(_05547_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21448_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .I1(_04850_),
    .S(_08869_),
    .Z(net221));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21449_ (.I0(net221),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .S(_05547_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21450_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .I1(_04849_),
    .S(_08869_),
    .Z(net222));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21451_ (.I0(net222),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .S(_05547_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21452_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .I1(_04873_),
    .S(_08869_),
    .Z(net223));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21453_ (.I0(net223),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .S(_05547_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21454_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .I1(_04871_),
    .S(_08869_),
    .Z(net224));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21455_ (.I0(net224),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .S(_05547_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21456_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .I1(_04882_),
    .S(_08869_),
    .Z(net225));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21457_ (.I0(net225),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .S(_05547_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21458_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .I1(_04891_),
    .S(_08869_),
    .Z(net226));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21459_ (.I0(net226),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .S(_05547_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21460_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .I1(_04901_),
    .S(_08869_),
    .Z(net227));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21461_ (.I0(net227),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .S(_05547_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21462_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .I1(_04910_),
    .S(_08869_),
    .Z(net228));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21463_ (.I0(net228),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .S(_05547_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input100 (.I(instr_rdata_i[13]),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21465_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .I1(_04924_),
    .S(_08869_),
    .Z(net229));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input99 (.I(instr_rdata_i[12]),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21467_ (.I0(net229),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .S(_05547_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21468_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .I1(_04932_),
    .S(_08869_),
    .Z(net230));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21469_ (.I0(net230),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .S(_05547_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21470_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .I1(_04942_),
    .S(_08869_),
    .Z(net231));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21471_ (.I0(net231),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .S(_05547_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21472_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .I1(_04953_),
    .S(_08869_),
    .Z(net232));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21473_ (.I0(net232),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .S(_05547_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21474_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .I1(_04976_),
    .S(_08869_),
    .Z(net233));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21475_ (.I0(net233),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .S(_05547_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21476_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .I1(_04975_),
    .S(_08869_),
    .Z(net234));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21477_ (.I0(net234),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .S(_05547_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21478_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .I1(_04997_),
    .S(_08869_),
    .Z(net235));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21479_ (.I0(net235),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .S(_05547_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21480_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .I1(_05009_),
    .S(_08869_),
    .Z(net236));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21481_ (.I0(net236),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .S(_05547_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21482_ (.I(_05008_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21483_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .I1(_05551_),
    .S(_08869_),
    .Z(net237));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21484_ (.I0(net237),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .S(_05547_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21485_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .I1(_05018_),
    .S(_08869_),
    .Z(net238));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21486_ (.I0(net238),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .S(_05547_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input98 (.I(instr_rdata_i[11]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21488_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .I1(_11660_[0]),
    .S(_08869_),
    .Z(net239));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input97 (.I(instr_rdata_i[10]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21490_ (.I0(net239),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .S(_05547_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21491_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .I1(_05028_),
    .S(_08869_),
    .Z(net240));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21492_ (.I0(net240),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .S(_05547_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21493_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .I1(_05038_),
    .S(_08869_),
    .Z(net241));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21494_ (.I0(net241),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .S(_05547_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21495_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .I1(_11663_[0]),
    .S(_08869_),
    .Z(net242));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21496_ (.I0(net242),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .S(_05547_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21497_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .I1(_05041_),
    .S(_08869_),
    .Z(net243));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21498_ (.I0(net243),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .S(_05547_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21499_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .I1(_05045_),
    .S(_08869_),
    .Z(net244));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21500_ (.I0(net244),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .S(_05547_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21501_ (.I(_04793_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21502_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .I1(_05554_),
    .S(_08869_),
    .Z(net245));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21503_ (.I0(net245),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .S(_05547_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21504_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .I1(_04799_),
    .S(_08869_),
    .Z(net246));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21505_ (.I0(net246),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .S(_05547_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21506_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .I1(_04778_),
    .S(_08869_),
    .Z(net247));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21507_ (.I0(net247),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .S(_05547_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21508_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .I1(_04769_),
    .S(_08869_),
    .Z(net248));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21509_ (.I0(net248),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .S(_05547_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21510_ (.A1(_06232_),
    .A2(net26),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21511_ (.A1(_06231_),
    .A2(net59),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _21512_ (.I(_05556_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21513_ (.A1(_08397_),
    .A2(_05557_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input96 (.I(instr_rdata_i[0]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21515_ (.A1(_08398_),
    .A2(_08885_),
    .B1(_05558_),
    .B2(\load_store_unit_i.ls_fsm_cs[1] ),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21516_ (.A1(_08885_),
    .A2(_08886_),
    .B1(_05558_),
    .B2(net3472),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _21517_ (.A1(_05555_),
    .A2(_05560_),
    .B1(_05561_),
    .B2(\load_store_unit_i.ls_fsm_cs[1] ),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input95 (.I(instr_gnt_i),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21519_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .I1(\alu_adder_result_ex[0] ),
    .S(_05562_),
    .Z(_01851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21520_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .I1(net151),
    .S(net3198),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21521_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .I1(net152),
    .S(net3198),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21522_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .I1(net153),
    .S(net3198),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21523_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .I1(net154),
    .S(net3198),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21524_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .I1(net364),
    .S(net3198),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21525_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .I1(net156),
    .S(net3198),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21526_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .I1(net403),
    .S(net3198),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21527_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .I1(net158),
    .S(net3198),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21528_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .I1(net360),
    .S(net3198),
    .Z(_01860_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input94 (.I(instr_err_i),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21530_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .I1(net160),
    .S(net3198),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21531_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .I1(\alu_adder_result_ex[1] ),
    .S(_05562_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21532_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .I1(net161),
    .S(net3198),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21533_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .I1(net162),
    .S(net3198),
    .Z(_01864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21534_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .I1(net163),
    .S(net3198),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21535_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .I1(net164),
    .S(net3198),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21536_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .I1(net165),
    .S(net3198),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21537_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .I1(net166),
    .S(net3198),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21538_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .I1(net167),
    .S(net3198),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21539_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .I1(net367),
    .S(net3198),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input93 (.I(hart_id_i[9]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21541_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .I1(net169),
    .S(net3198),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21542_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .I1(net338),
    .S(net3198),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21543_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .I1(net171),
    .S(_05562_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21544_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .I1(net256),
    .S(net3198),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21545_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .I1(net173),
    .S(_05562_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21546_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .I1(net174),
    .S(_05562_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21547_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .I1(net175),
    .S(_05562_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21548_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .I1(net176),
    .S(_05562_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21549_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .I1(net177),
    .S(net3198),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21550_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .I1(net178),
    .S(_05562_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21551_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .I1(net179),
    .S(net3198),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21552_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .I1(net180),
    .S(net3198),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21553_ (.A1(_06220_),
    .A2(net3417),
    .A3(_08880_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21554_ (.I0(_05566_),
    .I1(\load_store_unit_i.data_sign_ext_q ),
    .S(_08887_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21555_ (.A1(_06411_),
    .A2(_06757_),
    .A3(_06782_),
    .Z(net218));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21556_ (.I0(net218),
    .I1(\load_store_unit_i.data_we_q ),
    .S(_08887_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21557_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_08883_),
    .B(net26),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21558_ (.A1(net26),
    .A2(_05557_),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21559_ (.A1(_05567_),
    .A2(_05568_),
    .B(net3472),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21560_ (.A1(_06231_),
    .A2(_06340_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input92 (.I(hart_id_i[8]),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21562_ (.A1(net320),
    .A2(_11647_[0]),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21563_ (.A1(_06744_),
    .A2(_08880_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21564_ (.I0(_05572_),
    .I1(_08425_),
    .S(_05573_),
    .Z(_05574_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21565_ (.A1(net26),
    .A2(_05556_),
    .B(_06232_),
    .C(\load_store_unit_i.ls_fsm_cs[1] ),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21566_ (.A1(_05570_),
    .A2(_05574_),
    .B(_05575_),
    .C(_05569_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21567_ (.A1(_11641_[0]),
    .A2(_05569_),
    .B(_05576_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21568_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(net59),
    .B(_08884_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21569_ (.A1(_06231_),
    .A2(_05577_),
    .B(net26),
    .C(net3472),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21570_ (.A1(net26),
    .A2(_05574_),
    .B(\load_store_unit_i.ls_fsm_cs[0] ),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21571_ (.I0(_05556_),
    .I1(_05574_),
    .S(_06340_),
    .Z(_05579_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21572_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(_05578_),
    .B1(_05579_),
    .B2(net26),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21573_ (.A1(_06232_),
    .A2(_05580_),
    .Z(_05581_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21574_ (.I(net59),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21575_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(_05582_),
    .B(\load_store_unit_i.ls_fsm_cs[0] ),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21576_ (.I0(net59),
    .I1(_08883_),
    .S(_06232_),
    .Z(_05584_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _21577_ (.A1(net3472),
    .A2(net26),
    .A3(_05583_),
    .B1(_05584_),
    .B2(_05570_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21578_ (.I0(_05581_),
    .I1(\load_store_unit_i.ls_fsm_cs[1] ),
    .S(_05585_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21579_ (.I0(net3472),
    .I1(_08886_),
    .S(\load_store_unit_i.ls_fsm_cs[1] ),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21580_ (.A1(_06231_),
    .A2(_05582_),
    .A3(_05586_),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21581_ (.A1(net3472),
    .A2(\load_store_unit_i.ls_fsm_cs[1] ),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21582_ (.A1(_05557_),
    .A2(_05587_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21583_ (.A1(_06340_),
    .A2(net59),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21584_ (.I0(_05577_),
    .I1(_05589_),
    .S(net3472),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21585_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_05590_),
    .B(\load_store_unit_i.lsu_err_q ),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21586_ (.A1(_08397_),
    .A2(_05588_),
    .B(_05591_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21587_ (.I0(\alu_adder_result_ex[0] ),
    .I1(\load_store_unit_i.rdata_offset_q[0] ),
    .S(_08887_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21588_ (.I0(\alu_adder_result_ex[1] ),
    .I1(\load_store_unit_i.rdata_offset_q[1] ),
    .S(_08887_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21589_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_05588_),
    .Z(_05592_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input91 (.I(hart_id_i[7]),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21591_ (.I0(net57),
    .I1(\load_store_unit_i.rdata_q[0] ),
    .S(_05592_),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21592_ (.I0(net36),
    .I1(\load_store_unit_i.rdata_q[10] ),
    .S(_05592_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21593_ (.I0(net37),
    .I1(\load_store_unit_i.rdata_q[11] ),
    .S(_05592_),
    .Z(_01894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21594_ (.I0(net39),
    .I1(\load_store_unit_i.rdata_q[12] ),
    .S(_05592_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21595_ (.I0(net40),
    .I1(\load_store_unit_i.rdata_q[13] ),
    .S(_05592_),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21596_ (.I0(net41),
    .I1(\load_store_unit_i.rdata_q[14] ),
    .S(_05592_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21597_ (.I0(net42),
    .I1(\load_store_unit_i.rdata_q[15] ),
    .S(_05592_),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21598_ (.I0(net43),
    .I1(\load_store_unit_i.rdata_q[16] ),
    .S(_05592_),
    .Z(_01899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21599_ (.I0(net44),
    .I1(\load_store_unit_i.rdata_q[17] ),
    .S(_05592_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21600_ (.I0(net45),
    .I1(\load_store_unit_i.rdata_q[18] ),
    .S(_05592_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input90 (.I(hart_id_i[6]),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21602_ (.I0(net46),
    .I1(\load_store_unit_i.rdata_q[19] ),
    .S(_05592_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21603_ (.I0(net58),
    .I1(\load_store_unit_i.rdata_q[1] ),
    .S(_05592_),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21604_ (.I0(net47),
    .I1(\load_store_unit_i.rdata_q[20] ),
    .S(_05592_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21605_ (.I0(net48),
    .I1(\load_store_unit_i.rdata_q[21] ),
    .S(_05592_),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21606_ (.I0(net50),
    .I1(\load_store_unit_i.rdata_q[22] ),
    .S(_05592_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21607_ (.I0(net51),
    .I1(\load_store_unit_i.rdata_q[23] ),
    .S(_05592_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21608_ (.I0(net28),
    .I1(\load_store_unit_i.rdata_q[2] ),
    .S(_05592_),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21609_ (.I0(net29),
    .I1(\load_store_unit_i.rdata_q[3] ),
    .S(_05592_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21610_ (.I0(net30),
    .I1(\load_store_unit_i.rdata_q[4] ),
    .S(_05592_),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21611_ (.I0(net31),
    .I1(\load_store_unit_i.rdata_q[5] ),
    .S(_05592_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21612_ (.I0(net32),
    .I1(\load_store_unit_i.rdata_q[6] ),
    .S(_05592_),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21613_ (.I0(net33),
    .I1(\load_store_unit_i.rdata_q[7] ),
    .S(_05592_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21614_ (.I0(net34),
    .I1(\load_store_unit_i.rdata_q[8] ),
    .S(_05592_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21615_ (.I0(net35),
    .I1(\load_store_unit_i.rdata_q[9] ),
    .S(_05592_),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _21616_ (.A1(_04386_),
    .A2(_02535_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21617_ (.A1(_02217_),
    .A2(_02221_),
    .A3(_02678_),
    .B(_05595_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21618_ (.I(\cs_registers_i.mstatus_q[2] ),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21619_ (.A1(_05597_),
    .A2(_02678_),
    .Z(_05598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21620_ (.A1(\cs_registers_i.priv_mode_id_o[0] ),
    .A2(_02535_),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_q[0] ),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21621_ (.A1(_05596_),
    .A2(_05598_),
    .B(_05599_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21622_ (.A1(\cs_registers_i.priv_mode_id_o[1] ),
    .A2(_02535_),
    .B1(_02537_),
    .B2(\cs_registers_i.mstack_q[1] ),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21623_ (.I(\cs_registers_i.mstatus_q[3] ),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21624_ (.A1(_05601_),
    .A2(_02678_),
    .A3(_05595_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21625_ (.A1(_05596_),
    .A2(_05600_),
    .B(_05602_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21626_ (.A1(_08638_),
    .A2(\cs_registers_i.mstack_q[2] ),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21627_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(_02535_),
    .B1(_05603_),
    .B2(_04386_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21628_ (.A1(\cs_registers_i.mstatus_q[4] ),
    .A2(_02678_),
    .A3(_05595_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21629_ (.A1(_09593_),
    .A2(_02678_),
    .B(_05604_),
    .C(_05605_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21630_ (.A1(\cs_registers_i.mstatus_q[4] ),
    .A2(_04386_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21631_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(_02678_),
    .A3(_05595_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21632_ (.A1(_09491_),
    .A2(_02678_),
    .B(_05606_),
    .C(_05607_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21633_ (.I0(net104),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(net3652),
    .Z(_05608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21634_ (.I0(net107),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input89 (.I(hart_id_i[5]),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21636_ (.I0(_05608_),
    .I1(_05609_),
    .S(_08730_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input88 (.I(hart_id_i[4]),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input87 (.I(hart_id_i[3]),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21639_ (.I0(net112),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(net3652),
    .Z(_05614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21640_ (.I0(net126),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21641_ (.I0(_05614_),
    .I1(_05615_),
    .S(_08730_),
    .Z(_05616_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21642_ (.I(_05616_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21643_ (.I0(net115),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(net3652),
    .Z(_05618_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input86 (.I(hart_id_i[31]),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21645_ (.I0(net98),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21646_ (.I0(_05618_),
    .I1(_05620_),
    .S(_08730_),
    .Z(_05621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21647_ (.I0(net114),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S(net3652),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21648_ (.I0(net97),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21649_ (.I0(_05622_),
    .I1(_05623_),
    .S(_08730_),
    .Z(_05624_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21650_ (.A1(_05621_),
    .A2(_05624_),
    .Z(_05625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21651_ (.I0(net113),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .S(net3652),
    .Z(_05626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21652_ (.I0(net127),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21653_ (.I0(_05626_),
    .I1(_05627_),
    .S(_08730_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input85 (.I(hart_id_i[30]),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21655_ (.I0(net111),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S(net3652),
    .Z(_05630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21656_ (.I0(net125),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21657_ (.I0(_05630_),
    .I1(_05631_),
    .S(_08730_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input84 (.I(hart_id_i[2]),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _21659_ (.A1(_05625_),
    .A2(_05628_),
    .A3(_05632_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21660_ (.A1(_05617_),
    .A2(_05634_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21661_ (.I0(net103),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .S(net3652),
    .Z(_05636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21662_ (.I0(net96),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21663_ (.I0(_05636_),
    .I1(_05637_),
    .S(_08730_),
    .Z(_05638_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input83 (.I(hart_id_i[29]),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21665_ (.I0(net116),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(net3652),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21666_ (.I0(net99),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21667_ (.I0(_05640_),
    .I1(_05641_),
    .S(_08730_),
    .Z(_05642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21668_ (.I0(net110),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(net3652),
    .Z(_05643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21669_ (.I0(net124),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21670_ (.I0(_05643_),
    .I1(_05644_),
    .S(_08730_),
    .Z(_05645_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input82 (.I(hart_id_i[28]),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21672_ (.I0(net109),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(net3652),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21673_ (.I0(net123),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21674_ (.I0(_05647_),
    .I1(_05648_),
    .S(_08730_),
    .Z(_05649_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21675_ (.A1(_05645_),
    .A2(_05649_),
    .Z(_05650_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21676_ (.A1(_05642_),
    .A2(_05650_),
    .Z(_05651_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21677_ (.A1(_05638_),
    .A2(_05651_),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21678_ (.I0(net120),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .S(net3652),
    .Z(_05653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21679_ (.I0(net102),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05654_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21680_ (.A1(_08730_),
    .A2(_05654_),
    .Z(_05655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21681_ (.A1(net3653),
    .A2(_05653_),
    .B(_05655_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21682_ (.I0(net117),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .S(net3652),
    .Z(_05657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21683_ (.I0(net100),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05658_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21684_ (.A1(_08730_),
    .A2(_05658_),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21685_ (.A1(net3653),
    .A2(_05657_),
    .B(_05659_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21686_ (.A1(_05656_),
    .A2(_05660_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21687_ (.A1(_05635_),
    .A2(_05652_),
    .B(_05661_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21688_ (.A1(_08730_),
    .A2(_05641_),
    .Z(_05663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21689_ (.A1(net3653),
    .A2(_05640_),
    .B(_05663_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21690_ (.I0(net108),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(net3652),
    .Z(_05665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21691_ (.I0(net122),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21692_ (.I0(_05665_),
    .I1(_05666_),
    .S(_08730_),
    .Z(_05667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21693_ (.I0(net105),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .S(net3652),
    .Z(_05668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21694_ (.I0(net118),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21695_ (.I0(_05668_),
    .I1(_05669_),
    .S(_08730_),
    .Z(_05670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21696_ (.I0(net106),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .S(net3652),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21697_ (.I0(net121),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21698_ (.I0(_05671_),
    .I1(_05672_),
    .S(_08730_),
    .Z(_05673_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input81 (.I(hart_id_i[27]),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _21700_ (.A1(_05650_),
    .A2(_05670_),
    .A3(_05673_),
    .Z(_05675_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _21701_ (.A1(_05667_),
    .A2(_05675_),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input80 (.I(hart_id_i[26]),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21703_ (.I0(net119),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .S(net3652),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21704_ (.I0(net101),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21705_ (.I0(_05678_),
    .I1(_05679_),
    .S(_08730_),
    .Z(_05680_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input79 (.I(hart_id_i[25]),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21707_ (.A1(_05656_),
    .A2(_05680_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21708_ (.A1(_05660_),
    .A2(_05682_),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21709_ (.A1(_05664_),
    .A2(_05676_),
    .A3(_05683_),
    .Z(_05684_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input78 (.I(hart_id_i[24]),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21711_ (.A1(_08730_),
    .A2(_05623_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21712_ (.A1(net3653),
    .A2(_05622_),
    .B(_05686_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21713_ (.A1(_05621_),
    .A2(_05687_),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21714_ (.I0(_05653_),
    .I1(_05654_),
    .S(_08730_),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21715_ (.A1(_05689_),
    .A2(_05660_),
    .Z(_05690_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21716_ (.A1(_08730_),
    .A2(_05679_),
    .Z(_05691_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21717_ (.A1(net3653),
    .A2(_05678_),
    .B(_05691_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input77 (.I(hart_id_i[23]),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input76 (.I(hart_id_i[22]),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21720_ (.A1(_05692_),
    .A2(_05642_),
    .Z(_05695_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21721_ (.A1(_05688_),
    .A2(_05690_),
    .A3(_05695_),
    .Z(_05696_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21722_ (.A1(_05684_),
    .A2(_05696_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21723_ (.A1(net3395),
    .A2(_05660_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21724_ (.A1(_08730_),
    .A2(_05637_),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21725_ (.A1(net3653),
    .A2(_05636_),
    .B(_05699_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input75 (.I(hart_id_i[21]),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21727_ (.I0(_05697_),
    .I1(_05698_),
    .S(_05700_),
    .Z(_05702_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input74 (.I(hart_id_i[20]),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21729_ (.A1(_05656_),
    .A2(_05660_),
    .Z(_05704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21730_ (.A1(_05692_),
    .A2(_05704_),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input73 (.I(hart_id_i[1]),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21732_ (.A1(_05611_),
    .A2(_05700_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input72 (.I(hart_id_i[19]),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input71 (.I(hart_id_i[18]),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input70 (.I(hart_id_i[17]),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input69 (.I(hart_id_i[16]),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input68 (.I(hart_id_i[15]),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21738_ (.A1(_05692_),
    .A2(_05664_),
    .A3(_05676_),
    .Z(_05713_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21739_ (.A1(_05656_),
    .A2(_05713_),
    .B(_05635_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input67 (.I(hart_id_i[14]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21741_ (.A1(_05689_),
    .A2(_05680_),
    .B(_05714_),
    .C(_05660_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21742_ (.A1(_05642_),
    .A2(_05705_),
    .B(_05707_),
    .C(_05716_),
    .ZN(_05717_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21743_ (.A1(_05611_),
    .A2(_05662_),
    .A3(_05702_),
    .B(_05717_),
    .ZN(_05718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21744_ (.I0(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .I1(_05718_),
    .S(net3069),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21745_ (.A1(net94),
    .A2(_08743_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21746_ (.A1(_05070_),
    .A2(_05719_),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21747_ (.A1(net3653),
    .A2(_05720_),
    .B(_08744_),
    .ZN(_05721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21748_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .A2(_08745_),
    .ZN(_05722_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21749_ (.A1(net3653),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A3(_05083_),
    .A4(_05722_),
    .Z(_05723_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21750_ (.A1(_05721_),
    .A2(_05723_),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21751_ (.I0(\id_stage_i.controller_i.instr_fetch_err_i ),
    .I1(_05724_),
    .S(net3070),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input66 (.I(hart_id_i[13]),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21753_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .A2(_05070_),
    .A3(net94),
    .Z(_05726_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21754_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .B(_05726_),
    .ZN(_05727_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21755_ (.A1(_08730_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .A3(_05727_),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input65 (.I(hart_id_i[12]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21757_ (.I0(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .I1(_05728_),
    .S(net3070),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21758_ (.A1(_05611_),
    .A2(_05638_),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21759_ (.I0(\id_stage_i.controller_i.instr_is_compressed_i ),
    .I1(_05730_),
    .S(net3069),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21760_ (.I0(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .I1(_05638_),
    .S(net3069),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input64 (.I(hart_id_i[11]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21762_ (.I0(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .I1(_05624_),
    .S(net3069),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21763_ (.I0(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .I1(_05621_),
    .S(net3069),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21764_ (.I0(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .I1(_05642_),
    .S(net3069),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21765_ (.I0(_05657_),
    .I1(_05658_),
    .S(_08730_),
    .Z(_05732_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input63 (.I(hart_id_i[10]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input62 (.I(hart_id_i[0]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input61 (.I(fetch_enable_i),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21769_ (.I0(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .I1(_05732_),
    .S(net3069),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21770_ (.I0(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .I1(net3395),
    .S(net3069),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21771_ (.I0(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .I1(_05689_),
    .S(net3069),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21772_ (.I0(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .I1(_05611_),
    .S(net3069),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input60 (.I(debug_req_i),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input59 (.I(data_rvalid_i),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21775_ (.I0(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .I1(_05670_),
    .S(net3069),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21776_ (.I0(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .I1(_05673_),
    .S(net3069),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input58 (.I(data_rdata_i[9]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21778_ (.I0(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .I1(_05667_),
    .S(net3069),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input57 (.I(data_rdata_i[8]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21780_ (.I0(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .I1(_05649_),
    .S(net3069),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21781_ (.I0(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .I1(_05645_),
    .S(net3069),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21782_ (.I0(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .I1(_05632_),
    .S(net3069),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input56 (.I(data_rdata_i[7]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21784_ (.I0(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .I1(_05616_),
    .S(net3069),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21785_ (.I0(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .I1(_05628_),
    .S(net3069),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21786_ (.A1(_08730_),
    .A2(_05609_),
    .Z(_05741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21787_ (.A1(net3653),
    .A2(_05608_),
    .B(_05741_),
    .ZN(_05742_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input55 (.I(data_rdata_i[6]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21789_ (.A1(_05689_),
    .A2(_05692_),
    .Z(_05744_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21790_ (.A1(_05742_),
    .A2(_05744_),
    .B(_05732_),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21791_ (.A1(_05638_),
    .A2(_05745_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21792_ (.I0(\id_stage_i.controller_i.instr_i[0] ),
    .I1(_05746_),
    .S(net3069),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21793_ (.A1(_05692_),
    .A2(_05732_),
    .Z(_05747_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21794_ (.A1(_05660_),
    .A2(_05638_),
    .A3(_05744_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21795_ (.A1(_05624_),
    .A2(_05704_),
    .B(_05700_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21796_ (.A1(_05687_),
    .A2(_05747_),
    .B(_05748_),
    .C(_05749_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input54 (.I(data_rdata_i[5]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21798_ (.A1(_05692_),
    .A2(_05690_),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21799_ (.A1(_05676_),
    .A2(_05752_),
    .Z(_05753_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21800_ (.A1(_05700_),
    .A2(_05753_),
    .B(_05687_),
    .ZN(_05754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21801_ (.I0(_05750_),
    .I1(_05754_),
    .S(_05611_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21802_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .I1(_05755_),
    .S(net3069),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21803_ (.I0(_05704_),
    .I1(_05753_),
    .S(_05611_),
    .Z(_05756_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21804_ (.A1(_05621_),
    .A2(_05624_),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21805_ (.A1(_05642_),
    .A2(_05757_),
    .ZN(_05758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21806_ (.A1(_05689_),
    .A2(_05758_),
    .B(_05732_),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21807_ (.A1(_05742_),
    .A2(_05638_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input53 (.I(data_rdata_i[4]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21809_ (.A1(net3395),
    .A2(_05759_),
    .A3(_05760_),
    .B(_05621_),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21810_ (.A1(_05700_),
    .A2(_05756_),
    .B(_05762_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input52 (.I(data_rdata_i[3]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21812_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .I1(_05763_),
    .S(net3069),
    .Z(_01790_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21813_ (.A1(_05611_),
    .A2(_05700_),
    .ZN(_05765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21814_ (.A1(net3395),
    .A2(_05660_),
    .ZN(_05766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21815_ (.A1(_05661_),
    .A2(_05766_),
    .ZN(_05767_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21816_ (.A1(_05742_),
    .A2(_05700_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _21817_ (.A1(_05767_),
    .A2(_05768_),
    .B(_05730_),
    .ZN(_05769_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _21818_ (.A1(_05732_),
    .A2(_05707_),
    .B(_05769_),
    .ZN(_05770_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input51 (.I(data_rdata_i[31]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21820_ (.A1(_05616_),
    .A2(_05634_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21821_ (.A1(_05670_),
    .A2(_05772_),
    .B(_05682_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input50 (.I(data_rdata_i[30]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21823_ (.A1(_05692_),
    .A2(_05732_),
    .ZN(_05775_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21824_ (.A1(_05621_),
    .A2(_05624_),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21825_ (.A1(_05664_),
    .A2(_05645_),
    .Z(_05777_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21826_ (.A1(_05649_),
    .A2(_05777_),
    .Z(_05778_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21827_ (.A1(_05732_),
    .A2(_05776_),
    .A3(_05778_),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21828_ (.A1(_05775_),
    .A2(_05779_),
    .B(_05642_),
    .ZN(_05780_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21829_ (.A1(_05760_),
    .A2(_05767_),
    .A3(_05773_),
    .A4(_05780_),
    .Z(_05781_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21830_ (.A1(_05765_),
    .A2(_05705_),
    .B1(_05770_),
    .B2(_05664_),
    .C(_05781_),
    .ZN(_05782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21831_ (.I0(\id_stage_i.controller_i.instr_i[12] ),
    .I1(_05782_),
    .S(net3069),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21832_ (.A1(_05611_),
    .A2(_05638_),
    .Z(_05783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21833_ (.A1(_05689_),
    .A2(_05638_),
    .B(_05680_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21834_ (.A1(_05783_),
    .A2(_05784_),
    .Z(_05785_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21835_ (.A1(_05742_),
    .A2(_05638_),
    .Z(_05786_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input49 (.I(data_rdata_i[2]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21837_ (.A1(_05656_),
    .A2(_05680_),
    .A3(_05673_),
    .A4(_05772_),
    .Z(_05788_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21838_ (.A1(_05695_),
    .A2(_05788_),
    .B(_05732_),
    .ZN(_05789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21839_ (.A1(_05621_),
    .A2(_05752_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21840_ (.A1(_05687_),
    .A2(_05777_),
    .B(_05790_),
    .ZN(_05791_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21841_ (.A1(_05786_),
    .A2(_05789_),
    .A3(_05791_),
    .Z(_05792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21842_ (.A1(_05660_),
    .A2(_05785_),
    .B(_05792_),
    .ZN(_05793_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21843_ (.I0(\id_stage_i.controller_i.instr_i[13] ),
    .I1(_05793_),
    .S(net3069),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21844_ (.A1(_05660_),
    .A2(_05700_),
    .Z(_05794_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21845_ (.A1(_05683_),
    .A2(_05772_),
    .Z(_05795_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21846_ (.A1(_05689_),
    .A2(_05660_),
    .ZN(_05796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21847_ (.A1(_05664_),
    .A2(_05650_),
    .B(_05776_),
    .ZN(_05797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21848_ (.A1(_05642_),
    .A2(_05732_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21849_ (.A1(_05796_),
    .A2(_05797_),
    .B(_05798_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21850_ (.A1(_05667_),
    .A2(_05795_),
    .B1(_05799_),
    .B2(_05692_),
    .ZN(_05800_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21851_ (.A1(_05705_),
    .A2(_05786_),
    .ZN(_05801_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _21852_ (.A1(_05692_),
    .A2(_05786_),
    .A3(_05794_),
    .B1(_05800_),
    .B2(_05801_),
    .ZN(_05802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21853_ (.I0(\id_stage_i.controller_i.instr_i[14] ),
    .I1(_05802_),
    .S(net3069),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21854_ (.A1(_05632_),
    .A2(_05689_),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _21855_ (.I(_05632_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21856_ (.A1(_05732_),
    .A2(_05757_),
    .B(_05642_),
    .ZN(_05805_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21857_ (.A1(_05804_),
    .A2(_05689_),
    .A3(_05805_),
    .Z(_05806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21858_ (.A1(_05664_),
    .A2(_05747_),
    .B1(_05803_),
    .B2(net3395),
    .C(_05806_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21859_ (.A1(_05649_),
    .A2(_05795_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21860_ (.A1(_05692_),
    .A2(_05704_),
    .Z(_05809_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21861_ (.A1(_05804_),
    .A2(_05809_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21862_ (.A1(_05807_),
    .A2(_05808_),
    .B(_05810_),
    .C(_05786_),
    .ZN(_05811_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21863_ (.A1(_05632_),
    .A2(_05698_),
    .B(_05744_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21864_ (.A1(_05656_),
    .A2(_05660_),
    .B1(_05611_),
    .B2(_05812_),
    .ZN(_05813_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21865_ (.A1(_05689_),
    .A2(_05783_),
    .B1(_05813_),
    .B2(_05700_),
    .ZN(_05814_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21866_ (.A1(_05692_),
    .A2(_05660_),
    .Z(_05815_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _21867_ (.A1(_05656_),
    .A2(_05642_),
    .A3(_05676_),
    .Z(_05816_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21868_ (.A1(_05815_),
    .A2(_05816_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21869_ (.A1(_05804_),
    .A2(_05765_),
    .A3(_05817_),
    .Z(_05818_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21870_ (.A1(_05811_),
    .A2(_05814_),
    .A3(_05818_),
    .ZN(_05819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21871_ (.I0(net3607),
    .I1(_05819_),
    .S(net3069),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21872_ (.I0(_05258_),
    .I1(_05636_),
    .S(_08730_),
    .Z(_05820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21873_ (.A1(_05616_),
    .A2(_05816_),
    .ZN(_05821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21874_ (.A1(_05692_),
    .A2(_05821_),
    .ZN(_05822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21875_ (.I0(_05820_),
    .I1(_05822_),
    .S(_05794_),
    .Z(_05823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21876_ (.A1(_05651_),
    .A2(_05752_),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21877_ (.A1(_05642_),
    .A2(_05757_),
    .Z(_05825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21878_ (.A1(_05616_),
    .A2(_05778_),
    .B1(_05820_),
    .B2(_05825_),
    .ZN(_05826_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21879_ (.A1(_05661_),
    .A2(_05798_),
    .ZN(_05827_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21880_ (.A1(_05692_),
    .A2(_05827_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21881_ (.A1(_05645_),
    .A2(_05683_),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21882_ (.A1(_05824_),
    .A2(_05826_),
    .B(_05828_),
    .C(_05829_),
    .ZN(_05830_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21883_ (.A1(_05642_),
    .A2(_05778_),
    .B(_05757_),
    .ZN(_05831_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21884_ (.A1(_05660_),
    .A2(_05831_),
    .ZN(_05832_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21885_ (.A1(_05692_),
    .A2(_05832_),
    .B(_05656_),
    .ZN(_05833_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21886_ (.A1(_05634_),
    .A2(_05680_),
    .A3(_05732_),
    .Z(_05834_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21887_ (.A1(_05833_),
    .A2(_05830_),
    .A3(_05834_),
    .Z(_05835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21888_ (.A1(_05705_),
    .A2(_05830_),
    .B1(_05835_),
    .B2(_05616_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21889_ (.A1(_05616_),
    .A2(_05766_),
    .B1(_05767_),
    .B2(_05820_),
    .C(_05700_),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21890_ (.A1(_05700_),
    .A2(_05836_),
    .B(_05837_),
    .ZN(_05838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21891_ (.I0(_05823_),
    .I1(_05838_),
    .S(_05742_),
    .Z(_05839_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21892_ (.I0(net3605),
    .I1(_05839_),
    .S(net3069),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21893_ (.A1(_05742_),
    .A2(_05700_),
    .Z(_05840_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input48 (.I(data_rdata_i[29]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21895_ (.A1(_05628_),
    .A2(_05840_),
    .ZN(_05842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21896_ (.I0(_05360_),
    .I1(_05608_),
    .S(_08730_),
    .Z(_05843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21897_ (.A1(_05769_),
    .A2(_05843_),
    .ZN(_05844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21898_ (.A1(_05689_),
    .A2(net3395),
    .ZN(_05845_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21899_ (.A1(_05649_),
    .A2(_05752_),
    .A3(_05777_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21900_ (.A1(_05845_),
    .A2(_05846_),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21901_ (.A1(_05692_),
    .A2(_05690_),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21902_ (.A1(_05628_),
    .A2(_05831_),
    .B1(_05843_),
    .B2(_05825_),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21903_ (.A1(_05848_),
    .A2(_05849_),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21904_ (.A1(_05616_),
    .A2(_05634_),
    .Z(_05851_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21905_ (.A1(_05689_),
    .A2(_05851_),
    .A3(_05798_),
    .B(_05828_),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21906_ (.A1(_05628_),
    .A2(_05847_),
    .B(_05850_),
    .C(_05852_),
    .ZN(_05853_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _21907_ (.A1(_05760_),
    .A2(_05853_),
    .Z(_05854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21908_ (.A1(_05732_),
    .A2(_05843_),
    .ZN(_05855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21909_ (.A1(_05854_),
    .A2(_05855_),
    .B(_05809_),
    .ZN(_05856_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21910_ (.A1(_05817_),
    .A2(_05855_),
    .Z(_05857_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21911_ (.A1(_05765_),
    .A2(_05857_),
    .B(_05854_),
    .ZN(_05858_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21912_ (.A1(_05628_),
    .A2(_05856_),
    .B(_05858_),
    .ZN(_05859_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21913_ (.A1(_05766_),
    .A2(_05842_),
    .B(_05844_),
    .C(_05859_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21914_ (.I0(net3582),
    .I1(_05860_),
    .S(net3069),
    .Z(_01796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21915_ (.I0(_05431_),
    .I1(_05668_),
    .S(_08730_),
    .Z(_05861_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21916_ (.A1(_05758_),
    .A2(_05861_),
    .Z(_05862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21917_ (.A1(_05689_),
    .A2(_05680_),
    .Z(_05863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21918_ (.A1(_05752_),
    .A2(_05862_),
    .B(_05852_),
    .C(_05863_),
    .ZN(_05864_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21919_ (.A1(_05760_),
    .A2(_05864_),
    .ZN(_05865_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21920_ (.A1(_05732_),
    .A2(_05861_),
    .ZN(_05866_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21921_ (.A1(_05817_),
    .A2(_05866_),
    .B(_05765_),
    .ZN(_05867_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21922_ (.A1(_05760_),
    .A2(_05864_),
    .B(_05866_),
    .ZN(_05868_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21923_ (.A1(_05705_),
    .A2(_05868_),
    .Z(_05869_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21924_ (.A1(_05865_),
    .A2(_05867_),
    .B1(_05869_),
    .B2(_05624_),
    .ZN(_05870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21925_ (.A1(_05661_),
    .A2(_05861_),
    .B(_05698_),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21926_ (.A1(_05638_),
    .A2(_05861_),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21927_ (.A1(_05870_),
    .A2(_05872_),
    .ZN(_05873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21928_ (.A1(_05611_),
    .A2(_05873_),
    .ZN(_05874_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21929_ (.A1(_05700_),
    .A2(_05870_),
    .B1(_05871_),
    .B2(_05768_),
    .C(_05874_),
    .ZN(_05875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21930_ (.I0(net3580),
    .I1(_05875_),
    .S(net3069),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21931_ (.A1(_05661_),
    .A2(_05766_),
    .Z(_05876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21932_ (.A1(_05876_),
    .A2(_05840_),
    .B(_05783_),
    .ZN(_05877_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21933_ (.I(_05671_),
    .ZN(_05878_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21934_ (.I0(_05460_),
    .I1(_05878_),
    .S(_08730_),
    .Z(_05879_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21935_ (.A1(_05848_),
    .A2(_05758_),
    .A3(_05879_),
    .ZN(_05880_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21936_ (.A1(_05852_),
    .A2(_05880_),
    .Z(_05881_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21937_ (.A1(_05642_),
    .A2(_05676_),
    .B(_05790_),
    .ZN(_05882_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21938_ (.A1(_05660_),
    .A2(_05879_),
    .B(_05882_),
    .C(_05705_),
    .ZN(_05883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21939_ (.A1(_05786_),
    .A2(_05881_),
    .B1(_05883_),
    .B2(_05707_),
    .ZN(_05884_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21940_ (.A1(_05621_),
    .A2(_05705_),
    .ZN(_05885_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21941_ (.A1(_05877_),
    .A2(_05879_),
    .B1(_05884_),
    .B2(_05885_),
    .ZN(_05886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21942_ (.I0(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .I1(_05886_),
    .S(net3069),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21943_ (.A1(_05752_),
    .A2(_05825_),
    .Z(_05887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21944_ (.I0(_05876_),
    .I1(_05887_),
    .S(_05638_),
    .Z(_05888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21945_ (.A1(_05742_),
    .A2(_05888_),
    .ZN(_05889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21946_ (.I0(net398),
    .I1(_05889_),
    .S(net3069),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21947_ (.I0(_05479_),
    .I1(_05665_),
    .S(_08730_),
    .Z(_05890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21948_ (.A1(_05670_),
    .A2(_05698_),
    .B1(_05890_),
    .B2(_05692_),
    .ZN(_05891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21949_ (.A1(_05732_),
    .A2(_05890_),
    .ZN(_05892_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21950_ (.A1(_05656_),
    .A2(_05891_),
    .B(_05892_),
    .ZN(_05893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21951_ (.A1(_05783_),
    .A2(_05890_),
    .B1(_05893_),
    .B2(_05840_),
    .ZN(_05894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21952_ (.A1(_05656_),
    .A2(_05698_),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21953_ (.A1(_05848_),
    .A2(_05825_),
    .B(_05895_),
    .ZN(_05896_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21954_ (.A1(_05887_),
    .A2(_05890_),
    .B1(_05896_),
    .B2(_05670_),
    .C(_05852_),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21955_ (.A1(_05760_),
    .A2(_05897_),
    .ZN(_05898_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21956_ (.A1(_05635_),
    .A2(_05676_),
    .A3(_05695_),
    .Z(_05899_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21957_ (.A1(_05670_),
    .A2(_05899_),
    .B(_05682_),
    .C(_05660_),
    .ZN(_05900_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21958_ (.A1(_05892_),
    .A2(_05900_),
    .B(_05765_),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21959_ (.A1(_05670_),
    .A2(_05705_),
    .B1(_05898_),
    .B2(_05901_),
    .ZN(_05902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21960_ (.A1(_05894_),
    .A2(_05902_),
    .ZN(_05903_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input47 (.I(data_rdata_i[28]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21962_ (.I0(net3554),
    .I1(_05903_),
    .S(net3069),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21963_ (.I0(_05499_),
    .I1(_05647_),
    .S(_08730_),
    .Z(_05905_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21964_ (.A1(_05752_),
    .A2(_05757_),
    .A3(_05905_),
    .Z(_05906_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21965_ (.A1(_05795_),
    .A2(_05906_),
    .Z(_05907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21966_ (.A1(_05846_),
    .A2(_05895_),
    .ZN(_05908_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21967_ (.A1(_05642_),
    .A2(_05907_),
    .B1(_05908_),
    .B2(_05673_),
    .ZN(_05909_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21968_ (.I(_05673_),
    .ZN(_05910_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21969_ (.A1(_05796_),
    .A2(_05831_),
    .Z(_05911_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _21970_ (.A1(_05611_),
    .A2(_05794_),
    .Z(_05912_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21971_ (.A1(_05786_),
    .A2(_05911_),
    .B(_05912_),
    .ZN(_05913_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21972_ (.A1(net3395),
    .A2(_05910_),
    .A3(_05913_),
    .Z(_05914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _21973_ (.A1(_05689_),
    .A2(_05742_),
    .ZN(_05915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21974_ (.A1(_05673_),
    .A2(_05698_),
    .B1(_05905_),
    .B2(_05692_),
    .ZN(_05916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21975_ (.A1(_05732_),
    .A2(_05905_),
    .ZN(_05917_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21976_ (.A1(_05915_),
    .A2(_05916_),
    .B(_05917_),
    .ZN(_05918_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21977_ (.A1(_05673_),
    .A2(_05660_),
    .A3(_05707_),
    .A4(_05863_),
    .Z(_05919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21978_ (.A1(_05783_),
    .A2(_05905_),
    .B1(_05918_),
    .B2(_05700_),
    .C(_05919_),
    .ZN(_05920_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21979_ (.A1(_05801_),
    .A2(_05909_),
    .B(_05914_),
    .C(_05920_),
    .ZN(_05921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21980_ (.I0(net3552),
    .I1(_05921_),
    .S(net3069),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21981_ (.I0(_05511_),
    .I1(_05643_),
    .S(_08730_),
    .Z(_05922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _21982_ (.A1(_05642_),
    .A2(_05795_),
    .B1(_05887_),
    .B2(_05922_),
    .C1(_05896_),
    .C2(_05667_),
    .ZN(_05923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21983_ (.A1(_05796_),
    .A2(_05786_),
    .B(_05912_),
    .ZN(_05924_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21984_ (.A1(_05765_),
    .A2(_05661_),
    .B1(_05924_),
    .B2(net3395),
    .ZN(_05925_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21985_ (.A1(_05689_),
    .A2(_05698_),
    .A3(_05840_),
    .Z(_05926_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21986_ (.A1(_05925_),
    .A2(_05926_),
    .B(_05667_),
    .ZN(_05927_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21987_ (.A1(_05667_),
    .A2(_05863_),
    .Z(_05928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21988_ (.I0(_05922_),
    .I1(_05928_),
    .S(_05660_),
    .Z(_05929_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21989_ (.A1(_05645_),
    .A2(_05704_),
    .A3(_05840_),
    .Z(_05930_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21990_ (.A1(_05769_),
    .A2(_05922_),
    .B1(_05929_),
    .B2(_05707_),
    .C(_05930_),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21991_ (.A1(_05801_),
    .A2(_05923_),
    .B(_05927_),
    .C(_05931_),
    .ZN(_05932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21992_ (.I0(net3499),
    .I1(_05932_),
    .S(net3069),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21993_ (.A1(_05642_),
    .A2(_05795_),
    .ZN(_05933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21994_ (.I0(_05520_),
    .I1(_05630_),
    .S(_08730_),
    .Z(_05934_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21995_ (.A1(_05664_),
    .A2(_05934_),
    .Z(_05935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21996_ (.I0(_05649_),
    .I1(_05935_),
    .S(_05757_),
    .Z(_05936_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21997_ (.A1(_05656_),
    .A2(net3395),
    .A3(_05649_),
    .Z(_05937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21998_ (.A1(_05744_),
    .A2(_05936_),
    .B(_05937_),
    .ZN(_05938_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21999_ (.A1(_05732_),
    .A2(_05938_),
    .Z(_05939_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22000_ (.A1(_05933_),
    .A2(_05939_),
    .Z(_05940_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22001_ (.A1(_05624_),
    .A2(_05895_),
    .B1(_05934_),
    .B2(_05767_),
    .C(_05840_),
    .ZN(_05941_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22002_ (.I(_05941_),
    .ZN(_05942_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22003_ (.A1(_05925_),
    .A2(_05942_),
    .B(_05649_),
    .ZN(_05943_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22004_ (.A1(_05649_),
    .A2(_05863_),
    .Z(_05944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22005_ (.I0(_05934_),
    .I1(_05944_),
    .S(_05794_),
    .Z(_05945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22006_ (.A1(_05611_),
    .A2(_05945_),
    .B1(_05942_),
    .B2(_05705_),
    .ZN(_05946_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22007_ (.A1(_05801_),
    .A2(_05940_),
    .B(_05943_),
    .C(_05946_),
    .ZN(_05947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22008_ (.I0(net3498),
    .I1(_05947_),
    .S(net3069),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22009_ (.I0(_05529_),
    .I1(_05614_),
    .S(_08730_),
    .Z(_05948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22010_ (.A1(_05660_),
    .A2(_05700_),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22011_ (.I0(_05645_),
    .I1(_05948_),
    .S(_05949_),
    .Z(_05950_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22012_ (.I(_05950_),
    .ZN(_05951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22013_ (.A1(_05621_),
    .A2(_05704_),
    .B1(_05876_),
    .B2(_05948_),
    .C(_05768_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22014_ (.A1(_05642_),
    .A2(_05948_),
    .Z(_05953_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22015_ (.I0(_05645_),
    .I1(_05953_),
    .S(_05757_),
    .Z(_05954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22016_ (.A1(_05621_),
    .A2(_05747_),
    .B1(_05752_),
    .B2(_05954_),
    .C(_05760_),
    .ZN(_05955_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _22017_ (.I(_05645_),
    .ZN(_05956_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22018_ (.A1(net3395),
    .A2(_05851_),
    .B(_05660_),
    .ZN(_05957_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22019_ (.A1(_05689_),
    .A2(_05956_),
    .A3(_05957_),
    .Z(_05958_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22020_ (.A1(_05933_),
    .A2(_05955_),
    .A3(_05958_),
    .Z(_05959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22021_ (.A1(_05611_),
    .A2(_05951_),
    .B(_05952_),
    .C(_05959_),
    .ZN(_05960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22022_ (.I0(net3487),
    .I1(_05960_),
    .S(net3069),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22023_ (.I(_05626_),
    .ZN(_05961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22024_ (.I0(_05538_),
    .I1(_05961_),
    .S(_08730_),
    .Z(_05962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22025_ (.I0(_05664_),
    .I1(_05962_),
    .S(_05876_),
    .Z(_05963_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22026_ (.A1(_05664_),
    .A2(_05766_),
    .B(_05611_),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22027_ (.A1(_05611_),
    .A2(_05949_),
    .Z(_05965_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22028_ (.I(_05962_),
    .ZN(_05966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22029_ (.A1(_05700_),
    .A2(_05964_),
    .B1(_05965_),
    .B2(_05966_),
    .ZN(_05967_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22030_ (.A1(_05704_),
    .A2(_05795_),
    .B(_05642_),
    .ZN(_05968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22031_ (.A1(_05705_),
    .A2(_05968_),
    .ZN(_05969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22032_ (.A1(_05624_),
    .A2(_05962_),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22033_ (.A1(_05642_),
    .A2(_05790_),
    .A3(_05970_),
    .Z(_05971_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22034_ (.A1(_05692_),
    .A2(_05851_),
    .B(_05732_),
    .ZN(_05972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22035_ (.A1(_05845_),
    .A2(_05972_),
    .ZN(_05973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22036_ (.A1(_05670_),
    .A2(_05973_),
    .Z(_05974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22037_ (.A1(_05664_),
    .A2(_05809_),
    .B(_05760_),
    .ZN(_05975_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _22038_ (.A1(_05969_),
    .A2(_05971_),
    .A3(_05974_),
    .B(_05975_),
    .ZN(_05976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22039_ (.A1(_05840_),
    .A2(_05963_),
    .B1(_05967_),
    .B2(_05976_),
    .ZN(_05977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22040_ (.I0(\id_stage_i.controller_i.instr_i[25] ),
    .I1(_05977_),
    .S(net3069),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22041_ (.A1(_05656_),
    .A2(_05698_),
    .B(_05795_),
    .ZN(_05978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22042_ (.I0(_05273_),
    .I1(_05622_),
    .S(_08730_),
    .Z(_05979_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22043_ (.A1(_05687_),
    .A2(_05979_),
    .B(_05790_),
    .ZN(_05980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22044_ (.A1(_05978_),
    .A2(_05980_),
    .ZN(_05981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22045_ (.A1(_05642_),
    .A2(_05981_),
    .ZN(_05982_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22046_ (.A1(_05649_),
    .A2(_05851_),
    .Z(_05983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22047_ (.I0(_05632_),
    .I1(_05983_),
    .S(net3395),
    .Z(_05984_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22048_ (.A1(_05732_),
    .A2(_05984_),
    .B(_05944_),
    .C(_05809_),
    .ZN(_05985_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22049_ (.A1(_05642_),
    .A2(_05705_),
    .B(_05786_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22050_ (.A1(_05982_),
    .A2(_05985_),
    .B(_05986_),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22051_ (.A1(_05656_),
    .A2(_05670_),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22052_ (.A1(_05803_),
    .A2(_05988_),
    .B(_05765_),
    .C(_05766_),
    .ZN(_05989_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22053_ (.I(_05979_),
    .ZN(_05990_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22054_ (.A1(_05649_),
    .A2(_05766_),
    .B(_05840_),
    .C(_05810_),
    .ZN(_05991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22055_ (.A1(_05965_),
    .A2(_05979_),
    .ZN(_05992_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22056_ (.A1(_05876_),
    .A2(_05990_),
    .B1(_05991_),
    .B2(_05992_),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _22057_ (.A1(_05987_),
    .A2(_05989_),
    .A3(_05993_),
    .Z(_05994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22058_ (.I0(net3485),
    .I1(_05994_),
    .S(net3069),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22059_ (.I0(_05281_),
    .I1(_05618_),
    .S(_08730_),
    .Z(_05995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22060_ (.A1(_05616_),
    .A2(_05809_),
    .B1(_05876_),
    .B2(_05995_),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22061_ (.A1(_05687_),
    .A2(_05995_),
    .B(_05790_),
    .ZN(_05997_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22062_ (.A1(_05978_),
    .A2(_05997_),
    .Z(_05998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22063_ (.A1(_05645_),
    .A2(_05732_),
    .B(_05704_),
    .C(net3395),
    .ZN(_05999_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22064_ (.A1(_05656_),
    .A2(_05673_),
    .Z(_06000_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22065_ (.A1(_05732_),
    .A2(_05851_),
    .A3(_06000_),
    .Z(_06001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22066_ (.A1(_05689_),
    .A2(_05645_),
    .B(_06001_),
    .C(_05692_),
    .ZN(_06002_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _22067_ (.A1(_05664_),
    .A2(_05998_),
    .B1(_05999_),
    .B2(_06002_),
    .ZN(_06003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22068_ (.A1(_05616_),
    .A2(_05689_),
    .B(_06000_),
    .ZN(_06004_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22069_ (.A1(_05766_),
    .A2(_06004_),
    .B(_05611_),
    .ZN(_06005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22070_ (.A1(_05965_),
    .A2(_05995_),
    .B1(_06003_),
    .B2(_05975_),
    .C1(_06005_),
    .C2(_05700_),
    .ZN(_06006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22071_ (.A1(_05840_),
    .A2(_05996_),
    .B(_06006_),
    .ZN(_06007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22072_ (.I0(\id_stage_i.controller_i.instr_i[27] ),
    .I1(_06007_),
    .S(net3069),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22073_ (.A1(_05656_),
    .A2(_05667_),
    .A3(_05851_),
    .Z(_06008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22074_ (.I0(_05628_),
    .I1(_06008_),
    .S(net3395),
    .Z(_06009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22075_ (.I0(_05290_),
    .I1(_05640_),
    .S(_08730_),
    .Z(_06010_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22076_ (.A1(_05687_),
    .A2(_06010_),
    .B(_05790_),
    .ZN(_06011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22077_ (.A1(_05845_),
    .A2(_06011_),
    .B(_05664_),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22078_ (.A1(_05732_),
    .A2(_06009_),
    .B(_06012_),
    .C(_05969_),
    .ZN(_06013_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _22079_ (.I(_05770_),
    .ZN(_06014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22080_ (.A1(_06014_),
    .A2(_06010_),
    .ZN(_06015_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22081_ (.A1(_05705_),
    .A2(_05842_),
    .B1(_05986_),
    .B2(_06013_),
    .C(_06015_),
    .ZN(_06016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22082_ (.I0(net3483),
    .I1(_06016_),
    .S(net3069),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22083_ (.I0(_05298_),
    .I1(_05657_),
    .S(_08730_),
    .Z(_06017_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22084_ (.A1(_05687_),
    .A2(_06017_),
    .B(_05790_),
    .ZN(_06018_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22085_ (.A1(_05692_),
    .A2(_05661_),
    .A3(_06018_),
    .ZN(_06019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22086_ (.A1(_05624_),
    .A2(_05747_),
    .B1(_06019_),
    .B2(_05642_),
    .ZN(_06020_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22087_ (.A1(_05624_),
    .A2(_05809_),
    .A3(_05840_),
    .Z(_06021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22088_ (.A1(_06014_),
    .A2(_06017_),
    .B(_06021_),
    .ZN(_06022_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22089_ (.A1(_05760_),
    .A2(_06020_),
    .B(_06022_),
    .ZN(_06023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22090_ (.I0(net3482),
    .I1(_06023_),
    .S(net3069),
    .Z(_01809_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22091_ (.A1(_05747_),
    .A2(_05795_),
    .ZN(_06024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22092_ (.A1(_05635_),
    .A2(_05642_),
    .ZN(_06025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22093_ (.A1(_05670_),
    .A2(_05732_),
    .B1(_05753_),
    .B2(_06025_),
    .ZN(_06026_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22094_ (.A1(_05765_),
    .A2(_05809_),
    .A3(_06026_),
    .Z(_06027_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _22095_ (.A1(_05848_),
    .A2(_05758_),
    .A3(_05801_),
    .Z(_06028_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22096_ (.A1(_05877_),
    .A2(_06028_),
    .ZN(_06029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22097_ (.A1(_05670_),
    .A2(_06029_),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22098_ (.A1(_05801_),
    .A2(_06024_),
    .B(_06027_),
    .C(_06030_),
    .ZN(_06031_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input46 (.I(data_rdata_i[27]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22100_ (.I0(net3481),
    .I1(_06031_),
    .S(net3069),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22101_ (.I0(_05306_),
    .I1(_05678_),
    .S(_08730_),
    .Z(_06033_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22102_ (.A1(_05621_),
    .A2(_05650_),
    .B(_05687_),
    .ZN(_06034_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22103_ (.A1(_05642_),
    .A2(_06034_),
    .B1(_06033_),
    .B2(_05758_),
    .C(_05625_),
    .ZN(_06035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22104_ (.A1(_05617_),
    .A2(_05732_),
    .B1(_05690_),
    .B2(_06035_),
    .ZN(_06036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22105_ (.I0(_05642_),
    .I1(_06036_),
    .S(_05692_),
    .Z(_06037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22106_ (.A1(_06014_),
    .A2(_06033_),
    .B1(_06037_),
    .B2(_05975_),
    .C(_05112_),
    .ZN(_06038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22107_ (.A1(_06762_),
    .A2(_05112_),
    .B(_06038_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22108_ (.I0(_05314_),
    .I1(_05653_),
    .S(_08730_),
    .Z(_06039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22109_ (.I(_06039_),
    .ZN(_06040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22110_ (.A1(_05624_),
    .A2(_06040_),
    .ZN(_06041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22111_ (.A1(_05621_),
    .A2(_06041_),
    .B(_05848_),
    .ZN(_06042_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _22112_ (.A1(_05664_),
    .A2(_05760_),
    .A3(_06042_),
    .B1(_06040_),
    .B2(_05770_),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22113_ (.I0(net3479),
    .I1(_06043_),
    .S(net3069),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22114_ (.A1(_05770_),
    .A2(_06028_),
    .Z(_06044_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _22115_ (.A1(_05775_),
    .A2(_05801_),
    .B1(_06044_),
    .B2(_05910_),
    .ZN(_06045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22116_ (.I0(net3478),
    .I1(_06045_),
    .S(net3069),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22117_ (.A1(_05660_),
    .A2(_05915_),
    .B(_05667_),
    .ZN(_06046_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _22118_ (.A1(_05676_),
    .A2(_05611_),
    .A3(_05690_),
    .A4(_06025_),
    .Z(_06047_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _22119_ (.A1(_05638_),
    .A2(_05698_),
    .A3(_06046_),
    .A4(_06047_),
    .Z(_06048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22120_ (.A1(_05689_),
    .A2(_05825_),
    .B(_05611_),
    .ZN(_06049_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22121_ (.A1(_05775_),
    .A2(_05845_),
    .Z(_06050_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22122_ (.A1(_05667_),
    .A2(_06049_),
    .B1(_06050_),
    .B2(_05611_),
    .C(_05638_),
    .ZN(_06051_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22123_ (.A1(_06048_),
    .A2(_06051_),
    .ZN(_06052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22124_ (.I0(\id_stage_i.controller_i.instr_i[4] ),
    .I1(_06052_),
    .S(net3069),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22125_ (.A1(net3395),
    .A2(_05649_),
    .B(_05700_),
    .ZN(_06053_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22126_ (.A1(_05742_),
    .A2(_06053_),
    .ZN(_06054_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22127_ (.A1(_05638_),
    .A2(_05661_),
    .B1(_05794_),
    .B2(_05649_),
    .C(_06054_),
    .ZN(_06055_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22128_ (.A1(_05664_),
    .A2(_05649_),
    .B(_05757_),
    .ZN(_06056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22129_ (.A1(_05692_),
    .A2(_06056_),
    .B(_05656_),
    .ZN(_06057_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22130_ (.A1(_05682_),
    .A2(_05772_),
    .B1(_06057_),
    .B2(_05732_),
    .C(_05786_),
    .ZN(_06058_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22131_ (.A1(_06055_),
    .A2(_06058_),
    .ZN(_06059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22132_ (.I0(\id_stage_i.controller_i.instr_i[5] ),
    .I1(_06059_),
    .S(net3069),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22133_ (.A1(_05676_),
    .A2(_05744_),
    .A3(_05912_),
    .ZN(_06060_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22134_ (.A1(_05956_),
    .A2(_06044_),
    .B1(_06050_),
    .B2(_05760_),
    .C(_06060_),
    .ZN(_06061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22135_ (.I0(net354),
    .I1(_06061_),
    .S(net3069),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22136_ (.I(_05676_),
    .ZN(_06062_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _22137_ (.A1(_05635_),
    .A2(_05664_),
    .A3(_06062_),
    .B(_05689_),
    .ZN(_06063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22138_ (.A1(_05632_),
    .A2(_06062_),
    .B1(_05660_),
    .B2(_06063_),
    .ZN(_06064_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22139_ (.A1(_05804_),
    .A2(_05690_),
    .B1(_06064_),
    .B2(net3395),
    .C(_05700_),
    .ZN(_06065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22140_ (.A1(_05810_),
    .A2(_06065_),
    .ZN(_06066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22141_ (.A1(_05670_),
    .A2(_05704_),
    .B1(_05876_),
    .B2(_05632_),
    .C(_05768_),
    .ZN(_06067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22142_ (.I0(_05804_),
    .I1(_05689_),
    .S(_05732_),
    .Z(_06068_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _22143_ (.A1(_05664_),
    .A2(_05845_),
    .B1(_06068_),
    .B2(net3395),
    .ZN(_06069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22144_ (.A1(_05632_),
    .A2(_05915_),
    .B1(_06069_),
    .B2(_05742_),
    .C(_05700_),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22145_ (.A1(_05611_),
    .A2(_06066_),
    .B(_06067_),
    .C(_06070_),
    .ZN(_06071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22146_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .I1(_06071_),
    .S(net3069),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22147_ (.A1(net3395),
    .A2(_05676_),
    .B(_05690_),
    .ZN(_06072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22148_ (.A1(_05616_),
    .A2(_06072_),
    .ZN(_06073_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _22149_ (.A1(_05617_),
    .A2(_05689_),
    .B1(_05910_),
    .B2(_05915_),
    .ZN(_06074_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22150_ (.A1(_05611_),
    .A2(_05815_),
    .Z(_06075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22151_ (.A1(net3395),
    .A2(_06074_),
    .B1(_06075_),
    .B2(_05616_),
    .C(_05700_),
    .ZN(_06076_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22152_ (.A1(_05673_),
    .A2(_05704_),
    .B1(_05876_),
    .B2(_05616_),
    .C(_05768_),
    .ZN(_06077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22153_ (.A1(_05707_),
    .A2(_06073_),
    .B(_06076_),
    .C(_06077_),
    .ZN(_06078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22154_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .I1(_06078_),
    .S(net3069),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22155_ (.A1(net3395),
    .A2(_05742_),
    .ZN(_06079_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22156_ (.A1(net3395),
    .A2(_05675_),
    .A3(_05949_),
    .Z(_06080_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22157_ (.A1(_06079_),
    .A2(_06080_),
    .B(_05656_),
    .C(_05667_),
    .ZN(_06081_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22158_ (.A1(_05700_),
    .A2(_05747_),
    .B(_05742_),
    .ZN(_06082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22159_ (.A1(_05786_),
    .A2(_05863_),
    .B1(_06082_),
    .B2(_05628_),
    .ZN(_06083_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22160_ (.A1(net3395),
    .A2(_05956_),
    .ZN(_06084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22161_ (.I0(_05667_),
    .I1(_06084_),
    .S(_05689_),
    .Z(_06085_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22162_ (.A1(_05628_),
    .A2(_05767_),
    .B1(_06085_),
    .B2(_05732_),
    .C(_05840_),
    .ZN(_06086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22163_ (.A1(_06081_),
    .A2(_06083_),
    .B(_06086_),
    .ZN(_06087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22164_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .I1(_06087_),
    .S(net3069),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22165_ (.I0(\cs_registers_i.pc_id_i[10] ),
    .I1(\cs_registers_i.pc_if_i[10] ),
    .S(net3070),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input45 (.I(data_rdata_i[26]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22167_ (.I0(\cs_registers_i.pc_id_i[11] ),
    .I1(\cs_registers_i.pc_if_i[11] ),
    .S(net3070),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22168_ (.I0(\cs_registers_i.pc_id_i[12] ),
    .I1(\cs_registers_i.pc_if_i[12] ),
    .S(net3070),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22169_ (.I0(\cs_registers_i.pc_id_i[13] ),
    .I1(\cs_registers_i.pc_if_i[13] ),
    .S(net3070),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22170_ (.I0(\cs_registers_i.pc_id_i[14] ),
    .I1(\cs_registers_i.pc_if_i[14] ),
    .S(net3070),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22171_ (.I0(\cs_registers_i.pc_id_i[15] ),
    .I1(\cs_registers_i.pc_if_i[15] ),
    .S(net3070),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22172_ (.I0(\cs_registers_i.pc_id_i[16] ),
    .I1(\cs_registers_i.pc_if_i[16] ),
    .S(net3070),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22173_ (.I0(\cs_registers_i.pc_id_i[17] ),
    .I1(\cs_registers_i.pc_if_i[17] ),
    .S(net3070),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22174_ (.I0(\cs_registers_i.pc_id_i[18] ),
    .I1(\cs_registers_i.pc_if_i[18] ),
    .S(net3070),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22175_ (.I0(\cs_registers_i.pc_id_i[19] ),
    .I1(\cs_registers_i.pc_if_i[19] ),
    .S(net3070),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22176_ (.I0(\cs_registers_i.pc_id_i[1] ),
    .I1(net3653),
    .S(net3070),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input44 (.I(data_rdata_i[25]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22178_ (.I0(\cs_registers_i.pc_id_i[20] ),
    .I1(\cs_registers_i.pc_if_i[20] ),
    .S(net3070),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22179_ (.I0(\cs_registers_i.pc_id_i[21] ),
    .I1(\cs_registers_i.pc_if_i[21] ),
    .S(net3070),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22180_ (.I0(\cs_registers_i.pc_id_i[22] ),
    .I1(\cs_registers_i.pc_if_i[22] ),
    .S(net3070),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22181_ (.I0(\cs_registers_i.pc_id_i[23] ),
    .I1(\cs_registers_i.pc_if_i[23] ),
    .S(net3070),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22182_ (.I0(\cs_registers_i.pc_id_i[24] ),
    .I1(\cs_registers_i.pc_if_i[24] ),
    .S(net3070),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22183_ (.I0(\cs_registers_i.pc_id_i[25] ),
    .I1(\cs_registers_i.pc_if_i[25] ),
    .S(net3070),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22184_ (.I0(\cs_registers_i.pc_id_i[26] ),
    .I1(\cs_registers_i.pc_if_i[26] ),
    .S(net3070),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22185_ (.I0(\cs_registers_i.pc_id_i[27] ),
    .I1(\cs_registers_i.pc_if_i[27] ),
    .S(net3070),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22186_ (.I0(\cs_registers_i.pc_id_i[28] ),
    .I1(\cs_registers_i.pc_if_i[28] ),
    .S(net3070),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22187_ (.I0(\cs_registers_i.pc_id_i[29] ),
    .I1(\cs_registers_i.pc_if_i[29] ),
    .S(net3070),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input43 (.I(data_rdata_i[24]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22189_ (.I0(\cs_registers_i.pc_id_i[2] ),
    .I1(\cs_registers_i.pc_if_i[2] ),
    .S(net3070),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22190_ (.I0(\cs_registers_i.pc_id_i[30] ),
    .I1(\cs_registers_i.pc_if_i[30] ),
    .S(net3070),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22191_ (.I0(\cs_registers_i.pc_id_i[31] ),
    .I1(\cs_registers_i.pc_if_i[31] ),
    .S(net3070),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22192_ (.I0(\cs_registers_i.pc_id_i[3] ),
    .I1(\cs_registers_i.pc_if_i[3] ),
    .S(net3070),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22193_ (.I0(\cs_registers_i.pc_id_i[4] ),
    .I1(\cs_registers_i.pc_if_i[4] ),
    .S(net3070),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22194_ (.I0(\cs_registers_i.pc_id_i[5] ),
    .I1(\cs_registers_i.pc_if_i[5] ),
    .S(net3070),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22195_ (.I0(\cs_registers_i.pc_id_i[6] ),
    .I1(\cs_registers_i.pc_if_i[6] ),
    .S(net3070),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22196_ (.I0(\cs_registers_i.pc_id_i[7] ),
    .I1(\cs_registers_i.pc_if_i[7] ),
    .S(net3070),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22197_ (.I0(\cs_registers_i.pc_id_i[8] ),
    .I1(\cs_registers_i.pc_if_i[8] ),
    .S(net3070),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22198_ (.I0(\cs_registers_i.pc_id_i[9] ),
    .I1(\cs_registers_i.pc_if_i[9] ),
    .S(net3070),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _22199_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_08877_),
    .Z(net249));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _22200_ (.A1(net3472),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A4(_05570_),
    .Z(_06091_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22201_ (.A1(_04367_),
    .A2(net249),
    .A3(_06091_),
    .Z(core_busy_d));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22202_ (.A1(clknet_1_0__leaf_clk_i),
    .A2(net641),
    .Z(clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22203_ (.I(_11643_[0]),
    .ZN(_06092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22204_ (.I0(_11658_[0]),
    .I1(_06092_),
    .S(net320),
    .Z(_06093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22205_ (.I0(_06093_),
    .I1(_11644_[0]),
    .S(_05573_),
    .Z(net181));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input42 (.I(data_rdata_i[23]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input41 (.I(data_rdata_i[22]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22208_ (.A1(_11651_[0]),
    .A2(_11647_[0]),
    .B(_05573_),
    .ZN(_06096_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input40 (.I(data_rdata_i[21]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _22210_ (.A1(_11658_[0]),
    .A2(_11656_[0]),
    .A3(\load_store_unit_i.handle_misaligned_q ),
    .ZN(_06098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22211_ (.A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_06096_),
    .B(_06098_),
    .ZN(_06099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22212_ (.I0(_06099_),
    .I1(_11654_[0]),
    .S(_08888_),
    .Z(net182));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22213_ (.A1(net320),
    .A2(_11646_[0]),
    .ZN(_06100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22214_ (.I0(_06100_),
    .I1(_11645_[0]),
    .S(_05573_),
    .Z(_06101_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22215_ (.A1(_11647_[0]),
    .A2(\load_store_unit_i.handle_misaligned_q ),
    .A3(_05573_),
    .Z(_06102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22216_ (.A1(_11649_[0]),
    .A2(_08888_),
    .B(_06102_),
    .ZN(_06103_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22217_ (.A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_06101_),
    .B(_06103_),
    .ZN(net183));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22218_ (.A1(net320),
    .A2(_05573_),
    .Z(_06104_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22219_ (.A1(net320),
    .A2(_11651_[0]),
    .B(_11647_[0]),
    .C(_05573_),
    .ZN(_06105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22220_ (.A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_06104_),
    .B(_06105_),
    .ZN(net184));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22221_ (.A1(_05570_),
    .A2(_08883_),
    .Z(_06106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22222_ (.A1(_06232_),
    .A2(_06106_),
    .Z(net185));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input39 (.I(data_rdata_i[20]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22224_ (.A1(_11647_[0]),
    .A2(net413),
    .B1(_07544_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07936_),
    .ZN(_06108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22225_ (.I(_06108_),
    .ZN(_06109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22226_ (.I0(_06384_),
    .I1(_06109_),
    .S(_08425_),
    .Z(net186));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input38 (.I(data_rdata_i[1]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input37 (.I(data_rdata_i[19]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22229_ (.A1(_11656_[0]),
    .A2(net557),
    .B1(_07641_),
    .B2(_11647_[0]),
    .C1(_08017_),
    .C2(_11651_[0]),
    .ZN(_06112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22230_ (.I(_06112_),
    .ZN(_06113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22231_ (.I0(_06805_),
    .I1(_06113_),
    .S(_08425_),
    .Z(net187));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input36 (.I(data_rdata_i[18]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22233_ (.A1(_11656_[0]),
    .A2(_06487_),
    .B1(_07676_),
    .B2(_11647_[0]),
    .C1(_08055_),
    .C2(_11651_[0]),
    .ZN(_06115_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22234_ (.I(_06115_),
    .ZN(_06116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22235_ (.I0(_08543_),
    .I1(_06116_),
    .S(_08425_),
    .Z(net188));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22236_ (.A1(_11656_[0]),
    .A2(net330),
    .B1(_07732_),
    .B2(_11647_[0]),
    .C1(net530),
    .C2(_11651_[0]),
    .ZN(_06117_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22237_ (.I(_06117_),
    .ZN(_06118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22238_ (.I0(net420),
    .I1(_06118_),
    .S(_08425_),
    .Z(net189));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22239_ (.A1(_11656_[0]),
    .A2(net342),
    .B1(net442),
    .B2(_11647_[0]),
    .C1(_08145_),
    .C2(_11651_[0]),
    .ZN(_06119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22240_ (.I(_06119_),
    .ZN(_06120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22241_ (.I0(net424),
    .I1(_06120_),
    .S(_08425_),
    .Z(net190));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22242_ (.A1(_11656_[0]),
    .A2(net429),
    .B1(_07838_),
    .B2(_11647_[0]),
    .C1(_08193_),
    .C2(_11651_[0]),
    .ZN(_06121_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22243_ (.I(_06121_),
    .ZN(_06122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22244_ (.I0(_07449_),
    .I1(_06122_),
    .S(_08425_),
    .Z(net191));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22245_ (.A1(_11656_[0]),
    .A2(net427),
    .B1(_07875_),
    .B2(_11647_[0]),
    .C1(_08231_),
    .C2(_11651_[0]),
    .ZN(_06123_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22246_ (.I(_06123_),
    .ZN(_06124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22247_ (.I0(_07486_),
    .I1(_06124_),
    .S(_08425_),
    .Z(net192));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input35 (.I(data_rdata_i[17]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22249_ (.A1(_11651_[0]),
    .A2(_06384_),
    .B1(_07936_),
    .B2(_11647_[0]),
    .C1(net413),
    .C2(_11656_[0]),
    .ZN(_06126_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22250_ (.I(_06126_),
    .ZN(_06127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22251_ (.I0(_07544_),
    .I1(_06127_),
    .S(_08425_),
    .Z(net193));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22252_ (.A1(_11651_[0]),
    .A2(net468),
    .B1(_07973_),
    .B2(_11647_[0]),
    .C1(net407),
    .C2(_11656_[0]),
    .ZN(_06128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22253_ (.I(_06128_),
    .ZN(_06129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22254_ (.I0(_07582_),
    .I1(_06129_),
    .S(_08425_),
    .Z(net194));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22255_ (.A1(_11651_[0]),
    .A2(_06457_),
    .B1(_08017_),
    .B2(_11647_[0]),
    .C1(_06805_),
    .C2(_11656_[0]),
    .ZN(_06130_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22256_ (.I(_06130_),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input34 (.I(data_rdata_i[16]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22258_ (.I0(_07641_),
    .I1(_06131_),
    .S(_08425_),
    .Z(net195));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22259_ (.A1(_11651_[0]),
    .A2(net436),
    .B1(_08055_),
    .B2(_11647_[0]),
    .C1(net421),
    .C2(_11656_[0]),
    .ZN(_06133_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22260_ (.I(_06133_),
    .ZN(_06134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22261_ (.I0(_07676_),
    .I1(_06134_),
    .S(_08425_),
    .Z(net196));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input33 (.I(data_rdata_i[15]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22263_ (.A1(_11647_[0]),
    .A2(net407),
    .B1(_07582_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07973_),
    .ZN(_06136_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22264_ (.I(_06136_),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22265_ (.I0(net468),
    .I1(_06137_),
    .S(_08425_),
    .Z(net197));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22266_ (.A1(_11651_[0]),
    .A2(net330),
    .B1(net530),
    .B2(_11647_[0]),
    .C1(net420),
    .C2(_11656_[0]),
    .ZN(_06138_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22267_ (.I(_06138_),
    .ZN(_06139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22268_ (.I0(_07732_),
    .I1(_06139_),
    .S(_08425_),
    .Z(net198));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22269_ (.A1(_11651_[0]),
    .A2(net342),
    .B1(_08145_),
    .B2(_11647_[0]),
    .C1(net424),
    .C2(_11656_[0]),
    .ZN(_06140_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22270_ (.I(_06140_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22271_ (.I0(_07776_),
    .I1(_06141_),
    .S(_08425_),
    .Z(net199));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22272_ (.A1(_11651_[0]),
    .A2(net429),
    .B1(_08193_),
    .B2(_11647_[0]),
    .C1(_07449_),
    .C2(_11656_[0]),
    .ZN(_06142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22273_ (.I(_06142_),
    .ZN(_06143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22274_ (.I0(_07838_),
    .I1(_06143_),
    .S(_08425_),
    .Z(net200));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22275_ (.A1(_11651_[0]),
    .A2(net427),
    .B1(net430),
    .B2(_11647_[0]),
    .C1(_07486_),
    .C2(_11656_[0]),
    .ZN(_06144_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22276_ (.I(_06144_),
    .ZN(_06145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22277_ (.I0(_07875_),
    .I1(_06145_),
    .S(_08425_),
    .Z(net201));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22278_ (.A1(_11647_[0]),
    .A2(_06384_),
    .B1(net413),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07544_),
    .ZN(_06146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22279_ (.I(_06146_),
    .ZN(_06147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22280_ (.I0(_07936_),
    .I1(_06147_),
    .S(_08425_),
    .Z(net202));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22281_ (.A1(_11647_[0]),
    .A2(net468),
    .B1(net407),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07582_),
    .ZN(_06148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22282_ (.I(_06148_),
    .ZN(_06149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22283_ (.I0(_07973_),
    .I1(_06149_),
    .S(_08425_),
    .Z(net203));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22284_ (.A1(_11647_[0]),
    .A2(_06457_),
    .B1(_06805_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07641_),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22285_ (.I(_06150_),
    .ZN(_06151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22286_ (.I0(_08017_),
    .I1(_06151_),
    .S(_08425_),
    .Z(net204));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22287_ (.A1(_11647_[0]),
    .A2(_06487_),
    .B1(_08543_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07676_),
    .ZN(_06152_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22288_ (.I(_06152_),
    .ZN(_06153_));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input32 (.I(data_rdata_i[14]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22290_ (.I0(_08055_),
    .I1(_06153_),
    .S(_08425_),
    .Z(net205));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22291_ (.A1(_11647_[0]),
    .A2(net330),
    .B1(net420),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(net410),
    .ZN(_06155_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22292_ (.I(_06155_),
    .ZN(_06156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22293_ (.I0(net530),
    .I1(_06156_),
    .S(_08425_),
    .Z(net206));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22294_ (.A1(_11647_[0]),
    .A2(net342),
    .B1(net424),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07776_),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22295_ (.I(_06157_),
    .ZN(_06158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22296_ (.I0(_08145_),
    .I1(_06158_),
    .S(_08425_),
    .Z(net207));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22297_ (.A1(_11647_[0]),
    .A2(_06805_),
    .B1(net438),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_08017_),
    .ZN(_06159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22298_ (.I(_06159_),
    .ZN(_06160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22299_ (.I0(_06457_),
    .I1(_06160_),
    .S(_08425_),
    .Z(net208));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22300_ (.A1(_11647_[0]),
    .A2(net429),
    .B1(_07449_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07838_),
    .ZN(_06161_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22301_ (.I(_06161_),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22302_ (.I0(_08193_),
    .I1(_06162_),
    .S(_08425_),
    .Z(net209));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22303_ (.A1(_11647_[0]),
    .A2(net427),
    .B1(_07486_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_07875_),
    .ZN(_06163_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22304_ (.I(_06163_),
    .ZN(_06164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22305_ (.I0(_08231_),
    .I1(_06164_),
    .S(_08425_),
    .Z(net210));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22306_ (.A1(_11647_[0]),
    .A2(_08543_),
    .B1(_07676_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_08055_),
    .ZN(_06165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22307_ (.I(_06165_),
    .ZN(_06166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22308_ (.I0(_06487_),
    .I1(_06166_),
    .S(_08425_),
    .Z(net211));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22309_ (.A1(_11647_[0]),
    .A2(net420),
    .B1(_07732_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(net530),
    .ZN(_06167_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22310_ (.I(_06167_),
    .ZN(_06168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22311_ (.I0(net330),
    .I1(_06168_),
    .S(_08425_),
    .Z(net212));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22312_ (.A1(_11647_[0]),
    .A2(net424),
    .B1(net442),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_08145_),
    .ZN(_06169_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22313_ (.I(_06169_),
    .ZN(_06170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22314_ (.I0(net342),
    .I1(_06170_),
    .S(_08425_),
    .Z(net213));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22315_ (.A1(_11647_[0]),
    .A2(_07449_),
    .B1(_07838_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(_08193_),
    .ZN(_06171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22316_ (.I(_06171_),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22317_ (.I0(net429),
    .I1(_06172_),
    .S(_08425_),
    .Z(net214));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22318_ (.A1(_11647_[0]),
    .A2(_07486_),
    .B1(_07875_),
    .B2(_11651_[0]),
    .C1(_11656_[0]),
    .C2(net430),
    .ZN(_06173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22319_ (.I(_06173_),
    .ZN(_06174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22320_ (.I0(net427),
    .I1(_06174_),
    .S(_08425_),
    .Z(net215));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22321_ (.A1(_11656_[0]),
    .A2(_06384_),
    .B1(_07544_),
    .B2(_11647_[0]),
    .C1(_07936_),
    .C2(_11651_[0]),
    .ZN(_06175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22322_ (.I(_06175_),
    .ZN(_06176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22323_ (.I0(net413),
    .I1(_06176_),
    .S(_08425_),
    .Z(net216));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22324_ (.A1(_11656_[0]),
    .A2(net468),
    .B1(_07582_),
    .B2(_11647_[0]),
    .C1(_07973_),
    .C2(_11651_[0]),
    .ZN(_06177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22325_ (.I(_06177_),
    .ZN(_06178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22326_ (.I0(net407),
    .I1(_06178_),
    .S(_08425_),
    .Z(net217));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22327_ (.A1(_01960_),
    .A2(_04392_),
    .Z(\id_stage_i.branch_set_d ));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22328_ (.A1(net128),
    .A2(_08669_),
    .Z(_06179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22329_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(_06179_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .ZN(_06180_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22330_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(_08669_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .ZN(_06181_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22331_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net128),
    .A3(_06181_),
    .Z(_06182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22332_ (.A1(net95),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .ZN(_06183_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22333_ (.A1(_06180_),
    .A2(_06182_),
    .B(_06183_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _22334_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net95),
    .Z(_06184_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22335_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .A2(_06184_),
    .ZN(_06185_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22336_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net128),
    .B1(_06181_),
    .B2(_06185_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22337_ (.A1(_05064_),
    .A2(_05095_),
    .B(_05075_),
    .ZN(_06186_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _22338_ (.A1(_05327_),
    .A2(_05064_),
    .A3(_05328_),
    .Z(_06187_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22339_ (.A1(net3651),
    .A2(_06187_),
    .ZN(_06188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22340_ (.A1(_08736_),
    .A2(_06186_),
    .B(_06188_),
    .C(_08669_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22341_ (.A1(_05065_),
    .A2(_05095_),
    .B1(_06187_),
    .B2(net3651),
    .C(_05100_),
    .ZN(_06189_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22342_ (.A1(_08669_),
    .A2(_06189_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22343_ (.A1(net3651),
    .A2(_05064_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .ZN(_06190_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _22344_ (.A1(_08669_),
    .A2(net3071),
    .A3(_06190_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22345_ (.A1(_08870_),
    .A2(net128),
    .ZN(_06191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22346_ (.A1(net95),
    .A2(net249),
    .B1(_06191_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .ZN(_06192_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22347_ (.I(_06192_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22348_ (.A1(net249),
    .A2(_06184_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .ZN(_06193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22349_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net128),
    .B(_06193_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22350_ (.A1(_05546_),
    .A2(net249),
    .Z(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22351_ (.A1(_08391_),
    .A2(_04372_),
    .Z(_06194_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _22352_ (.A1(_06345_),
    .A2(_04351_),
    .A3(_04381_),
    .A4(_06194_),
    .ZN(_06195_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22353_ (.A1(_08669_),
    .A2(_05069_),
    .ZN(_06196_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22354_ (.A1(_02019_),
    .A2(_04364_),
    .ZN(_06197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22355_ (.I0(_06195_),
    .I1(_06196_),
    .S(_06197_),
    .Z(\if_stage_i.instr_valid_id_d ));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22356_ (.A(_09746_[0]),
    .B(_09744_[0]),
    .CI(_09745_[0]),
    .CO(_09747_[0]),
    .S(_09748_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22357_ (.A(_09749_[0]),
    .B(_09750_[0]),
    .CI(_09751_[0]),
    .CO(_09752_[0]),
    .S(_09753_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22358_ (.A(_09754_[0]),
    .B(_09755_[0]),
    .CI(_09756_[0]),
    .CO(_09757_[0]),
    .S(_09758_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22359_ (.A(_09759_[0]),
    .B(_09760_[0]),
    .CI(_09761_[0]),
    .CO(_09762_[0]),
    .S(_09763_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22360_ (.A(_09764_[0]),
    .B(_09765_[0]),
    .CI(_09766_[0]),
    .CO(_09767_[0]),
    .S(_09768_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22361_ (.A(_09769_[0]),
    .B(_09757_[0]),
    .CI(_09768_[0]),
    .CO(_09770_[0]),
    .S(_09771_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22362_ (.A(_09772_[0]),
    .B(_09773_[0]),
    .CI(_09774_[0]),
    .CO(_09775_[0]),
    .S(_09776_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22363_ (.A(_09777_[0]),
    .B(_09778_[0]),
    .CI(_09779_[0]),
    .CO(_09780_[0]),
    .S(_09781_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22364_ (.A(_09782_[0]),
    .B(_09767_[0]),
    .CI(_09776_[0]),
    .CO(_09783_[0]),
    .S(_09784_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22365_ (.A(_09785_[0]),
    .B(_09786_[0]),
    .CI(_09787_[0]),
    .CO(_09788_[0]),
    .S(_09789_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22366_ (.A(_09790_[0]),
    .B(_09791_[0]),
    .CI(_09792_[0]),
    .CO(_09793_[0]),
    .S(_09794_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22367_ (.A(_09795_[0]),
    .B(_09796_[0]),
    .CI(_09797_[0]),
    .CO(_09798_[0]),
    .S(_09799_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22368_ (.A(_09799_[0]),
    .B(_09775_[0]),
    .CI(_09794_[0]),
    .CO(_09800_[0]),
    .S(_09801_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22369_ (.A(_09802_[0]),
    .B(_09783_[0]),
    .CI(_09801_[0]),
    .CO(_09803_[0]),
    .S(_09804_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22370_ (.A(_09806_[0]),
    .B(_09805_[0]),
    .CI(_09807_[0]),
    .CO(_09808_[0]),
    .S(_09809_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22371_ (.A(_09810_[0]),
    .B(_09811_[0]),
    .CI(_09812_[0]),
    .CO(_09813_[0]),
    .S(_09814_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22372_ (.A(_09809_[0]),
    .B(_09793_[0]),
    .CI(_09815_[0]),
    .CO(_09816_[0]),
    .S(_09817_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22373_ (.A(_09818_[0]),
    .B(_09800_[0]),
    .CI(_09817_[0]),
    .CO(_09819_[0]),
    .S(_09820_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22374_ (.A(_09821_[0]),
    .B(_09822_[0]),
    .CI(_09823_[0]),
    .CO(_09824_[0]),
    .S(_09825_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22375_ (.A(_09826_[0]),
    .B(_09827_[0]),
    .CI(_09828_[0]),
    .CO(_09829_[0]),
    .S(_09830_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22376_ (.A(_09831_[0]),
    .B(_09832_[0]),
    .CI(_09833_[0]),
    .CO(_09834_[0]),
    .S(_09835_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22377_ (.A(_09836_[0]),
    .B(_09808_[0]),
    .CI(_09830_[0]),
    .CO(_09837_[0]),
    .S(_09838_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22378_ (.A(_09839_[0]),
    .B(_09840_[0]),
    .CI(_09841_[0]),
    .CO(_09842_[0]),
    .S(_09843_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22379_ (.A(_09844_[0]),
    .B(_09845_[0]),
    .CI(_09813_[0]),
    .CO(_09846_[0]),
    .S(_09847_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22380_ (.A(_09848_[0]),
    .B(_09816_[0]),
    .CI(_09838_[0]),
    .CO(_09849_[0]),
    .S(_09850_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22381_ (.A(_09851_[0]),
    .B(_09852_[0]),
    .CI(_09853_[0]),
    .CO(_09854_[0]),
    .S(_09855_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22382_ (.A(_09858_[0]),
    .B(_09857_[0]),
    .CI(_09856_[0]),
    .CO(_09859_[0]),
    .S(_09860_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22383_ (.A(_09861_[0]),
    .B(_09862_[0]),
    .CI(_09863_[0]),
    .CO(_09864_[0]),
    .S(_09865_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22384_ (.A(_09866_[0]),
    .B(_09867_[0]),
    .CI(_09868_[0]),
    .CO(_09869_[0]),
    .S(_09870_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22385_ (.A(_09871_[0]),
    .B(_09829_[0]),
    .CI(_09865_[0]),
    .CO(_09872_[0]),
    .S(_09873_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22386_ (.A(_09874_[0]),
    .B(_09875_[0]),
    .CI(_09876_[0]),
    .CO(_09877_[0]),
    .S(_09878_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22387_ (.A(_09879_[0]),
    .B(_09880_[0]),
    .CI(_09834_[0]),
    .CO(_09881_[0]),
    .S(_09882_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22388_ (.A(_09883_[0]),
    .B(_09837_[0]),
    .CI(_09873_[0]),
    .CO(_09884_[0]),
    .S(_09885_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22389_ (.A(_09886_[0]),
    .B(_09849_[0]),
    .CI(_09885_[0]),
    .CO(_09887_[0]),
    .S(_09888_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22390_ (.A(_09889_[0]),
    .B(_09890_[0]),
    .CI(_09891_[0]),
    .CO(_09892_[0]),
    .S(_09893_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22391_ (.A(_09894_[0]),
    .B(_09895_[0]),
    .CI(_09896_[0]),
    .CO(_09897_[0]),
    .S(_09898_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22392_ (.A(_09899_[0]),
    .B(_09864_[0]),
    .CI(_09893_[0]),
    .CO(_09900_[0]),
    .S(_09901_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22393_ (.A(_09902_[0]),
    .B(_09903_[0]),
    .CI(_09904_[0]),
    .CO(_09905_[0]),
    .S(_09906_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22394_ (.A(_09907_[0]),
    .B(_09908_[0]),
    .CI(_09869_[0]),
    .CO(_09909_[0]),
    .S(_09910_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22395_ (.A(_09911_[0]),
    .B(_09872_[0]),
    .CI(_09901_[0]),
    .CO(_09912_[0]),
    .S(_09913_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22396_ (.A(_09914_[0]),
    .B(_09884_[0]),
    .CI(_09913_[0]),
    .CO(_09915_[0]),
    .S(_09916_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22397_ (.A(_09917_[0]),
    .B(_09918_[0]),
    .CI(_09919_[0]),
    .CO(_09920_[0]),
    .S(_09921_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22398_ (.A(_09922_[0]),
    .B(_09923_[0]),
    .CI(_09924_[0]),
    .CO(_09925_[0]),
    .S(_09926_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22399_ (.A(_09927_[0]),
    .B(_09928_[0]),
    .CI(_09929_[0]),
    .CO(_09930_[0]),
    .S(_09931_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22400_ (.A(_09932_[0]),
    .B(_09892_[0]),
    .CI(_09926_[0]),
    .CO(_09933_[0]),
    .S(_09934_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22401_ (.A(_09935_[0]),
    .B(_09936_[0]),
    .CI(_09937_[0]),
    .CO(_09938_[0]),
    .S(_09939_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22402_ (.A(_09905_[0]),
    .B(_09939_[0]),
    .CI(_09940_[0]),
    .CO(_09941_[0]),
    .S(_09942_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22403_ (.A(_09942_[0]),
    .B(_09900_[0]),
    .CI(_09934_[0]),
    .CO(_09943_[0]),
    .S(_09944_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22404_ (.A(_09945_[0]),
    .B(_09946_[0]),
    .CI(_09947_[0]),
    .CO(_09948_[0]),
    .S(_09949_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22405_ (.A(_09950_[0]),
    .B(_09912_[0]),
    .CI(_09944_[0]),
    .CO(_09951_[0]),
    .S(_09952_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22406_ (.A(_09953_[0]),
    .B(_09954_[0]),
    .CI(_09955_[0]),
    .CO(_09956_[0]),
    .S(_09957_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22407_ (.A(_09958_[0]),
    .B(_09959_[0]),
    .CI(_09960_[0]),
    .CO(_09961_[0]),
    .S(_09962_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22408_ (.A(_09963_[0]),
    .B(_09964_[0]),
    .CI(_09965_[0]),
    .CO(_09966_[0]),
    .S(_09967_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22409_ (.A(_09968_[0]),
    .B(_09925_[0]),
    .CI(_09962_[0]),
    .CO(_09969_[0]),
    .S(_09970_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22410_ (.A(_09971_[0]),
    .B(_09972_[0]),
    .CI(_09973_[0]),
    .CO(_09974_[0]),
    .S(_09975_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22411_ (.A(_09938_[0]),
    .B(_09975_[0]),
    .CI(_09976_[0]),
    .CO(_09977_[0]),
    .S(_09978_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22412_ (.A(_09978_[0]),
    .B(_09933_[0]),
    .CI(_09970_[0]),
    .CO(_09979_[0]),
    .S(_09980_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22413_ (.A(_09981_[0]),
    .B(_09982_[0]),
    .CI(_09983_[0]),
    .CO(_09984_[0]),
    .S(_09985_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22414_ (.A(_09986_[0]),
    .B(_09987_[0]),
    .CI(_09988_[0]),
    .CO(_09989_[0]),
    .S(_09990_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22415_ (.A(_09991_[0]),
    .B(_09990_[0]),
    .CI(_09992_[0]),
    .CO(_09993_[0]),
    .S(_09994_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22416_ (.A(_09995_[0]),
    .B(_09943_[0]),
    .CI(_09980_[0]),
    .CO(_09996_[0]),
    .S(_09997_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22417_ (.A(_09998_[0]),
    .B(_09999_[0]),
    .CI(_10000_[0]),
    .CO(_10001_[0]),
    .S(_10002_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22418_ (.A(_10003_[0]),
    .B(_10004_[0]),
    .CI(_10005_[0]),
    .CO(_10006_[0]),
    .S(_10007_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22419_ (.A(_10008_[0]),
    .B(_10009_[0]),
    .CI(_10010_[0]),
    .CO(_10011_[0]),
    .S(_10012_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22420_ (.A(_10013_[0]),
    .B(_09961_[0]),
    .CI(_10007_[0]),
    .CO(_10014_[0]),
    .S(_10015_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22421_ (.A(_10016_[0]),
    .B(_10017_[0]),
    .CI(_10018_[0]),
    .CO(_10019_[0]),
    .S(_10020_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22422_ (.A(_09974_[0]),
    .B(_10020_[0]),
    .CI(_10021_[0]),
    .CO(_10022_[0]),
    .S(_10023_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22423_ (.A(_10023_[0]),
    .B(_09969_[0]),
    .CI(_10015_[0]),
    .CO(_10024_[0]),
    .S(_10025_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22424_ (.A(_10026_[0]),
    .B(_10027_[0]),
    .CI(_10028_[0]),
    .CO(_10029_[0]),
    .S(_10030_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22425_ (.A(_10031_[0]),
    .B(_09984_[0]),
    .CI(_10030_[0]),
    .CO(_10032_[0]),
    .S(_10033_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22426_ (.A(_10034_[0]),
    .B(_10033_[0]),
    .CI(_09977_[0]),
    .CO(_10035_[0]),
    .S(_10036_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22427_ (.A(_10036_[0]),
    .B(_09979_[0]),
    .CI(_10025_[0]),
    .CO(_10037_[0]),
    .S(_10038_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22428_ (.A(_10039_[0]),
    .B(_09996_[0]),
    .CI(_10038_[0]),
    .CO(_10040_[0]),
    .S(_10041_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22429_ (.A(_10042_[0]),
    .B(_10043_[0]),
    .CI(_10044_[0]),
    .CO(_10045_[0]),
    .S(_10046_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22430_ (.A(_10047_[0]),
    .B(_10048_[0]),
    .CI(_10049_[0]),
    .CO(_10050_[0]),
    .S(_10051_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22431_ (.A(_10006_[0]),
    .B(_10046_[0]),
    .CI(_10052_[0]),
    .CO(_10053_[0]),
    .S(_10054_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22432_ (.A(_10055_[0]),
    .B(_10056_[0]),
    .CI(_10057_[0]),
    .CO(_10058_[0]),
    .S(_10059_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22433_ (.A(_10019_[0]),
    .B(_10059_[0]),
    .CI(_10060_[0]),
    .CO(_10061_[0]),
    .S(_10062_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22434_ (.A(_10062_[0]),
    .B(_10014_[0]),
    .CI(_10054_[0]),
    .CO(_10063_[0]),
    .S(_10064_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22435_ (.A(_10065_[0]),
    .B(_10066_[0]),
    .CI(_10067_[0]),
    .CO(_10068_[0]),
    .S(_10069_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22436_ (.A(_10070_[0]),
    .B(_10071_[0]),
    .CI(_10072_[0]),
    .CO(_10073_[0]),
    .S(_10074_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22437_ (.A(_10069_[0]),
    .B(_10029_[0]),
    .CI(_10075_[0]),
    .CO(_10076_[0]),
    .S(_10077_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22438_ (.A(_10078_[0]),
    .B(_10080_[0]),
    .CI(_10079_[0]),
    .CO(_10081_[0]),
    .S(_10082_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22439_ (.A(_10083_[0]),
    .B(_10024_[0]),
    .CI(_10064_[0]),
    .CO(_10084_[0]),
    .S(_10085_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22440_ (.A(_10086_[0]),
    .B(_10037_[0]),
    .CI(_10085_[0]),
    .CO(_10087_[0]),
    .S(_10088_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22441_ (.A(_10089_[0]),
    .B(_10090_[0]),
    .CI(_10091_[0]),
    .CO(_10092_[0]),
    .S(_10093_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22442_ (.A(_10094_[0]),
    .B(_10095_[0]),
    .CI(_10096_[0]),
    .CO(_10097_[0]),
    .S(_10098_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22443_ (.A(_10098_[0]),
    .B(_10045_[0]),
    .CI(_10093_[0]),
    .CO(_10099_[0]),
    .S(_10100_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22444_ (.A(_10101_[0]),
    .B(_10102_[0]),
    .CI(_10103_[0]),
    .CO(_10104_[0]),
    .S(_10105_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22445_ (.A(_10058_[0]),
    .B(_10105_[0]),
    .CI(_10106_[0]),
    .CO(_10107_[0]),
    .S(_10108_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22446_ (.A(_10053_[0]),
    .B(_10108_[0]),
    .CI(_10100_[0]),
    .CO(_10109_[0]),
    .S(_10110_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22447_ (.A(_10111_[0]),
    .B(_10112_[0]),
    .CI(_10113_[0]),
    .CO(_10114_[0]),
    .S(_10115_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22448_ (.A(_10118_[0]),
    .B(_10117_[0]),
    .CI(_10116_[0]),
    .CO(_10119_[0]),
    .S(_10120_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22449_ (.A(_10115_[0]),
    .B(_10068_[0]),
    .CI(_10121_[0]),
    .CO(_10122_[0]),
    .S(_10123_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22450_ (.A(_10124_[0]),
    .B(_10126_[0]),
    .CI(_10125_[0]),
    .CO(_10127_[0]),
    .S(_10128_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22451_ (.A(_10110_[0]),
    .B(_10063_[0]),
    .CI(_10129_[0]),
    .CO(_10130_[0]),
    .S(_10131_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22452_ (.A(_10131_[0]),
    .B(_10084_[0]),
    .CI(_10132_[0]),
    .CO(_10133_[0]),
    .S(_10134_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22453_ (.A(_10137_[0]),
    .B(_10136_[0]),
    .CI(_10135_[0]),
    .CO(_10138_[0]),
    .S(_10139_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22454_ (.A(_10140_[0]),
    .B(_10141_[0]),
    .CI(_10142_[0]),
    .CO(_10143_[0]),
    .S(_10144_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22455_ (.A(_10145_[0]),
    .B(_10146_[0]),
    .CI(_10147_[0]),
    .CO(_10148_[0]),
    .S(_10149_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22456_ (.A(_10150_[0]),
    .B(_10092_[0]),
    .CI(_10144_[0]),
    .CO(_10151_[0]),
    .S(_10152_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22457_ (.A(_10153_[0]),
    .B(_10154_[0]),
    .CI(_10155_[0]),
    .CO(_10156_[0]),
    .S(_10157_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22458_ (.A(_10104_[0]),
    .B(_10157_[0]),
    .CI(_10097_[0]),
    .CO(_10158_[0]),
    .S(_10159_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22459_ (.A(_10159_[0]),
    .B(_10099_[0]),
    .CI(_10152_[0]),
    .CO(_10160_[0]),
    .S(_10161_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22460_ (.A(_10162_[0]),
    .B(_10163_[0]),
    .CI(_10164_[0]),
    .CO(_10165_[0]),
    .S(_10166_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22461_ (.A(_10167_[0]),
    .B(_10168_[0]),
    .CI(_10169_[0]),
    .CO(_10170_[0]),
    .S(_10171_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22462_ (.A(_10172_[0]),
    .B(_10114_[0]),
    .CI(_10166_[0]),
    .CO(_10173_[0]),
    .S(_10174_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22463_ (.A(_10122_[0]),
    .B(_10174_[0]),
    .CI(_10107_[0]),
    .CO(_10175_[0]),
    .S(_10176_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22464_ (.A(_10176_[0]),
    .B(_10109_[0]),
    .CI(_10161_[0]),
    .CO(_10177_[0]),
    .S(_10178_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22465_ (.A(_10179_[0]),
    .B(_10130_[0]),
    .CI(_10178_[0]),
    .CO(_10180_[0]),
    .S(_10181_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22466_ (.A(_10182_[0]),
    .B(_10183_[0]),
    .CI(_10184_[0]),
    .CO(_10185_[0]),
    .S(_10186_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22467_ (.A(_10187_[0]),
    .B(_10188_[0]),
    .CI(_10189_[0]),
    .CO(_10190_[0]),
    .S(_10191_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22468_ (.A(_10192_[0]),
    .B(_10193_[0]),
    .CI(_10194_[0]),
    .CO(_10195_[0]),
    .S(_10196_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22469_ (.A(_10197_[0]),
    .B(_10143_[0]),
    .CI(_10198_[0]),
    .CO(_10199_[0]),
    .S(_10200_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22470_ (.A(_10201_[0]),
    .B(_10202_[0]),
    .CI(_10203_[0]),
    .CO(_10204_[0]),
    .S(_10205_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22471_ (.A(_10156_[0]),
    .B(_10205_[0]),
    .CI(_10206_[0]),
    .CO(_10207_[0]),
    .S(_10208_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22472_ (.A(_10208_[0]),
    .B(_10151_[0]),
    .CI(_10200_[0]),
    .CO(_10209_[0]),
    .S(_10210_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22473_ (.A(_10211_[0]),
    .B(_10212_[0]),
    .CI(_10213_[0]),
    .CO(_10214_[0]),
    .S(_10215_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22474_ (.A(_10216_[0]),
    .B(_10217_[0]),
    .CI(_10218_[0]),
    .CO(_10219_[0]),
    .S(_10220_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22475_ (.A(_10221_[0]),
    .B(_10165_[0]),
    .CI(_10215_[0]),
    .CO(_10222_[0]),
    .S(_10223_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22476_ (.A(_10223_[0]),
    .B(_10173_[0]),
    .CI(_10158_[0]),
    .CO(_10224_[0]),
    .S(_10225_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22477_ (.A(_10225_[0]),
    .B(_10160_[0]),
    .CI(_10210_[0]),
    .CO(_10226_[0]),
    .S(_10227_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22478_ (.A(_10228_[0]),
    .B(_10229_[0]),
    .CI(_10230_[0]),
    .CO(_10231_[0]),
    .S(_10232_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22479_ (.A(_10233_[0]),
    .B(_10234_[0]),
    .CI(_10170_[0]),
    .CO(_10235_[0]),
    .S(_10236_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22480_ (.A(_10237_[0]),
    .B(_10238_[0]),
    .CI(_10239_[0]),
    .CO(_10240_[0]),
    .S(_10241_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22481_ (.A(_10242_[0]),
    .B(_10243_[0]),
    .CI(_10244_[0]),
    .CO(_10245_[0]),
    .S(_10246_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22482_ (.A(_10177_[0]),
    .B(_10227_[0]),
    .CI(_10247_[0]),
    .CO(_10248_[0]),
    .S(_10249_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22483_ (.A(_10250_[0]),
    .B(_10251_[0]),
    .CI(_10252_[0]),
    .CO(_10253_[0]),
    .S(_10254_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22484_ (.A(_10255_[0]),
    .B(_10256_[0]),
    .CI(_10187_[0]),
    .CO(_10257_[0]),
    .S(_10258_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22485_ (.A(_10259_[0]),
    .B(_10260_[0]),
    .CI(_10261_[0]),
    .CO(_10262_[0]),
    .S(_10263_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22486_ (.A(_10264_[0]),
    .B(_10265_[0]),
    .CI(_10266_[0]),
    .CO(_10267_[0]),
    .S(_10268_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22487_ (.A(_10269_[0]),
    .B(_10270_[0]),
    .CI(_10271_[0]),
    .CO(_10272_[0]),
    .S(_10273_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22488_ (.A(_10204_[0]),
    .B(_10273_[0]),
    .CI(_10274_[0]),
    .CO(_10275_[0]),
    .S(_10276_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22489_ (.A(_10276_[0]),
    .B(_10199_[0]),
    .CI(_10268_[0]),
    .CO(_10277_[0]),
    .S(_10278_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22490_ (.A(_10279_[0]),
    .B(_10280_[0]),
    .CI(_10281_[0]),
    .CO(_10282_[0]),
    .S(_10283_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22491_ (.A(_10284_[0]),
    .B(_10285_[0]),
    .CI(_10286_[0]),
    .CO(_10287_[0]),
    .S(_10288_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22492_ (.A(_10289_[0]),
    .B(_10214_[0]),
    .CI(_10283_[0]),
    .CO(_10290_[0]),
    .S(_10291_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22493_ (.A(_10222_[0]),
    .B(_10291_[0]),
    .CI(_10207_[0]),
    .CO(_10292_[0]),
    .S(_10293_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22494_ (.A(_10293_[0]),
    .B(_10209_[0]),
    .CI(_10278_[0]),
    .CO(_10294_[0]),
    .S(_10295_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22495_ (.A(_10296_[0]),
    .B(_10297_[0]),
    .CI(_10298_[0]),
    .CO(_10299_[0]),
    .S(_10300_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22496_ (.A(_10231_[0]),
    .B(_10300_[0]),
    .CI(_10301_[0]),
    .CO(_10302_[0]),
    .S(_10303_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22497_ (.A(_10240_[0]),
    .B(_10304_[0]),
    .CI(_10224_[0]),
    .CO(_10305_[0]),
    .S(_10306_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22498_ (.A(_10226_[0]),
    .B(_10295_[0]),
    .CI(_10306_[0]),
    .CO(_10307_[0]),
    .S(_10308_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22499_ (.A(_10309_[0]),
    .B(_10248_[0]),
    .CI(_10308_[0]),
    .CO(_10310_[0]),
    .S(_10311_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22500_ (.A(_10255_[0]),
    .B(_10187_[0]),
    .CI(_10312_[0]),
    .CO(_10313_[0]),
    .S(_10314_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22501_ (.A(_10315_[0]),
    .B(_10316_[0]),
    .CI(_10317_[0]),
    .CO(_10318_[0]),
    .S(_10319_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22502_ (.A(_10320_[0]),
    .B(_10321_[0]),
    .CI(_10322_[0]),
    .CO(_10323_[0]),
    .S(_10324_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22503_ (.A(_10325_[0]),
    .B(_10326_[0]),
    .CI(_10327_[0]),
    .CO(_10328_[0]),
    .S(_10329_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22504_ (.A(_10272_[0]),
    .B(_10329_[0]),
    .CI(_10330_[0]),
    .CO(_10331_[0]),
    .S(_10332_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22505_ (.A(_10332_[0]),
    .B(_10267_[0]),
    .CI(_10324_[0]),
    .CO(_10333_[0]),
    .S(_10334_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22506_ (.A(_10335_[0]),
    .B(_10336_[0]),
    .CI(_10337_[0]),
    .CO(_10338_[0]),
    .S(_10339_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22507_ (.A(_10340_[0]),
    .B(_10341_[0]),
    .CI(_10342_[0]),
    .CO(_10343_[0]),
    .S(_10344_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22508_ (.A(_10345_[0]),
    .B(_10282_[0]),
    .CI(_10339_[0]),
    .CO(_10346_[0]),
    .S(_10347_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22509_ (.A(_10290_[0]),
    .B(_10347_[0]),
    .CI(_10275_[0]),
    .CO(_10348_[0]),
    .S(_10349_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22510_ (.A(_10349_[0]),
    .B(_10277_[0]),
    .CI(_10334_[0]),
    .CO(_10350_[0]),
    .S(_10351_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22511_ (.A(_10352_[0]),
    .B(_10353_[0]),
    .CI(_10354_[0]),
    .CO(_10355_[0]),
    .S(_10356_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22512_ (.A(_10299_[0]),
    .B(_10356_[0]),
    .CI(_10357_[0]),
    .CO(_10358_[0]),
    .S(_10359_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22513_ (.A(_10360_[0]),
    .B(_10361_[0]),
    .CI(_10362_[0]),
    .CO(_10363_[0]),
    .S(_10364_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22514_ (.A(_10294_[0]),
    .B(_10351_[0]),
    .CI(_10365_[0]),
    .CO(_10366_[0]),
    .S(_10367_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22515_ (.A(_10305_[0]),
    .B(_10307_[0]),
    .CI(_10367_[0]),
    .CO(_10368_[0]),
    .S(_10369_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22516_ (.A(_10255_[0]),
    .B(net476),
    .CI(_10370_[0]),
    .CO(_10371_[0]),
    .S(_10372_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22517_ (.A(_10373_[0]),
    .B(_10374_[0]),
    .CI(_10317_[0]),
    .CO(_10375_[0]),
    .S(_10376_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22518_ (.A(_10377_[0]),
    .B(_10378_[0]),
    .CI(_10379_[0]),
    .CO(_10380_[0]),
    .S(_10381_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22519_ (.A(_10382_[0]),
    .B(_10383_[0]),
    .CI(_10384_[0]),
    .CO(_10385_[0]),
    .S(_10386_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22520_ (.A(_10328_[0]),
    .B(_10386_[0]),
    .CI(_10387_[0]),
    .CO(_10388_[0]),
    .S(_10389_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22521_ (.A(_10389_[0]),
    .B(_10323_[0]),
    .CI(_10381_[0]),
    .CO(_10390_[0]),
    .S(_10391_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22522_ (.A(_10392_[0]),
    .B(_10393_[0]),
    .CI(_10394_[0]),
    .CO(_10395_[0]),
    .S(_10396_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22523_ (.A(_10397_[0]),
    .B(_10398_[0]),
    .CI(_10399_[0]),
    .CO(_10400_[0]),
    .S(_10401_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22524_ (.A(_10402_[0]),
    .B(_10338_[0]),
    .CI(_10396_[0]),
    .CO(_10403_[0]),
    .S(_10404_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22525_ (.A(_10331_[0]),
    .B(_10346_[0]),
    .CI(_10404_[0]),
    .CO(_10405_[0]),
    .S(_10406_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22526_ (.A(_10333_[0]),
    .B(_10391_[0]),
    .CI(_10406_[0]),
    .CO(_10407_[0]),
    .S(_10408_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22527_ (.A(_10409_[0]),
    .B(_10410_[0]),
    .CI(_10411_[0]),
    .CO(_10412_[0]),
    .S(_10413_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22528_ (.A(_10355_[0]),
    .B(_10413_[0]),
    .CI(_10414_[0]),
    .CO(_10415_[0]),
    .S(_10416_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22529_ (.A(_10417_[0]),
    .B(_10418_[0]),
    .CI(_10419_[0]),
    .CO(_10420_[0]),
    .S(_10421_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22530_ (.A(_10422_[0]),
    .B(_10350_[0]),
    .CI(_10408_[0]),
    .CO(_10423_[0]),
    .S(_10424_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22531_ (.A(_10425_[0]),
    .B(_10366_[0]),
    .CI(_10424_[0]),
    .CO(_10426_[0]),
    .S(_10427_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22532_ (.A(net3227),
    .B(net476),
    .CI(_10428_[0]),
    .CO(_10429_[0]),
    .S(_10430_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22533_ (.A(_10374_[0]),
    .B(_10431_[0]),
    .CI(_10317_[0]),
    .CO(_10432_[0]),
    .S(_10433_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22534_ (.A(_10433_[0]),
    .B(_10371_[0]),
    .CI(_10430_[0]),
    .CO(_10434_[0]),
    .S(_10435_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22535_ (.A(_10437_[0]),
    .B(_10438_[0]),
    .CI(_10439_[0]),
    .CO(_10440_[0]),
    .S(_10441_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22536_ (.A(_10385_[0]),
    .B(_10441_[0]),
    .CI(_10442_[0]),
    .CO(_10443_[0]),
    .S(_10444_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22537_ (.A(_10444_[0]),
    .B(_10380_[0]),
    .CI(_10445_[0]),
    .CO(_10446_[0]),
    .S(_10447_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22538_ (.A(_10448_[0]),
    .B(_10449_[0]),
    .CI(_10450_[0]),
    .CO(_10451_[0]),
    .S(_10452_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22539_ (.A(_10453_[0]),
    .B(_10454_[0]),
    .CI(_10455_[0]),
    .CO(_10456_[0]),
    .S(_10457_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22540_ (.A(_10395_[0]),
    .B(_10452_[0]),
    .CI(_10458_[0]),
    .CO(_10459_[0]),
    .S(_10460_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22541_ (.A(_10388_[0]),
    .B(_10403_[0]),
    .CI(_10460_[0]),
    .CO(_10461_[0]),
    .S(_10462_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22542_ (.A(_10390_[0]),
    .B(_10447_[0]),
    .CI(_10462_[0]),
    .CO(_10463_[0]),
    .S(_10464_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22543_ (.A(_10465_[0]),
    .B(_10466_[0]),
    .CI(_10467_[0]),
    .CO(_10468_[0]),
    .S(_10469_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22544_ (.A(_10412_[0]),
    .B(_10469_[0]),
    .CI(_10470_[0]),
    .CO(_10471_[0]),
    .S(_10472_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22545_ (.A(_10473_[0]),
    .B(_10474_[0]),
    .CI(_10475_[0]),
    .CO(_10476_[0]),
    .S(_10477_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22546_ (.A(_10478_[0]),
    .B(_10407_[0]),
    .CI(_10464_[0]),
    .CO(_10479_[0]),
    .S(_10480_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22547_ (.A(_10481_[0]),
    .B(_10423_[0]),
    .CI(_10480_[0]),
    .CO(_10482_[0]),
    .S(_10483_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22548_ (.A(net3228),
    .B(net3232),
    .CI(_10484_[0]),
    .CO(_10485_[0]),
    .S(_10486_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22549_ (.A(_10488_[0]),
    .B(_10487_[0]),
    .CI(_10436_[0]),
    .CO(_10489_[0]),
    .S(_10490_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22550_ (.A(_10491_[0]),
    .B(_10492_[0]),
    .CI(net3226),
    .CO(_10494_[0]),
    .S(_10495_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22551_ (.A(_10496_[0]),
    .B(net3212),
    .CI(_10440_[0]),
    .CO(_10498_[0]),
    .S(_10499_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22552_ (.A(_10490_[0]),
    .B(_10500_[0]),
    .CI(_10499_[0]),
    .CO(_10501_[0]),
    .S(_10502_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22553_ (.A(_10503_[0]),
    .B(_10504_[0]),
    .CI(_10505_[0]),
    .CO(_10506_[0]),
    .S(_10507_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22554_ (.A(_10508_[0]),
    .B(_10509_[0]),
    .CI(_10510_[0]),
    .CO(_10511_[0]),
    .S(_10512_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22555_ (.A(_10513_[0]),
    .B(_10451_[0]),
    .CI(_10507_[0]),
    .CO(_10514_[0]),
    .S(_10515_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22556_ (.A(_10459_[0]),
    .B(_10515_[0]),
    .CI(_10443_[0]),
    .CO(_10516_[0]),
    .S(_10517_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22557_ (.A(_10502_[0]),
    .B(_10446_[0]),
    .CI(_10517_[0]),
    .CO(_10518_[0]),
    .S(_10519_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22558_ (.A(_10520_[0]),
    .B(_10521_[0]),
    .CI(_10522_[0]),
    .CO(_10523_[0]),
    .S(_10524_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22559_ (.A(_10468_[0]),
    .B(_10524_[0]),
    .CI(_10525_[0]),
    .CO(_10526_[0]),
    .S(_10527_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22560_ (.A(_10528_[0]),
    .B(_10529_[0]),
    .CI(_10530_[0]),
    .CO(_10531_[0]),
    .S(_10532_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22561_ (.A(_10533_[0]),
    .B(_10463_[0]),
    .CI(_10519_[0]),
    .CO(_10534_[0]),
    .S(_10535_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22562_ (.A(_10536_[0]),
    .B(_10479_[0]),
    .CI(_10535_[0]),
    .CO(_10537_[0]),
    .S(_10538_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22563_ (.A(net3228),
    .B(net3232),
    .CI(_10539_[0]),
    .CO(_10540_[0]),
    .S(_10541_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22564_ (.A(net3216),
    .B(_10485_[0]),
    .CI(_10541_[0]),
    .CO(_10542_[0]),
    .S(_10543_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22565_ (.A(net3226),
    .B(_10544_[0]),
    .CI(net3225),
    .CO(_10546_[0]),
    .S(_10547_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22566_ (.A(net3212),
    .B(_10548_[0]),
    .CI(_10549_[0]),
    .CO(_10550_[0]),
    .S(_10551_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22567_ (.A(_10551_[0]),
    .B(_10489_[0]),
    .CI(_10552_[0]),
    .CO(_10553_[0]),
    .S(_10554_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22568_ (.A(_10555_[0]),
    .B(_10556_[0]),
    .CI(_10557_[0]),
    .CO(_10558_[0]),
    .S(_10559_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22569_ (.A(_10560_[0]),
    .B(_10561_[0]),
    .CI(_10562_[0]),
    .CO(_10563_[0]),
    .S(_10564_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22570_ (.A(_10565_[0]),
    .B(_10506_[0]),
    .CI(_10559_[0]),
    .CO(_10566_[0]),
    .S(_10567_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22571_ (.A(_10514_[0]),
    .B(_10567_[0]),
    .CI(_10498_[0]),
    .CO(_10568_[0]),
    .S(_10569_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22572_ (.A(_10569_[0]),
    .B(_10501_[0]),
    .CI(_10554_[0]),
    .CO(_10570_[0]),
    .S(_10571_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22573_ (.A(_10572_[0]),
    .B(_10573_[0]),
    .CI(_10574_[0]),
    .CO(_10575_[0]),
    .S(_10576_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22574_ (.A(_10523_[0]),
    .B(_10576_[0]),
    .CI(_10577_[0]),
    .CO(_10578_[0]),
    .S(_10579_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22575_ (.A(_10580_[0]),
    .B(_10581_[0]),
    .CI(_10582_[0]),
    .CO(_10583_[0]),
    .S(_10584_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22576_ (.A(_10585_[0]),
    .B(_10518_[0]),
    .CI(_10571_[0]),
    .CO(_10586_[0]),
    .S(_10587_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22577_ (.A(_10588_[0]),
    .B(_10534_[0]),
    .CI(_10587_[0]),
    .CO(_10589_[0]),
    .S(_10590_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22578_ (.A(net3228),
    .B(net3232),
    .CI(_10591_[0]),
    .CO(_10592_[0]),
    .S(_10593_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22579_ (.A(_10594_[0]),
    .B(_10595_[0]),
    .CI(_10436_[0]),
    .CO(_10596_[0]),
    .S(_10597_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22580_ (.A(_10598_[0]),
    .B(_10493_[0]),
    .CI(_10545_[0]),
    .CO(_10599_[0]),
    .S(_10600_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22581_ (.A(_10601_[0]),
    .B(net3213),
    .CI(net3212),
    .CO(_10603_[0]),
    .S(_10604_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22582_ (.A(_10605_[0]),
    .B(_10597_[0]),
    .CI(_10604_[0]),
    .CO(_10606_[0]),
    .S(_10607_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22583_ (.A(_10608_[0]),
    .B(_10609_[0]),
    .CI(_10610_[0]),
    .CO(_10611_[0]),
    .S(_10612_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22584_ (.A(_10613_[0]),
    .B(_10614_[0]),
    .CI(_10615_[0]),
    .CO(_10616_[0]),
    .S(_10617_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22585_ (.A(_10618_[0]),
    .B(_10558_[0]),
    .CI(_10612_[0]),
    .CO(_10619_[0]),
    .S(_10620_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22586_ (.A(_10566_[0]),
    .B(_10620_[0]),
    .CI(_10550_[0]),
    .CO(_10621_[0]),
    .S(_10622_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22587_ (.A(_10622_[0]),
    .B(_10553_[0]),
    .CI(_10607_[0]),
    .CO(_10623_[0]),
    .S(_10624_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22588_ (.A(_10625_[0]),
    .B(_10626_[0]),
    .CI(_10627_[0]),
    .CO(_10628_[0]),
    .S(_10629_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22589_ (.A(_10575_[0]),
    .B(_10629_[0]),
    .CI(_10630_[0]),
    .CO(_10631_[0]),
    .S(_10632_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22590_ (.A(_10633_[0]),
    .B(_10634_[0]),
    .CI(_10635_[0]),
    .CO(_10636_[0]),
    .S(_10637_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22591_ (.A(_10638_[0]),
    .B(_10570_[0]),
    .CI(_10624_[0]),
    .CO(_10639_[0]),
    .S(_10640_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22592_ (.A(_10641_[0]),
    .B(_10586_[0]),
    .CI(_10640_[0]),
    .CO(_10642_[0]),
    .S(_10643_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22593_ (.A(net3228),
    .B(net3232),
    .CI(_10644_[0]),
    .CO(_10645_[0]),
    .S(_10646_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22594_ (.A(net3216),
    .B(_10592_[0]),
    .CI(_10646_[0]),
    .CO(_10647_[0]),
    .S(_10648_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22595_ (.A(_10602_[0]),
    .B(_10497_[0]),
    .CI(_10649_[0]),
    .CO(_10650_[0]),
    .S(_10651_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22596_ (.A(_10652_[0]),
    .B(_10653_[0]),
    .CI(_10648_[0]),
    .CO(_10654_[0]),
    .S(_10655_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22597_ (.A(_10656_[0]),
    .B(_10657_[0]),
    .CI(_10658_[0]),
    .CO(_10659_[0]),
    .S(_10660_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22598_ (.A(_10661_[0]),
    .B(_10662_[0]),
    .CI(_10663_[0]),
    .CO(_10664_[0]),
    .S(_10665_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22599_ (.A(_10666_[0]),
    .B(_10611_[0]),
    .CI(_10667_[0]),
    .CO(_10668_[0]),
    .S(_10669_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22600_ (.A(_10669_[0]),
    .B(_10603_[0]),
    .CI(_10619_[0]),
    .CO(_10670_[0]),
    .S(_10671_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22601_ (.A(_10606_[0]),
    .B(_10672_[0]),
    .CI(_10671_[0]),
    .CO(_10673_[0]),
    .S(_10674_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22602_ (.A(_10675_[0]),
    .B(_10676_[0]),
    .CI(_10677_[0]),
    .CO(_10678_[0]),
    .S(_10679_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22603_ (.A(_10628_[0]),
    .B(_10679_[0]),
    .CI(_10680_[0]),
    .CO(_10681_[0]),
    .S(_10682_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22604_ (.A(_10683_[0]),
    .B(_10684_[0]),
    .CI(_10685_[0]),
    .CO(_10686_[0]),
    .S(_10687_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22605_ (.A(_10688_[0]),
    .B(_10623_[0]),
    .CI(_10674_[0]),
    .CO(_10689_[0]),
    .S(_10690_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22606_ (.A(_10691_[0]),
    .B(_10639_[0]),
    .CI(_10690_[0]),
    .CO(_10692_[0]),
    .S(_10693_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22607_ (.A(net3228),
    .B(net3234),
    .CI(_10694_[0]),
    .CO(_10695_[0]),
    .S(_10696_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22608_ (.A(net3216),
    .B(_10645_[0]),
    .CI(_10696_[0]),
    .CO(_10697_[0]),
    .S(_10698_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22609_ (.A(_10699_[0]),
    .B(_10700_[0]),
    .CI(net3203),
    .CO(_10701_[0]),
    .S(_10702_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22610_ (.A(_10703_[0]),
    .B(_10704_[0]),
    .CI(_10658_[0]),
    .CO(_10705_[0]),
    .S(_10706_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22611_ (.A(_10707_[0]),
    .B(_10708_[0]),
    .CI(_10709_[0]),
    .CO(_10710_[0]),
    .S(_10711_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22612_ (.A(_10712_[0]),
    .B(_10713_[0]),
    .CI(_10714_[0]),
    .CO(_10715_[0]),
    .S(_10716_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22613_ (.A(_10650_[0]),
    .B(_10668_[0]),
    .CI(_10716_[0]),
    .CO(_10717_[0]),
    .S(_10718_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22614_ (.A(_10719_[0]),
    .B(_10702_[0]),
    .CI(_10718_[0]),
    .CO(_10720_[0]),
    .S(_10721_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22615_ (.A(_10722_[0]),
    .B(_10723_[0]),
    .CI(_10724_[0]),
    .CO(_10725_[0]),
    .S(_10726_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22616_ (.A(_10678_[0]),
    .B(_10726_[0]),
    .CI(_10727_[0]),
    .CO(_10728_[0]),
    .S(_10729_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22617_ (.A(_10730_[0]),
    .B(_10731_[0]),
    .CI(_10732_[0]),
    .CO(_10733_[0]),
    .S(_10734_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22618_ (.A(_10735_[0]),
    .B(_10673_[0]),
    .CI(_10721_[0]),
    .CO(_10736_[0]),
    .S(_10737_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22619_ (.A(_10738_[0]),
    .B(_10689_[0]),
    .CI(_10737_[0]),
    .CO(_10739_[0]),
    .S(_10740_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22620_ (.A(net3229),
    .B(net3233),
    .CI(_10741_[0]),
    .CO(_10742_[0]),
    .S(_10743_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22621_ (.A(net3217),
    .B(_10695_[0]),
    .CI(_10743_[0]),
    .CO(_10744_[0]),
    .S(_10745_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22622_ (.A(net3202),
    .B(_10697_[0]),
    .CI(_10745_[0]),
    .CO(_10746_[0]),
    .S(_10747_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22623_ (.A(_10704_[0]),
    .B(_10658_[0]),
    .CI(_10748_[0]),
    .CO(_10749_[0]),
    .S(_10750_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22624_ (.A(_10751_[0]),
    .B(_10752_[0]),
    .CI(_10753_[0]),
    .CO(_10754_[0]),
    .S(_10755_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22625_ (.A(_10756_[0]),
    .B(_10757_[0]),
    .CI(_10758_[0]),
    .CO(_10759_[0]),
    .S(_10760_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22626_ (.A(net3205),
    .B(_10715_[0]),
    .CI(_10760_[0]),
    .CO(_10761_[0]),
    .S(_10762_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22627_ (.A(_10762_[0]),
    .B(_10701_[0]),
    .CI(_10763_[0]),
    .CO(_10764_[0]),
    .S(_10765_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22628_ (.A(_10766_[0]),
    .B(_10767_[0]),
    .CI(_10768_[0]),
    .CO(_10769_[0]),
    .S(_10770_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22629_ (.A(_10725_[0]),
    .B(_10770_[0]),
    .CI(_10771_[0]),
    .CO(_10772_[0]),
    .S(_10773_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22630_ (.A(_10774_[0]),
    .B(_10775_[0]),
    .CI(_10776_[0]),
    .CO(_10777_[0]),
    .S(_10778_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22631_ (.A(_10720_[0]),
    .B(_10765_[0]),
    .CI(_10779_[0]),
    .CO(_10780_[0]),
    .S(_10781_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22632_ (.A(_10782_[0]),
    .B(_10736_[0]),
    .CI(_10781_[0]),
    .CO(_10783_[0]),
    .S(_10784_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22633_ (.A(net3229),
    .B(net3233),
    .CI(_10785_[0]),
    .CO(_10786_[0]),
    .S(_10787_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22634_ (.A(net3217),
    .B(_10742_[0]),
    .CI(_10787_[0]),
    .CO(_10788_[0]),
    .S(_10789_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22635_ (.A(net3202),
    .B(_10744_[0]),
    .CI(_10789_[0]),
    .CO(_10790_[0]),
    .S(_10791_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22636_ (.A(_10792_[0]),
    .B(_10793_[0]),
    .CI(_10794_[0]),
    .CO(_10795_[0]),
    .S(_10796_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22637_ (.A(_10797_[0]),
    .B(_10758_[0]),
    .CI(_10798_[0]),
    .CO(_10799_[0]),
    .S(_10800_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22638_ (.A(net3205),
    .B(_10759_[0]),
    .CI(_10800_[0]),
    .CO(_10801_[0]),
    .S(_10802_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22639_ (.A(_10802_[0]),
    .B(_10803_[0]),
    .CI(_10804_[0]),
    .CO(_10805_[0]),
    .S(_10806_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22640_ (.A(_10807_[0]),
    .B(_10808_[0]),
    .CI(_10809_[0]),
    .CO(_10810_[0]),
    .S(_10811_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22641_ (.A(_10769_[0]),
    .B(_10811_[0]),
    .CI(_10812_[0]),
    .CO(_10813_[0]),
    .S(_10814_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22642_ (.A(_10815_[0]),
    .B(_10816_[0]),
    .CI(_10817_[0]),
    .CO(_10818_[0]),
    .S(_10819_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22643_ (.A(_10820_[0]),
    .B(_10764_[0]),
    .CI(_10806_[0]),
    .CO(_10821_[0]),
    .S(_10822_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22644_ (.A(_10823_[0]),
    .B(_10780_[0]),
    .CI(_10822_[0]),
    .CO(_10824_[0]),
    .S(_10825_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22645_ (.A(net3229),
    .B(net3233),
    .CI(_10826_[0]),
    .CO(_10827_[0]),
    .S(_10828_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22646_ (.A(net3217),
    .B(_10786_[0]),
    .CI(_10828_[0]),
    .CO(_10829_[0]),
    .S(_10830_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22647_ (.A(net3202),
    .B(_10788_[0]),
    .CI(_10830_[0]),
    .CO(_10831_[0]),
    .S(_10832_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22648_ (.A(_10794_[0]),
    .B(_10833_[0]),
    .CI(_10834_[0]),
    .CO(_10835_[0]),
    .S(_10836_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22649_ (.A(_10758_[0]),
    .B(_10798_[0]),
    .CI(_10837_[0]),
    .CO(_10838_[0]),
    .S(_10839_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22650_ (.A(net3205),
    .B(_10799_[0]),
    .CI(_10839_[0]),
    .CO(_10840_[0]),
    .S(_10841_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22651_ (.A(_10841_[0]),
    .B(_10842_[0]),
    .CI(_10843_[0]),
    .CO(_10844_[0]),
    .S(_10845_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22652_ (.A(_10846_[0]),
    .B(_10847_[0]),
    .CI(_10848_[0]),
    .CO(_10849_[0]),
    .S(_10850_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22653_ (.A(_10810_[0]),
    .B(_10850_[0]),
    .CI(_10851_[0]),
    .CO(_10852_[0]),
    .S(_10853_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22654_ (.A(_10854_[0]),
    .B(_10855_[0]),
    .CI(_10856_[0]),
    .CO(_10857_[0]),
    .S(_10858_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22655_ (.A(_10859_[0]),
    .B(_10805_[0]),
    .CI(_10845_[0]),
    .CO(_10860_[0]),
    .S(_10861_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22656_ (.A(_10862_[0]),
    .B(_10821_[0]),
    .CI(_10861_[0]),
    .CO(_10863_[0]),
    .S(_10864_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22657_ (.A(net3229),
    .B(net3233),
    .CI(_10865_[0]),
    .CO(_10866_[0]),
    .S(_10867_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22658_ (.A(net3217),
    .B(_10827_[0]),
    .CI(_10867_[0]),
    .CO(_10868_[0]),
    .S(_10869_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22659_ (.A(net3202),
    .B(_10829_[0]),
    .CI(_10869_[0]),
    .CO(_10870_[0]),
    .S(_10871_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22660_ (.A(_10794_[0]),
    .B(_10834_[0]),
    .CI(_10872_[0]),
    .CO(_10873_[0]),
    .S(_10874_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22661_ (.A(_10758_[0]),
    .B(_10798_[0]),
    .CI(_10875_[0]),
    .CO(_10876_[0]),
    .S(_10877_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22662_ (.A(net3205),
    .B(_10838_[0]),
    .CI(_10877_[0]),
    .CO(_10878_[0]),
    .S(_10879_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22663_ (.A(_10879_[0]),
    .B(_10880_[0]),
    .CI(_10881_[0]),
    .CO(_10882_[0]),
    .S(_10883_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22664_ (.A(_10884_[0]),
    .B(_10885_[0]),
    .CI(_10886_[0]),
    .CO(_10887_[0]),
    .S(_10888_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22665_ (.A(_10849_[0]),
    .B(_10888_[0]),
    .CI(_10889_[0]),
    .CO(_10890_[0]),
    .S(_10891_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22666_ (.A(_10892_[0]),
    .B(_10893_[0]),
    .CI(_10894_[0]),
    .CO(_10895_[0]),
    .S(_10896_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22667_ (.A(_10897_[0]),
    .B(_10844_[0]),
    .CI(_10883_[0]),
    .CO(_10898_[0]),
    .S(_10899_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22668_ (.A(_10900_[0]),
    .B(_10860_[0]),
    .CI(_10899_[0]),
    .CO(_10901_[0]),
    .S(_10902_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22669_ (.A(net3229),
    .B(net3233),
    .CI(_10903_[0]),
    .CO(_10904_[0]),
    .S(_10905_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22670_ (.A(net3214),
    .B(_10906_[0]),
    .CI(_10907_[0]),
    .CO(_10908_[0]),
    .S(_10909_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22671_ (.A(_10910_[0]),
    .B(_10909_[0]),
    .CI(net3204),
    .CO(_10911_[0]),
    .S(_10912_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22672_ (.A(_10876_[0]),
    .B(net3205),
    .CI(_10877_[0]),
    .CO(_10913_[0]),
    .S(_10914_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22673_ (.A(_10915_[0]),
    .B(_10870_[0]),
    .CI(_10916_[0]),
    .CO(_10917_[0]),
    .S(_10918_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22674_ (.A(_10919_[0]),
    .B(_10920_[0]),
    .CI(_10921_[0]),
    .CO(_10922_[0]),
    .S(_10923_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22675_ (.A(_10887_[0]),
    .B(_10924_[0]),
    .CI(_10925_[0]),
    .CO(_10926_[0]),
    .S(_10927_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22676_ (.A(_10928_[0]),
    .B(_10929_[0]),
    .CI(_10930_[0]),
    .CO(_10931_[0]),
    .S(_10932_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22677_ (.A(_10933_[0]),
    .B(_10882_[0]),
    .CI(_10934_[0]),
    .CO(_10935_[0]),
    .S(_10936_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22678_ (.A(_10937_[0]),
    .B(_10898_[0]),
    .CI(_10936_[0]),
    .CO(_10938_[0]),
    .S(_10939_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22679_ (.A(_10940_[0]),
    .B(net3229),
    .CI(net3233),
    .CO(_10941_[0]),
    .S(_10942_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22680_ (.A(_10943_[0]),
    .B(_10944_[0]),
    .CI(net3214),
    .CO(_10945_[0]),
    .S(_10946_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22681_ (.A(_10908_[0]),
    .B(_10946_[0]),
    .CI(net3204),
    .CO(_10947_[0]),
    .S(_10948_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22682_ (.A(_10911_[0]),
    .B(_10948_[0]),
    .CI(_10914_[0]),
    .CO(_10949_[0]),
    .S(_10950_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22683_ (.A(_10951_[0]),
    .B(_10952_[0]),
    .CI(_10921_[0]),
    .CO(_10953_[0]),
    .S(_10954_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22684_ (.A(_10955_[0]),
    .B(_10956_[0]),
    .CI(_10925_[0]),
    .CO(_10957_[0]),
    .S(_10958_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22685_ (.A(_10959_[0]),
    .B(_10960_[0]),
    .CI(_10961_[0]),
    .CO(_10962_[0]),
    .S(_10963_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22686_ (.A(_10964_[0]),
    .B(_10965_[0]),
    .CI(_10950_[0]),
    .CO(_10966_[0]),
    .S(_10967_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22687_ (.A(_10968_[0]),
    .B(_10935_[0]),
    .CI(_10967_[0]),
    .CO(_10969_[0]),
    .S(_10970_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22688_ (.A(_10971_[0]),
    .B(net3229),
    .CI(net3233),
    .CO(_10972_[0]),
    .S(_10973_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22689_ (.A(_10974_[0]),
    .B(_10975_[0]),
    .CI(net3214),
    .CO(_10976_[0]),
    .S(_10977_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22690_ (.A(_10945_[0]),
    .B(_10977_[0]),
    .CI(net3204),
    .CO(_10978_[0]),
    .S(_10979_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22691_ (.A(_10947_[0]),
    .B(_10979_[0]),
    .CI(_10914_[0]),
    .CO(_10980_[0]),
    .S(_10981_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22692_ (.A(_10982_[0]),
    .B(_10952_[0]),
    .CI(_10921_[0]),
    .CO(_10983_[0]),
    .S(_10984_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22693_ (.A(_10953_[0]),
    .B(_10984_[0]),
    .CI(_10873_[0]),
    .CO(_10985_[0]),
    .S(_10986_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22694_ (.A(_10987_[0]),
    .B(_10988_[0]),
    .CI(_10961_[0]),
    .CO(_10989_[0]),
    .S(_10990_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22695_ (.A(_10991_[0]),
    .B(_10949_[0]),
    .CI(_10981_[0]),
    .CO(_10992_[0]),
    .S(_10993_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22696_ (.A(_10994_[0]),
    .B(_10966_[0]),
    .CI(_10993_[0]),
    .CO(_10995_[0]),
    .S(_10996_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addf_4 _22697_ (.A(_10997_[0]),
    .B(_10998_[0]),
    .CI(_10999_[0]),
    .CO(_11000_[0]),
    .S(_11001_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22698_ (.A(_11002_[0]),
    .B(net3286),
    .CO(_11004_[0]),
    .S(_11005_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22699_ (.A(_11002_[0]),
    .B(_11006_[0]),
    .CO(_11007_[0]),
    .S(_11008_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22700_ (.A(net463),
    .B(net3286),
    .CO(_11010_[0]),
    .S(_11011_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22701_ (.A(_11009_[0]),
    .B(_11006_[0]),
    .CO(_11012_[0]),
    .S(_11013_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22702_ (.A(net474),
    .B(_11015_[0]),
    .CO(_11016_[0]),
    .S(_11017_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22703_ (.A(_11018_[0]),
    .B(_11019_[0]),
    .CO(_11020_[0]),
    .S(_11021_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22704_ (.A(_11022_[0]),
    .B(_11023_[0]),
    .CO(_11024_[0]),
    .S(_11025_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22705_ (.A(_11027_[0]),
    .B(_11026_[0]),
    .CO(_11028_[0]),
    .S(_11029_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22706_ (.A(_11031_[0]),
    .B(_11030_[0]),
    .CO(_11032_[0]),
    .S(_11033_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22707_ (.A(_11035_[0]),
    .B(_11034_[0]),
    .CO(_11036_[0]),
    .S(_11037_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22708_ (.A(_11038_[0]),
    .B(_11039_[0]),
    .CO(_11040_[0]),
    .S(_11041_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22709_ (.A(_11043_[0]),
    .B(_11042_[0]),
    .CO(_11044_[0]),
    .S(_11045_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22710_ (.A(_11047_[0]),
    .B(_11046_[0]),
    .CO(_11048_[0]),
    .S(_11049_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22711_ (.A(_11051_[0]),
    .B(_11050_[0]),
    .CO(_11052_[0]),
    .S(_11053_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22712_ (.A(_11055_[0]),
    .B(_11054_[0]),
    .CO(_11056_[0]),
    .S(_11057_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22713_ (.A(_11058_[0]),
    .B(_11059_[0]),
    .CO(_11060_[0]),
    .S(_11061_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22714_ (.A(_11062_[0]),
    .B(_11063_[0]),
    .CO(_11064_[0]),
    .S(_11065_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22715_ (.A(_11066_[0]),
    .B(_11067_[0]),
    .CO(_11068_[0]),
    .S(_11069_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22716_ (.A(_11070_[0]),
    .B(_11071_[0]),
    .CO(_11072_[0]),
    .S(_11073_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22717_ (.A(_11075_[0]),
    .B(_11074_[0]),
    .CO(_11076_[0]),
    .S(_11077_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22718_ (.A(_11078_[0]),
    .B(_11079_[0]),
    .CO(_11080_[0]),
    .S(_11081_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22719_ (.A(_11082_[0]),
    .B(_11083_[0]),
    .CO(_11084_[0]),
    .S(_11085_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22720_ (.A(_11086_[0]),
    .B(_11087_[0]),
    .CO(_11088_[0]),
    .S(_11089_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22721_ (.A(_11090_[0]),
    .B(_11091_[0]),
    .CO(_11092_[0]),
    .S(_11093_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22722_ (.A(_11094_[0]),
    .B(_11095_[0]),
    .CO(_11096_[0]),
    .S(_11097_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22723_ (.A(_11099_[0]),
    .B(_11098_[0]),
    .CO(_11100_[0]),
    .S(_11101_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22724_ (.A(_11102_[0]),
    .B(_11103_[0]),
    .CO(_11104_[0]),
    .S(_11105_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22725_ (.A(_11106_[0]),
    .B(_11107_[0]),
    .CO(_11108_[0]),
    .S(_11109_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22726_ (.A(_11110_[0]),
    .B(_11111_[0]),
    .CO(_11112_[0]),
    .S(_11113_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22727_ (.A(_11114_[0]),
    .B(_11115_[0]),
    .CO(_11116_[0]),
    .S(_11117_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22728_ (.A(_11118_[0]),
    .B(_11119_[0]),
    .CO(_11120_[0]),
    .S(_11121_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22729_ (.A(_11122_[0]),
    .B(_11123_[0]),
    .CO(_11124_[0]),
    .S(_11125_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22730_ (.A(_11126_[0]),
    .B(_11127_[0]),
    .CO(_11128_[0]),
    .S(_11129_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22731_ (.A(_11130_[0]),
    .B(_11131_[0]),
    .CO(_11132_[0]),
    .S(_11133_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22732_ (.A(_11134_[0]),
    .B(_11135_[0]),
    .CO(_11136_[0]),
    .S(_11137_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22733_ (.A(_11138_[0]),
    .B(_11139_[0]),
    .CO(_11140_[0]),
    .S(_11141_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22734_ (.A(_11142_[0]),
    .B(_11143_[0]),
    .CO(_11144_[0]),
    .S(_11145_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22735_ (.A(_11146_[0]),
    .B(_11147_[0]),
    .CO(_11148_[0]),
    .S(_11149_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22736_ (.A(_11146_[0]),
    .B(_11150_[0]),
    .CO(_11151_[0]),
    .S(_11152_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22737_ (.A(_06849_),
    .B(_11147_[0]),
    .CO(_11154_[0]),
    .S(_11155_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22738_ (.A(_11156_[0]),
    .B(_11157_[0]),
    .CO(_11158_[0]),
    .S(_11159_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22739_ (.A(\cs_registers_i.priv_mode_id_o[0] ),
    .B(_11160_[0]),
    .CO(_11161_[0]),
    .S(_11162_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22740_ (.A(\cs_registers_i.mhpmcounter[1856] ),
    .B(\cs_registers_i.mhpmcounter[1857] ),
    .CO(_11163_[0]),
    .S(_11164_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22741_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .CO(_11165_[0]),
    .S(_11166_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22742_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .CO(_11167_[0]),
    .S(_11168_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22743_ (.A(_11169_[0]),
    .B(_11170_[0]),
    .CO(_11171_[0]),
    .S(_11172_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22744_ (.A(_11169_[0]),
    .B(_11170_[0]),
    .CO(_11173_[0]),
    .S(_11174_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22745_ (.A(_11169_[0]),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CO(_11175_[0]),
    .S(_11176_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22746_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_11170_[0]),
    .CO(_11177_[0]),
    .S(_11178_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22747_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CO(_11179_[0]),
    .S(_11180_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22748_ (.A(_11181_[0]),
    .B(_11182_[0]),
    .CO(_11183_[0]),
    .S(_11184_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22749_ (.A(_11183_[0]),
    .B(_11185_[0]),
    .CO(_11186_[0]),
    .S(_11187_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22750_ (.A(_11186_[0]),
    .B(_09763_[0]),
    .CO(_11188_[0]),
    .S(_11189_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22751_ (.A(_11190_[0]),
    .B(_11191_[0]),
    .CO(_09785_[0]),
    .S(_11192_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22752_ (.A(_09762_[0]),
    .B(_11193_[0]),
    .CO(_11194_[0]),
    .S(_11195_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22753_ (.A(_11188_[0]),
    .B(_11195_[0]),
    .CO(_11196_[0]),
    .S(_11197_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22754_ (.A(_11194_[0]),
    .B(_09789_[0]),
    .CO(_11198_[0]),
    .S(_11199_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22755_ (.A(_11196_[0]),
    .B(_11199_[0]),
    .CO(_11200_[0]),
    .S(_11201_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22756_ (.A(_11202_[0]),
    .B(_09780_[0]),
    .CO(_09821_[0]),
    .S(_11203_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22757_ (.A(_11204_[0]),
    .B(_09788_[0]),
    .CO(_11205_[0]),
    .S(_11206_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22758_ (.A(_11198_[0]),
    .B(_11206_[0]),
    .CO(_11207_[0]),
    .S(_11208_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22759_ (.A(_11200_[0]),
    .B(_11208_[0]),
    .CO(_11209_[0]),
    .S(_11210_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22760_ (.A(_11211_[0]),
    .B(_11212_[0]),
    .CO(_09844_[0]),
    .S(_11213_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22761_ (.A(_11213_[0]),
    .B(_11214_[0]),
    .CO(_09851_[0]),
    .S(_11215_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22762_ (.A(_11205_[0]),
    .B(_09825_[0]),
    .CO(_11216_[0]),
    .S(_11217_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22763_ (.A(_11207_[0]),
    .B(_11217_[0]),
    .CO(_11218_[0]),
    .S(_11219_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22764_ (.A(_11209_[0]),
    .B(_11219_[0]),
    .CO(_11220_[0]),
    .S(_11221_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22765_ (.A(_09824_[0]),
    .B(_09855_[0]),
    .CO(_11222_[0]),
    .S(_11223_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22766_ (.A(_11216_[0]),
    .B(_11223_[0]),
    .CO(_11224_[0]),
    .S(_11225_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22767_ (.A(_11218_[0]),
    .B(_11225_[0]),
    .CO(_11226_[0]),
    .S(_11227_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22768_ (.A(_11228_[0]),
    .B(_09846_[0]),
    .CO(_09917_[0]),
    .S(_11229_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22769_ (.A(_09854_[0]),
    .B(_11230_[0]),
    .CO(_11231_[0]),
    .S(_11232_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22770_ (.A(_11222_[0]),
    .B(_11232_[0]),
    .CO(_11233_[0]),
    .S(_11234_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22771_ (.A(_11224_[0]),
    .B(_11234_[0]),
    .CO(_11235_[0]),
    .S(_11236_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22772_ (.A(_11237_[0]),
    .B(_11238_[0]),
    .CO(_11239_[0]),
    .S(_11240_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22773_ (.A(_11240_[0]),
    .B(_09881_[0]),
    .CO(_09953_[0]),
    .S(_11241_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22774_ (.A(_11231_[0]),
    .B(_09921_[0]),
    .CO(_11242_[0]),
    .S(_11243_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22775_ (.A(_11233_[0]),
    .B(_11243_[0]),
    .CO(_11244_[0]),
    .S(_11245_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22776_ (.A(_11239_[0]),
    .B(_11246_[0]),
    .CO(_09991_[0]),
    .S(_11247_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22777_ (.A(_11247_[0]),
    .B(_09909_[0]),
    .CO(_09998_[0]),
    .S(_11248_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22778_ (.A(_09920_[0]),
    .B(_09957_[0]),
    .CO(_11249_[0]),
    .S(_11250_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22779_ (.A(_11242_[0]),
    .B(_11250_[0]),
    .CO(_11251_[0]),
    .S(_11252_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22780_ (.A(_09956_[0]),
    .B(_10002_[0]),
    .CO(_11253_[0]),
    .S(_11254_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22781_ (.A(_11249_[0]),
    .B(_11254_[0]),
    .CO(_11255_[0]),
    .S(_11256_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22782_ (.A(_11257_[0]),
    .B(_11258_[0]),
    .CO(_11259_[0]),
    .S(_11260_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22783_ (.A(_10001_[0]),
    .B(_11261_[0]),
    .CO(_11262_[0]),
    .S(_11263_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22784_ (.A(_11253_[0]),
    .B(_11263_[0]),
    .CO(_11264_[0]),
    .S(_11265_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22785_ (.A(_11259_[0]),
    .B(_11266_[0]),
    .CO(_10135_[0]),
    .S(_11267_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22786_ (.A(_11268_[0]),
    .B(_11269_[0]),
    .CO(_11270_[0]),
    .S(_11271_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22787_ (.A(_11262_[0]),
    .B(_11271_[0]),
    .CO(_11272_[0]),
    .S(_11273_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22788_ (.A(_11274_[0]),
    .B(_10073_[0]),
    .CO(_11275_[0]),
    .S(_11276_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22789_ (.A(_11276_[0]),
    .B(_10081_[0]),
    .CO(_10182_[0]),
    .S(_11277_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22790_ (.A(_10139_[0]),
    .B(_11270_[0]),
    .CO(_11278_[0]),
    .S(_11279_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22791_ (.A(_11280_[0]),
    .B(_11281_[0]),
    .CO(_10233_[0]),
    .S(_11282_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22792_ (.A(_11282_[0]),
    .B(_10119_[0]),
    .CO(_11283_[0]),
    .S(_11284_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22793_ (.A(_11275_[0]),
    .B(_11284_[0]),
    .CO(_10243_[0]),
    .S(_11285_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22794_ (.A(_11285_[0]),
    .B(_10127_[0]),
    .CO(_10250_[0]),
    .S(_11286_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22795_ (.A(_10138_[0]),
    .B(_10186_[0]),
    .CO(_11287_[0]),
    .S(_11288_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22796_ (.A(_10185_[0]),
    .B(_10254_[0]),
    .CO(_11289_[0]),
    .S(_11290_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22797_ (.A(_10235_[0]),
    .B(_11291_[0]),
    .CO(_10361_[0]),
    .S(_11292_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22798_ (.A(_10253_[0]),
    .B(_11293_[0]),
    .CO(_11294_[0]),
    .S(_11295_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22799_ (.A(_11296_[0]),
    .B(_11297_[0]),
    .CO(_10417_[0]),
    .S(_10362_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22800_ (.A(_11298_[0]),
    .B(_11299_[0]),
    .CO(_11300_[0]),
    .S(_11301_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22801_ (.A(_11302_[0]),
    .B(_11303_[0]),
    .CO(_10473_[0]),
    .S(_10418_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22802_ (.A(_11304_[0]),
    .B(_11305_[0]),
    .CO(_11306_[0]),
    .S(_11307_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22803_ (.A(_11308_[0]),
    .B(_11309_[0]),
    .CO(_10528_[0]),
    .S(_10474_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22804_ (.A(_11310_[0]),
    .B(_11311_[0]),
    .CO(_11312_[0]),
    .S(_11313_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22805_ (.A(_11314_[0]),
    .B(_11315_[0]),
    .CO(_10580_[0]),
    .S(_10529_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22806_ (.A(_11316_[0]),
    .B(_11317_[0]),
    .CO(_11318_[0]),
    .S(_11319_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22807_ (.A(_11320_[0]),
    .B(_11321_[0]),
    .CO(_10633_[0]),
    .S(_10581_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22808_ (.A(_11322_[0]),
    .B(_11323_[0]),
    .CO(_11324_[0]),
    .S(_11325_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22809_ (.A(_11326_[0]),
    .B(_11327_[0]),
    .CO(_10683_[0]),
    .S(_10634_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22810_ (.A(_11328_[0]),
    .B(_11329_[0]),
    .CO(_11330_[0]),
    .S(_11331_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22811_ (.A(_11332_[0]),
    .B(_11333_[0]),
    .CO(_10730_[0]),
    .S(_10684_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22812_ (.A(_11334_[0]),
    .B(_11335_[0]),
    .CO(_11336_[0]),
    .S(_11337_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22813_ (.A(_11338_[0]),
    .B(_11339_[0]),
    .CO(_10776_[0]),
    .S(_10731_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22814_ (.A(_11340_[0]),
    .B(_11341_[0]),
    .CO(_11342_[0]),
    .S(_11343_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22815_ (.A(_11344_[0]),
    .B(_11345_[0]),
    .CO(_10815_[0]),
    .S(_10774_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22816_ (.A(_11346_[0]),
    .B(_11347_[0]),
    .CO(_11348_[0]),
    .S(_11349_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22817_ (.A(_11350_[0]),
    .B(_11351_[0]),
    .CO(_10854_[0]),
    .S(_10816_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22818_ (.A(_11352_[0]),
    .B(_11353_[0]),
    .CO(_11354_[0]),
    .S(_11355_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22819_ (.A(_11356_[0]),
    .B(_11357_[0]),
    .CO(_10892_[0]),
    .S(_10855_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22820_ (.A(_11358_[0]),
    .B(_11359_[0]),
    .CO(_11360_[0]),
    .S(_11361_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22821_ (.A(_11362_[0]),
    .B(_11363_[0]),
    .CO(_10928_[0]),
    .S(_10893_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22822_ (.A(_11364_[0]),
    .B(_11365_[0]),
    .CO(_11366_[0]),
    .S(_11367_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22823_ (.A(_11368_[0]),
    .B(_11369_[0]),
    .CO(_10959_[0]),
    .S(_10929_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22824_ (.A(_11370_[0]),
    .B(_11371_[0]),
    .CO(_11372_[0]),
    .S(_11373_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22825_ (.A(_11374_[0]),
    .B(_11375_[0]),
    .CO(_10987_[0]),
    .S(_10960_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22826_ (.A(_11376_[0]),
    .B(_11377_[0]),
    .CO(_11378_[0]),
    .S(_11379_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22827_ (.A(_10984_[0]),
    .B(_10873_[0]),
    .CO(_11380_[0]),
    .S(_11381_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22828_ (.A(_11382_[0]),
    .B(_10986_[0]),
    .CO(_11383_[0]),
    .S(_10988_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22829_ (.A(_11384_[0]),
    .B(_11385_[0]),
    .CO(_11386_[0]),
    .S(_11387_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22830_ (.A(\cs_registers_i.pc_if_i[2] ),
    .B(_11388_[0]),
    .CO(_11389_[0]),
    .S(_11390_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22831_ (.A(net264),
    .B(net302),
    .CO(_11393_[0]),
    .S(_11394_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22832_ (.A(_11395_[0]),
    .B(_06388_),
    .CO(_11397_[0]),
    .S(_11398_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22833_ (.A(_11399_[0]),
    .B(net3253),
    .CO(_11400_[0]),
    .S(_11401_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22834_ (.A(_11402_[0]),
    .B(_06440_),
    .CO(_11404_[0]),
    .S(_11405_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22835_ (.A(_11406_[0]),
    .B(net264),
    .CO(_11407_[0]),
    .S(_11408_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22836_ (.A(_11409_[0]),
    .B(_11410_[0]),
    .CO(_11411_[0]),
    .S(_11412_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22837_ (.A(_11413_[0]),
    .B(_11414_[0]),
    .CO(_11415_[0]),
    .S(_11416_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22838_ (.A(_11417_[0]),
    .B(_11418_[0]),
    .CO(_11419_[0]),
    .S(_11420_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22839_ (.A(_11421_[0]),
    .B(net3288),
    .CO(_11423_[0]),
    .S(_11424_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22840_ (.A(net3252),
    .B(_06530_),
    .CO(_11427_[0]),
    .S(_11428_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22841_ (.A(_11429_[0]),
    .B(net3287),
    .CO(_11431_[0]),
    .S(_11432_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22842_ (.A(_11433_[0]),
    .B(_11434_[0]),
    .CO(_11435_[0]),
    .S(_11436_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22843_ (.A(_11437_[0]),
    .B(_11438_[0]),
    .CO(_11439_[0]),
    .S(_11440_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22844_ (.A(_11441_[0]),
    .B(_11442_[0]),
    .CO(_11443_[0]),
    .S(_11444_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22845_ (.A(_11445_[0]),
    .B(_11446_[0]),
    .CO(_11447_[0]),
    .S(_11448_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22846_ (.A(_11449_[0]),
    .B(_11450_[0]),
    .CO(_11451_[0]),
    .S(_11452_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22847_ (.A(_11453_[0]),
    .B(_11454_[0]),
    .CO(_11455_[0]),
    .S(_11456_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22848_ (.A(_11457_[0]),
    .B(_11458_[0]),
    .CO(_11459_[0]),
    .S(_11460_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22849_ (.A(_11461_[0]),
    .B(_11462_[0]),
    .CO(_11463_[0]),
    .S(_11464_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22850_ (.A(_11465_[0]),
    .B(_11466_[0]),
    .CO(_11467_[0]),
    .S(_11468_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22851_ (.A(_11469_[0]),
    .B(_11470_[0]),
    .CO(_11471_[0]),
    .S(_11472_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22852_ (.A(_11473_[0]),
    .B(_11474_[0]),
    .CO(_11475_[0]),
    .S(_11476_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22853_ (.A(_11477_[0]),
    .B(_11478_[0]),
    .CO(_11479_[0]),
    .S(_11480_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22854_ (.A(_11481_[0]),
    .B(_11482_[0]),
    .CO(_11483_[0]),
    .S(_11484_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22855_ (.A(_11485_[0]),
    .B(_11486_[0]),
    .CO(_11487_[0]),
    .S(_11488_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22856_ (.A(_11489_[0]),
    .B(_11490_[0]),
    .CO(_11491_[0]),
    .S(_11492_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22857_ (.A(_11493_[0]),
    .B(_11494_[0]),
    .CO(_11495_[0]),
    .S(_11496_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22858_ (.A(_11497_[0]),
    .B(_11498_[0]),
    .CO(_11499_[0]),
    .S(_11500_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22859_ (.A(_11501_[0]),
    .B(_11502_[0]),
    .CO(_11503_[0]),
    .S(_11504_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22860_ (.A(_11505_[0]),
    .B(_11506_[0]),
    .CO(_11507_[0]),
    .S(_11508_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22861_ (.A(_11509_[0]),
    .B(_11510_[0]),
    .CO(_11511_[0]),
    .S(_11512_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22862_ (.A(_11513_[0]),
    .B(_11514_[0]),
    .CO(_11515_[0]),
    .S(_11516_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22863_ (.A(_11517_[0]),
    .B(_11518_[0]),
    .CO(_11519_[0]),
    .S(_11520_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22864_ (.A(_11521_[0]),
    .B(_11522_[0]),
    .CO(_11523_[0]),
    .S(_11524_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22865_ (.A(_11525_[0]),
    .B(_11526_[0]),
    .CO(_11527_[0]),
    .S(_11528_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22866_ (.A(_11529_[0]),
    .B(_11530_[0]),
    .CO(_11531_[0]),
    .S(_11532_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22867_ (.A(_11533_[0]),
    .B(_11534_[0]),
    .CO(_11535_[0]),
    .S(_11536_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22868_ (.A(_11537_[0]),
    .B(_11538_[0]),
    .CO(_11539_[0]),
    .S(_11540_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22869_ (.A(_11541_[0]),
    .B(_11542_[0]),
    .CO(_11543_[0]),
    .S(_11544_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22870_ (.A(_11545_[0]),
    .B(_11546_[0]),
    .CO(_11547_[0]),
    .S(_11548_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22871_ (.A(_11549_[0]),
    .B(_11550_[0]),
    .CO(_11551_[0]),
    .S(_11552_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22872_ (.A(_11553_[0]),
    .B(_11554_[0]),
    .CO(_11555_[0]),
    .S(_11556_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22873_ (.A(_11557_[0]),
    .B(_11558_[0]),
    .CO(_11559_[0]),
    .S(_11560_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22874_ (.A(_11561_[0]),
    .B(_11562_[0]),
    .CO(_11563_[0]),
    .S(_11564_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22875_ (.A(_11565_[0]),
    .B(_11566_[0]),
    .CO(_11567_[0]),
    .S(_11568_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22876_ (.A(_11569_[0]),
    .B(_11570_[0]),
    .CO(_11571_[0]),
    .S(_11572_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22877_ (.A(_11573_[0]),
    .B(_11574_[0]),
    .CO(_11575_[0]),
    .S(_11576_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22878_ (.A(_11577_[0]),
    .B(_11578_[0]),
    .CO(_11579_[0]),
    .S(_11580_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22879_ (.A(_11581_[0]),
    .B(_11582_[0]),
    .CO(_11583_[0]),
    .S(_11584_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22880_ (.A(_11585_[0]),
    .B(_11586_[0]),
    .CO(_11587_[0]),
    .S(_11588_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22881_ (.A(_11589_[0]),
    .B(_11590_[0]),
    .CO(_11591_[0]),
    .S(_11592_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22882_ (.A(_11593_[0]),
    .B(_11594_[0]),
    .CO(_11595_[0]),
    .S(_11596_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22883_ (.A(_11597_[0]),
    .B(_11598_[0]),
    .CO(_11599_[0]),
    .S(_11600_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22884_ (.A(_11601_[0]),
    .B(_11602_[0]),
    .CO(_11603_[0]),
    .S(_11604_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22885_ (.A(_11605_[0]),
    .B(_11606_[0]),
    .CO(_11607_[0]),
    .S(_11608_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22886_ (.A(_11609_[0]),
    .B(_11610_[0]),
    .CO(_11611_[0]),
    .S(_11612_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22887_ (.A(_11613_[0]),
    .B(_11614_[0]),
    .CO(_11615_[0]),
    .S(_11616_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22888_ (.A(_11617_[0]),
    .B(_11618_[0]),
    .CO(_11619_[0]),
    .S(_11620_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22889_ (.A(_11621_[0]),
    .B(_11622_[0]),
    .CO(_11623_[0]),
    .S(_11624_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22890_ (.A(_11625_[0]),
    .B(_11626_[0]),
    .CO(_11627_[0]),
    .S(_11628_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22891_ (.A(_11629_[0]),
    .B(_11630_[0]),
    .CO(_11631_[0]),
    .S(_11632_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22892_ (.A(_11633_[0]),
    .B(_11634_[0]),
    .CO(_11635_[0]),
    .S(_11636_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22893_ (.A(_11637_[0]),
    .B(_11638_[0]),
    .CO(_11639_[0]),
    .S(_11640_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22894_ (.A(_11641_[0]),
    .B(_08425_),
    .CO(_11643_[0]),
    .S(_11644_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22895_ (.A(\alu_adder_result_ex[1] ),
    .B(\alu_adder_result_ex[0] ),
    .CO(_11645_[0]),
    .S(_11646_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22896_ (.A(\alu_adder_result_ex[1] ),
    .B(\alu_adder_result_ex[0] ),
    .CO(_11647_[0]),
    .S(_11648_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22897_ (.A(\alu_adder_result_ex[1] ),
    .B(_09748_[0]),
    .CO(_11649_[0]),
    .S(_11650_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22898_ (.A(\alu_adder_result_ex[1] ),
    .B(_09748_[0]),
    .CO(_11651_[0]),
    .S(_11652_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22899_ (.A(_11653_[0]),
    .B(\alu_adder_result_ex[0] ),
    .CO(_11654_[0]),
    .S(_11655_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22900_ (.A(_11653_[0]),
    .B(\alu_adder_result_ex[0] ),
    .CO(_11656_[0]),
    .S(_11657_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22901_ (.A(_11653_[0]),
    .B(_09748_[0]),
    .CO(_11658_[0]),
    .S(_11659_[0]));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22902_ (.A(_11660_[0]),
    .B(_11661_[0]),
    .CO(_11662_[0]),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22903_ (.A(_11663_[0]),
    .B(_11662_[0]),
    .CO(_11664_[0]),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22904_ (.D(_00007_),
    .RN(net148),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22905_ (.D(_00008_),
    .RN(net148),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22906_ (.D(_00009_),
    .RN(net3660),
    .CLK(clknet_leaf_382_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22907_ (.D(_00010_),
    .RN(net3660),
    .CLK(clknet_leaf_382_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 _22908_ (.D(_00011_),
    .SETN(net3660),
    .CLK(clknet_leaf_384_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22909_ (.D(_00012_),
    .RN(net3663),
    .CLK(clknet_leaf_475_clk),
    .Q(\load_store_unit_i.data_type_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22910_ (.D(_00013_),
    .RN(net3663),
    .CLK(clknet_leaf_476_clk),
    .Q(\load_store_unit_i.data_type_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_regs_0_core_clock (.I(clk_i),
    .Z(delaynet_0_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input31 (.I(data_rdata_i[13]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _22913_ (.I(net251),
    .Z(alert_minor_o));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _22914_ (.I(net252),
    .Z(data_addr_o[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _22915_ (.I(net253),
    .Z(data_addr_o[1]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input30 (.I(data_rdata_i[12]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input29 (.I(data_rdata_i[11]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input28 (.I(data_rdata_i[10]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input27 (.I(data_rdata_i[0]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 input26 (.I(data_gnt_i),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input25 (.I(data_err_i),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input24 (.I(boot_addr_i[9]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input23 (.I(boot_addr_i[8]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input22 (.I(boot_addr_i[31]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input21 (.I(boot_addr_i[30]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input20 (.I(boot_addr_i[29]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input19 (.I(boot_addr_i[28]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input18 (.I(boot_addr_i[27]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input17 (.I(boot_addr_i[26]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input16 (.I(boot_addr_i[25]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input15 (.I(boot_addr_i[24]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input14 (.I(boot_addr_i[23]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input13 (.I(boot_addr_i[22]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(boot_addr_i[21]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input11 (.I(boot_addr_i[20]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input10 (.I(boot_addr_i[19]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input9 (.I(boot_addr_i[18]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input8 (.I(boot_addr_i[17]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input7 (.I(boot_addr_i[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input6 (.I(boot_addr_i[15]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input5 (.I(boot_addr_i[14]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input4 (.I(boot_addr_i[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input3 (.I(boot_addr_i[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input2 (.I(boot_addr_i[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(boot_addr_i[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _22946_ (.I(net254),
    .Z(instr_addr_o[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlya_4 _22947_ (.I(net255),
    .Z(instr_addr_o[1]));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \core_busy_q$_DFF_PN0_  (.D(core_busy_d),
    .RN(net148),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(core_busy_q));
 gf180mcu_fd_sc_mcu9t5v0__latsnq_2 \core_clock_gate_i.en_latch$_DLATCH_N_  (.D(_00006_),
    .E(clknet_leaf_8_clk_i_regs),
    .Q(\core_clock_gate_i.en_latch ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.D(_00014_),
    .RN(net148),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.mcountinhibit_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.D(_00015_),
    .RN(net148),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mcountinhibit_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.D(_00016_),
    .RN(net148),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.D(_00017_),
    .RN(net148),
    .CLK(clknet_leaf_129_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.D(_00018_),
    .RN(net148),
    .CLK(clknet_leaf_128_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.D(_00019_),
    .RN(net148),
    .CLK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.D(_00020_),
    .RN(net148),
    .CLK(clknet_leaf_130_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.D(_00021_),
    .RN(net148),
    .CLK(clknet_leaf_135_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.D(_00022_),
    .RN(net148),
    .CLK(clknet_leaf_135_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.D(_00023_),
    .RN(net148),
    .CLK(clknet_leaf_140_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.D(_00024_),
    .RN(net148),
    .CLK(clknet_leaf_140_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.D(_00025_),
    .RN(net148),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.D(_00026_),
    .RN(net148),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.D(_00027_),
    .RN(net148),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.D(_00028_),
    .RN(net148),
    .CLK(clknet_leaf_168_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.D(_00029_),
    .RN(net148),
    .CLK(clknet_leaf_168_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.D(_00030_),
    .RN(net148),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.D(_00031_),
    .RN(net148),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.D(_00032_),
    .RN(net148),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.D(_00033_),
    .RN(net148),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.D(_00034_),
    .RN(net148),
    .CLK(clknet_leaf_173_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.D(_00035_),
    .RN(net148),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.D(_00036_),
    .RN(net148),
    .CLK(clknet_leaf_173_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.D(_00037_),
    .RN(net148),
    .CLK(clknet_leaf_175_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.D(_00038_),
    .RN(net148),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.D(_00039_),
    .RN(net148),
    .CLK(clknet_leaf_173_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.D(_00040_),
    .RN(net148),
    .CLK(clknet_leaf_175_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.D(_00041_),
    .RN(net148),
    .CLK(clknet_leaf_129_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.D(_00042_),
    .RN(net148),
    .CLK(clknet_leaf_612_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.D(_00043_),
    .RN(net148),
    .CLK(clknet_leaf_612_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.D(_00044_),
    .RN(net148),
    .CLK(clknet_leaf_612_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.D(_00045_),
    .RN(net148),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.D(_00046_),
    .RN(net148),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.D(_00047_),
    .RN(net148),
    .CLK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.D(_00048_),
    .RN(net148),
    .CLK(clknet_leaf_128_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.D(_00049_),
    .RN(net148),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.D(_00050_),
    .RN(net148),
    .CLK(clknet_leaf_117_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.D(_00051_),
    .RN(net148),
    .CLK(clknet_leaf_117_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.D(_00052_),
    .RN(net148),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.D(_00053_),
    .RN(net148),
    .CLK(clknet_6_32__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.D(_00054_),
    .RN(net148),
    .CLK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.D(_00055_),
    .RN(net148),
    .CLK(clknet_leaf_132_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.D(_00056_),
    .RN(net148),
    .CLK(clknet_6_32__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.D(_00057_),
    .RN(net148),
    .CLK(clknet_leaf_146_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.D(_00058_),
    .RN(net148),
    .CLK(clknet_leaf_149_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.D(_00059_),
    .RN(net148),
    .CLK(clknet_leaf_139_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.D(_00060_),
    .RN(net148),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.D(_00061_),
    .RN(net148),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.D(_00062_),
    .RN(net148),
    .CLK(clknet_leaf_138_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.D(_00063_),
    .RN(net148),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.D(_00064_),
    .RN(net148),
    .CLK(clknet_leaf_139_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.D(_00065_),
    .RN(net148),
    .CLK(clknet_leaf_181_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.D(_00066_),
    .RN(net148),
    .CLK(clknet_leaf_181_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.D(_00067_),
    .RN(net148),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.D(_00068_),
    .RN(net148),
    .CLK(clknet_leaf_178_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.D(_00069_),
    .RN(net148),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.D(_00070_),
    .RN(net148),
    .CLK(clknet_leaf_178_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.D(_00071_),
    .RN(net148),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.D(_00072_),
    .RN(net148),
    .CLK(clknet_leaf_174_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.D(_00073_),
    .RN(net148),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.D(_00074_),
    .RN(net148),
    .CLK(clknet_leaf_174_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.D(_00075_),
    .RN(net148),
    .CLK(clknet_leaf_175_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.D(_00076_),
    .RN(net148),
    .CLK(clknet_leaf_125_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.D(_00077_),
    .RN(net148),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.D(_00078_),
    .RN(net148),
    .CLK(clknet_leaf_127_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.D(_00079_),
    .RN(net148),
    .CLK(clknet_leaf_127_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.D(_00080_),
    .RN(net148),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1856] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.D(_00081_),
    .RN(net148),
    .CLK(clknet_leaf_131_clk),
    .Q(\cs_registers_i.mhpmcounter[1866] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.D(_00082_),
    .RN(net148),
    .CLK(clknet_leaf_131_clk),
    .Q(\cs_registers_i.mhpmcounter[1867] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.D(_00083_),
    .RN(net148),
    .CLK(clknet_6_32__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1868] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.D(_00084_),
    .RN(net148),
    .CLK(clknet_6_32__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1869] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.D(_00085_),
    .RN(net148),
    .CLK(clknet_leaf_146_clk),
    .Q(\cs_registers_i.mhpmcounter[1870] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.D(_00086_),
    .RN(net148),
    .CLK(clknet_6_32__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1871] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.D(_00087_),
    .RN(net148),
    .CLK(clknet_leaf_138_clk),
    .Q(\cs_registers_i.mhpmcounter[1872] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.D(_00088_),
    .RN(net148),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1873] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.D(_00089_),
    .RN(net148),
    .CLK(clknet_leaf_143_clk),
    .Q(\cs_registers_i.mhpmcounter[1874] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.D(_00090_),
    .RN(net148),
    .CLK(clknet_leaf_143_clk),
    .Q(\cs_registers_i.mhpmcounter[1875] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.D(_00091_),
    .RN(net148),
    .CLK(clknet_leaf_611_clk),
    .Q(\cs_registers_i.mhpmcounter[1857] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.D(_00092_),
    .RN(net148),
    .CLK(clknet_6_34__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1876] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.D(_00093_),
    .RN(net148),
    .CLK(clknet_leaf_167_clk),
    .Q(\cs_registers_i.mhpmcounter[1877] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.D(_00094_),
    .RN(net148),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1878] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.D(_00095_),
    .RN(net148),
    .CLK(clknet_leaf_167_clk),
    .Q(\cs_registers_i.mhpmcounter[1879] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.D(_00096_),
    .RN(net148),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1880] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.D(_00097_),
    .RN(net148),
    .CLK(clknet_leaf_165_clk),
    .Q(\cs_registers_i.mhpmcounter[1881] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.D(_00098_),
    .RN(net148),
    .CLK(clknet_leaf_165_clk),
    .Q(\cs_registers_i.mhpmcounter[1882] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.D(_00099_),
    .RN(net148),
    .CLK(clknet_leaf_160_clk),
    .Q(\cs_registers_i.mhpmcounter[1883] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.D(_00100_),
    .RN(net148),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1884] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.D(_00101_),
    .RN(net148),
    .CLK(clknet_6_40__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1885] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.D(_00102_),
    .RN(net148),
    .CLK(clknet_leaf_611_clk),
    .Q(\cs_registers_i.mhpmcounter[1858] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.D(_00103_),
    .RN(net148),
    .CLK(clknet_leaf_162_clk),
    .Q(\cs_registers_i.mhpmcounter[1886] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.D(_00104_),
    .RN(net148),
    .CLK(clknet_leaf_162_clk),
    .Q(\cs_registers_i.mhpmcounter[1887] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.D(_00105_),
    .RN(net148),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1888] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.D(_00106_),
    .RN(net148),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1889] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.D(_00107_),
    .RN(net148),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mhpmcounter[1890] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.D(_00108_),
    .RN(net148),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1891] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.D(_00109_),
    .RN(net148),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1892] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.D(_00110_),
    .RN(net148),
    .CLK(clknet_6_14__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1893] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.D(_00111_),
    .RN(net148),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1894] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.D(_00112_),
    .RN(net148),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1895] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.D(_00113_),
    .RN(net148),
    .CLK(clknet_6_8__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1859] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.D(_00114_),
    .RN(net148),
    .CLK(clknet_6_14__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1896] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.D(_00115_),
    .RN(net148),
    .CLK(clknet_6_14__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1897] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.D(_00116_),
    .RN(net148),
    .CLK(clknet_6_14__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1898] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.D(_00117_),
    .RN(net148),
    .CLK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.mhpmcounter[1899] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.D(_00118_),
    .RN(net148),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1900] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.D(_00119_),
    .RN(net148),
    .CLK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[1901] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.D(_00120_),
    .RN(net148),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1902] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.D(_00121_),
    .RN(net148),
    .CLK(clknet_leaf_98_clk),
    .Q(\cs_registers_i.mhpmcounter[1903] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.D(_00122_),
    .RN(net148),
    .CLK(clknet_leaf_157_clk),
    .Q(\cs_registers_i.mhpmcounter[1904] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.D(_00123_),
    .RN(net148),
    .CLK(clknet_leaf_149_clk),
    .Q(\cs_registers_i.mhpmcounter[1905] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.D(_00124_),
    .RN(net148),
    .CLK(clknet_leaf_620_clk),
    .Q(\cs_registers_i.mhpmcounter[1860] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.D(_00125_),
    .RN(net148),
    .CLK(clknet_leaf_151_clk),
    .Q(\cs_registers_i.mhpmcounter[1906] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.D(_00126_),
    .RN(net148),
    .CLK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.mhpmcounter[1907] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.D(_00127_),
    .RN(net148),
    .CLK(clknet_leaf_150_clk),
    .Q(\cs_registers_i.mhpmcounter[1908] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.D(_00128_),
    .RN(net148),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1909] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.D(_00129_),
    .RN(net148),
    .CLK(clknet_leaf_183_clk),
    .Q(\cs_registers_i.mhpmcounter[1910] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.D(_00130_),
    .RN(net148),
    .CLK(clknet_leaf_183_clk),
    .Q(\cs_registers_i.mhpmcounter[1911] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.D(_00131_),
    .RN(net148),
    .CLK(clknet_leaf_183_clk),
    .Q(\cs_registers_i.mhpmcounter[1912] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.D(_00132_),
    .RN(net148),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1913] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.D(_00133_),
    .RN(net148),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1914] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.D(_00134_),
    .RN(net148),
    .CLK(clknet_leaf_186_clk),
    .Q(\cs_registers_i.mhpmcounter[1915] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.D(_00135_),
    .RN(net148),
    .CLK(clknet_leaf_620_clk),
    .Q(\cs_registers_i.mhpmcounter[1861] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.D(_00136_),
    .RN(net148),
    .CLK(clknet_leaf_186_clk),
    .Q(\cs_registers_i.mhpmcounter[1916] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.D(_00137_),
    .RN(net148),
    .CLK(clknet_leaf_197_clk),
    .Q(\cs_registers_i.mhpmcounter[1917] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.D(_00138_),
    .RN(net148),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1918] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.D(_00139_),
    .RN(net148),
    .CLK(clknet_6_42__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1919] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.D(_00140_),
    .RN(net148),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1862] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.D(_00141_),
    .RN(net148),
    .CLK(clknet_6_10__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1863] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.D(_00142_),
    .RN(net148),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1864] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.D(_00143_),
    .RN(net148),
    .CLK(clknet_6_11__leaf_clk),
    .Q(\cs_registers_i.mhpmcounter[1865] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \cs_registers_i.priv_mode_id_o[0]$_DFFE_PN1P_  (.D(_00144_),
    .SETN(net3661),
    .CLK(clknet_leaf_29_clk),
    .Q(\cs_registers_i.priv_mode_id_o[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \cs_registers_i.priv_mode_id_o[1]$_DFFE_PN1P_  (.D(_00145_),
    .SETN(net3661),
    .CLK(clknet_leaf_29_clk),
    .Q(\cs_registers_i.priv_mode_id_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \cs_registers_i.u_dcsr_csr.rd_data_o[0]$_DFFE_PN1P_  (.D(_00146_),
    .SETN(net3661),
    .CLK(clknet_leaf_34_clk),
    .Q(\cs_registers_i.dcsr_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00147_),
    .RN(net3660),
    .CLK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.dcsr_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00148_),
    .RN(net3660),
    .CLK(clknet_6_15__leaf_clk),
    .Q(\cs_registers_i.dcsr_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00149_),
    .RN(net3660),
    .CLK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.dcsr_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00150_),
    .RN(net3660),
    .CLK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.dcsr_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \cs_registers_i.u_dcsr_csr.rd_data_o[1]$_DFFE_PN1P_  (.D(_00151_),
    .SETN(net3661),
    .CLK(clknet_leaf_34_clk),
    .Q(\cs_registers_i.dcsr_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00152_),
    .RN(net148),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.dcsr_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00153_),
    .RN(net3661),
    .CLK(clknet_leaf_32_clk),
    .Q(\cs_registers_i.dcsr_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00154_),
    .RN(net3661),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\cs_registers_i.dcsr_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00155_),
    .RN(net3661),
    .CLK(clknet_leaf_32_clk),
    .Q(\cs_registers_i.dcsr_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00156_),
    .RN(net148),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00157_),
    .RN(net3660),
    .CLK(clknet_6_15__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00158_),
    .RN(net3660),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00159_),
    .RN(net3660),
    .CLK(clknet_leaf_298_clk),
    .Q(\cs_registers_i.csr_depc_o[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00160_),
    .RN(net3660),
    .CLK(clknet_leaf_258_clk),
    .Q(\cs_registers_i.csr_depc_o[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00161_),
    .RN(net148),
    .CLK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.csr_depc_o[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00162_),
    .RN(net3660),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00163_),
    .RN(net3660),
    .CLK(clknet_leaf_272_clk),
    .Q(\cs_registers_i.csr_depc_o[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00164_),
    .RN(net3660),
    .CLK(clknet_leaf_192_clk),
    .Q(\cs_registers_i.csr_depc_o[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00165_),
    .RN(net3660),
    .CLK(clknet_leaf_286_clk),
    .Q(\cs_registers_i.csr_depc_o[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00166_),
    .RN(net148),
    .CLK(clknet_leaf_37_clk),
    .Q(\cs_registers_i.csr_depc_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00167_),
    .RN(net148),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00168_),
    .RN(net3660),
    .CLK(clknet_leaf_275_clk),
    .Q(\cs_registers_i.csr_depc_o[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00169_),
    .RN(net3660),
    .CLK(clknet_leaf_215_clk),
    .Q(\cs_registers_i.csr_depc_o[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00170_),
    .RN(net3660),
    .CLK(clknet_leaf_233_clk),
    .Q(\cs_registers_i.csr_depc_o[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00171_),
    .RN(net3660),
    .CLK(clknet_leaf_220_clk),
    .Q(\cs_registers_i.csr_depc_o[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00172_),
    .RN(net3660),
    .CLK(clknet_leaf_215_clk),
    .Q(\cs_registers_i.csr_depc_o[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00173_),
    .RN(net3660),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00174_),
    .RN(net3660),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00175_),
    .RN(net3660),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00176_),
    .RN(net3660),
    .CLK(clknet_leaf_214_clk),
    .Q(\cs_registers_i.csr_depc_o[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00177_),
    .RN(net3661),
    .CLK(clknet_leaf_33_clk),
    .Q(\cs_registers_i.csr_depc_o[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00178_),
    .RN(net3660),
    .CLK(clknet_leaf_296_clk),
    .Q(\cs_registers_i.csr_depc_o[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00179_),
    .RN(net148),
    .CLK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.csr_depc_o[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00180_),
    .RN(net148),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00181_),
    .RN(net3660),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00182_),
    .RN(net3660),
    .CLK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_depc_o[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00183_),
    .RN(net148),
    .CLK(clknet_leaf_54_clk),
    .Q(\cs_registers_i.csr_depc_o[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00184_),
    .RN(net148),
    .CLK(clknet_6_26__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00185_),
    .RN(net3660),
    .CLK(clknet_6_26__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00186_),
    .RN(net3660),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.csr_depc_o[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00187_),
    .RN(net148),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\cs_registers_i.dscratch0_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00188_),
    .RN(net148),
    .CLK(clknet_leaf_57_clk),
    .Q(\cs_registers_i.dscratch0_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00189_),
    .RN(net148),
    .CLK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.dscratch0_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00190_),
    .RN(net148),
    .CLK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.dscratch0_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00191_),
    .RN(net3660),
    .CLK(clknet_leaf_74_clk),
    .Q(\cs_registers_i.dscratch0_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00192_),
    .RN(net3660),
    .CLK(clknet_leaf_265_clk),
    .Q(\cs_registers_i.dscratch0_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00193_),
    .RN(net148),
    .CLK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.dscratch0_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00194_),
    .RN(net3660),
    .CLK(clknet_leaf_269_clk),
    .Q(\cs_registers_i.dscratch0_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00195_),
    .RN(net3660),
    .CLK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.dscratch0_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00196_),
    .RN(net148),
    .CLK(clknet_leaf_157_clk),
    .Q(\cs_registers_i.dscratch0_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00197_),
    .RN(net3660),
    .CLK(clknet_leaf_284_clk),
    .Q(\cs_registers_i.dscratch0_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00198_),
    .RN(net148),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\cs_registers_i.dscratch0_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00199_),
    .RN(net148),
    .CLK(clknet_leaf_152_clk),
    .Q(\cs_registers_i.dscratch0_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00200_),
    .RN(net3660),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\cs_registers_i.dscratch0_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00201_),
    .RN(net3660),
    .CLK(clknet_leaf_206_clk),
    .Q(\cs_registers_i.dscratch0_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00202_),
    .RN(net3660),
    .CLK(clknet_leaf_264_clk),
    .Q(\cs_registers_i.dscratch0_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00203_),
    .RN(net148),
    .CLK(clknet_leaf_161_clk),
    .Q(\cs_registers_i.dscratch0_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00204_),
    .RN(net148),
    .CLK(clknet_leaf_156_clk),
    .Q(\cs_registers_i.dscratch0_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00205_),
    .RN(net148),
    .CLK(clknet_leaf_160_clk),
    .Q(\cs_registers_i.dscratch0_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00206_),
    .RN(net148),
    .CLK(clknet_leaf_160_clk),
    .Q(\cs_registers_i.dscratch0_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00207_),
    .RN(net148),
    .CLK(clknet_leaf_156_clk),
    .Q(\cs_registers_i.dscratch0_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00208_),
    .RN(net148),
    .CLK(clknet_leaf_156_clk),
    .Q(\cs_registers_i.dscratch0_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00209_),
    .RN(net148),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\cs_registers_i.dscratch0_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00210_),
    .RN(net3660),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\cs_registers_i.dscratch0_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00211_),
    .RN(net148),
    .CLK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.dscratch0_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00212_),
    .RN(net148),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.dscratch0_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00213_),
    .RN(net148),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.dscratch0_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00214_),
    .RN(net3660),
    .CLK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.dscratch0_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00215_),
    .RN(net148),
    .CLK(clknet_leaf_44_clk),
    .Q(\cs_registers_i.dscratch0_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00216_),
    .RN(net148),
    .CLK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.dscratch0_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00217_),
    .RN(net148),
    .CLK(clknet_leaf_56_clk),
    .Q(\cs_registers_i.dscratch0_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00218_),
    .RN(net3660),
    .CLK(clknet_leaf_277_clk),
    .Q(\cs_registers_i.dscratch0_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00219_),
    .RN(net148),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00220_),
    .RN(net148),
    .CLK(clknet_leaf_57_clk),
    .Q(\cs_registers_i.dscratch1_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00221_),
    .RN(net3660),
    .CLK(clknet_6_15__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00222_),
    .RN(net3660),
    .CLK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.dscratch1_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00223_),
    .RN(net3660),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00224_),
    .RN(net3660),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00225_),
    .RN(net148),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00226_),
    .RN(net3660),
    .CLK(clknet_leaf_207_clk),
    .Q(\cs_registers_i.dscratch1_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00227_),
    .RN(net3660),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00228_),
    .RN(net148),
    .CLK(clknet_leaf_199_clk),
    .Q(\cs_registers_i.dscratch1_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00229_),
    .RN(net3660),
    .CLK(clknet_leaf_284_clk),
    .Q(\cs_registers_i.dscratch1_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00230_),
    .RN(net148),
    .CLK(clknet_leaf_37_clk),
    .Q(\cs_registers_i.dscratch1_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00231_),
    .RN(net148),
    .CLK(clknet_leaf_151_clk),
    .Q(\cs_registers_i.dscratch1_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00232_),
    .RN(net3660),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00233_),
    .RN(net3660),
    .CLK(clknet_leaf_213_clk),
    .Q(\cs_registers_i.dscratch1_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00234_),
    .RN(net3660),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00235_),
    .RN(net148),
    .CLK(clknet_leaf_198_clk),
    .Q(\cs_registers_i.dscratch1_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00236_),
    .RN(net3660),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00237_),
    .RN(net148),
    .CLK(clknet_leaf_198_clk),
    .Q(\cs_registers_i.dscratch1_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00238_),
    .RN(net148),
    .CLK(clknet_leaf_192_clk),
    .Q(\cs_registers_i.dscratch1_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00239_),
    .RN(net3660),
    .CLK(clknet_leaf_202_clk),
    .Q(\cs_registers_i.dscratch1_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00240_),
    .RN(net3660),
    .CLK(clknet_leaf_214_clk),
    .Q(\cs_registers_i.dscratch1_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00241_),
    .RN(net3661),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00242_),
    .RN(net3660),
    .CLK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.dscratch1_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00243_),
    .RN(net148),
    .CLK(clknet_leaf_100_clk),
    .Q(\cs_registers_i.dscratch1_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00244_),
    .RN(net3660),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00245_),
    .RN(net148),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00246_),
    .RN(net3660),
    .CLK(clknet_6_15__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00247_),
    .RN(net148),
    .CLK(clknet_leaf_44_clk),
    .Q(\cs_registers_i.dscratch1_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00248_),
    .RN(net148),
    .CLK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.dscratch1_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00249_),
    .RN(net148),
    .CLK(clknet_leaf_56_clk),
    .Q(\cs_registers_i.dscratch1_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00250_),
    .RN(net3660),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\cs_registers_i.dscratch1_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00251_),
    .RN(net148),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.mcause_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00252_),
    .RN(net148),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcause_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00253_),
    .RN(net148),
    .CLK(clknet_leaf_42_clk),
    .Q(\cs_registers_i.mcause_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00254_),
    .RN(net148),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcause_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00255_),
    .RN(net148),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\cs_registers_i.mcause_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00256_),
    .RN(net148),
    .CLK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mcause_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00257_),
    .RN(net148),
    .CLK(clknet_leaf_610_clk),
    .Q(\cs_registers_i.csr_mepc_o[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00258_),
    .RN(net148),
    .CLK(clknet_leaf_298_clk),
    .Q(\cs_registers_i.csr_mepc_o[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00259_),
    .RN(net3660),
    .CLK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.csr_mepc_o[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00260_),
    .RN(net3660),
    .CLK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.csr_mepc_o[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00261_),
    .RN(net3660),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00262_),
    .RN(net3660),
    .CLK(clknet_leaf_258_clk),
    .Q(\cs_registers_i.csr_mepc_o[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00263_),
    .RN(net148),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00264_),
    .RN(net3660),
    .CLK(clknet_leaf_209_clk),
    .Q(\cs_registers_i.csr_mepc_o[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00265_),
    .RN(net3660),
    .CLK(clknet_leaf_266_clk),
    .Q(\cs_registers_i.csr_mepc_o[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00266_),
    .RN(net3660),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00267_),
    .RN(net3660),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00268_),
    .RN(net148),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.csr_mepc_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00269_),
    .RN(net148),
    .CLK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.csr_mepc_o[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00270_),
    .RN(net3660),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00271_),
    .RN(net3660),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00272_),
    .RN(net3660),
    .CLK(clknet_leaf_233_clk),
    .Q(\cs_registers_i.csr_mepc_o[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00273_),
    .RN(net3660),
    .CLK(clknet_leaf_188_clk),
    .Q(\cs_registers_i.csr_mepc_o[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00274_),
    .RN(net3660),
    .CLK(clknet_leaf_229_clk),
    .Q(\cs_registers_i.csr_mepc_o[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00275_),
    .RN(net3660),
    .CLK(clknet_leaf_188_clk),
    .Q(\cs_registers_i.csr_mepc_o[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00276_),
    .RN(net3660),
    .CLK(clknet_leaf_195_clk),
    .Q(\cs_registers_i.csr_mepc_o[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00277_),
    .RN(net3660),
    .CLK(clknet_leaf_220_clk),
    .Q(\cs_registers_i.csr_mepc_o[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00278_),
    .RN(net3660),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00279_),
    .RN(net148),
    .CLK(clknet_leaf_38_clk),
    .Q(\cs_registers_i.csr_mepc_o[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00280_),
    .RN(net3660),
    .CLK(clknet_leaf_281_clk),
    .Q(\cs_registers_i.csr_mepc_o[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00281_),
    .RN(net148),
    .CLK(clknet_6_14__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00282_),
    .RN(net148),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00283_),
    .RN(net148),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\cs_registers_i.csr_mepc_o[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00284_),
    .RN(net3660),
    .CLK(clknet_leaf_64_clk),
    .Q(\cs_registers_i.csr_mepc_o[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00285_),
    .RN(net148),
    .CLK(clknet_leaf_54_clk),
    .Q(\cs_registers_i.csr_mepc_o[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00286_),
    .RN(net148),
    .CLK(clknet_leaf_53_clk),
    .Q(\cs_registers_i.csr_mepc_o[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00287_),
    .RN(net3660),
    .CLK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.csr_mepc_o[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00288_),
    .RN(net3660),
    .CLK(clknet_leaf_281_clk),
    .Q(\cs_registers_i.csr_mepc_o[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00289_),
    .RN(net3660),
    .CLK(clknet_leaf_269_clk),
    .Q(\cs_registers_i.mie_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00290_),
    .RN(net148),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\cs_registers_i.mie_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00291_),
    .RN(net148),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\cs_registers_i.mie_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00292_),
    .RN(net148),
    .CLK(clknet_leaf_155_clk),
    .Q(\cs_registers_i.mie_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00293_),
    .RN(net148),
    .CLK(clknet_leaf_155_clk),
    .Q(\cs_registers_i.mie_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00294_),
    .RN(net3660),
    .CLK(clknet_leaf_78_clk),
    .Q(\cs_registers_i.mie_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00295_),
    .RN(net148),
    .CLK(clknet_6_14__leaf_clk),
    .Q(\cs_registers_i.mie_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00296_),
    .RN(net148),
    .CLK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.mie_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00297_),
    .RN(net148),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.mie_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00298_),
    .RN(net3660),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\cs_registers_i.mie_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00299_),
    .RN(net148),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\cs_registers_i.mie_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00300_),
    .RN(net3660),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\cs_registers_i.mie_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00301_),
    .RN(net148),
    .CLK(clknet_leaf_150_clk),
    .Q(\cs_registers_i.mie_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00302_),
    .RN(net3660),
    .CLK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mie_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00303_),
    .RN(net3660),
    .CLK(clknet_leaf_211_clk),
    .Q(\cs_registers_i.mie_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00304_),
    .RN(net3660),
    .CLK(clknet_leaf_264_clk),
    .Q(\cs_registers_i.mie_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00305_),
    .RN(net148),
    .CLK(clknet_leaf_161_clk),
    .Q(\cs_registers_i.mie_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00306_),
    .RN(net3660),
    .CLK(clknet_leaf_206_clk),
    .Q(\cs_registers_i.mie_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00307_),
    .RN(net148),
    .CLK(clknet_6_12__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00308_),
    .RN(net148),
    .CLK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.mscratch_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00309_),
    .RN(net148),
    .CLK(clknet_leaf_107_clk),
    .Q(\cs_registers_i.mscratch_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00310_),
    .RN(net148),
    .CLK(clknet_leaf_102_clk),
    .Q(\cs_registers_i.mscratch_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00311_),
    .RN(net3660),
    .CLK(clknet_6_15__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00312_),
    .RN(net3660),
    .CLK(clknet_leaf_265_clk),
    .Q(\cs_registers_i.mscratch_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00313_),
    .RN(net148),
    .CLK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mscratch_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00314_),
    .RN(net3660),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00315_),
    .RN(net3660),
    .CLK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mscratch_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00316_),
    .RN(net148),
    .CLK(clknet_leaf_199_clk),
    .Q(\cs_registers_i.mscratch_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00317_),
    .RN(net3660),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00318_),
    .RN(net148),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00319_),
    .RN(net148),
    .CLK(clknet_leaf_152_clk),
    .Q(\cs_registers_i.mscratch_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00320_),
    .RN(net3660),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00321_),
    .RN(net3660),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00322_),
    .RN(net3660),
    .CLK(clknet_leaf_264_clk),
    .Q(\cs_registers_i.mscratch_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00323_),
    .RN(net148),
    .CLK(clknet_leaf_198_clk),
    .Q(\cs_registers_i.mscratch_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00324_),
    .RN(net3660),
    .CLK(clknet_leaf_211_clk),
    .Q(\cs_registers_i.mscratch_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00325_),
    .RN(net148),
    .CLK(clknet_leaf_198_clk),
    .Q(\cs_registers_i.mscratch_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00326_),
    .RN(net148),
    .CLK(clknet_leaf_197_clk),
    .Q(\cs_registers_i.mscratch_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00327_),
    .RN(net3660),
    .CLK(clknet_leaf_202_clk),
    .Q(\cs_registers_i.mscratch_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00328_),
    .RN(net3660),
    .CLK(clknet_leaf_213_clk),
    .Q(\cs_registers_i.mscratch_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00329_),
    .RN(net148),
    .CLK(clknet_6_24__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00330_),
    .RN(net3660),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00331_),
    .RN(net148),
    .CLK(clknet_6_33__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00332_),
    .RN(net148),
    .CLK(clknet_leaf_0_clk),
    .Q(\cs_registers_i.mscratch_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00333_),
    .RN(net148),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mscratch_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00334_),
    .RN(net3660),
    .CLK(clknet_leaf_66_clk),
    .Q(\cs_registers_i.mscratch_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00335_),
    .RN(net148),
    .CLK(clknet_leaf_44_clk),
    .Q(\cs_registers_i.mscratch_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00336_),
    .RN(net148),
    .CLK(clknet_leaf_48_clk),
    .Q(\cs_registers_i.mscratch_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00337_),
    .RN(net148),
    .CLK(clknet_6_26__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00338_),
    .RN(net3660),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.mscratch_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00339_),
    .RN(net148),
    .CLK(clknet_leaf_25_clk),
    .Q(\cs_registers_i.mstack_cause_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00340_),
    .RN(net148),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mstack_cause_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00341_),
    .RN(net148),
    .CLK(clknet_leaf_42_clk),
    .Q(\cs_registers_i.mstack_cause_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00342_),
    .RN(net148),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mstack_cause_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00343_),
    .RN(net148),
    .CLK(clknet_leaf_0_clk),
    .Q(\cs_registers_i.mstack_cause_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00344_),
    .RN(net148),
    .CLK(clknet_leaf_109_clk),
    .Q(\cs_registers_i.mstack_cause_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00345_),
    .RN(net3661),
    .CLK(clknet_leaf_35_clk),
    .Q(\cs_registers_i.mstack_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00346_),
    .RN(net148),
    .CLK(clknet_leaf_35_clk),
    .Q(\cs_registers_i.mstack_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \cs_registers_i.u_mstack_csr.rd_data_o[2]$_DFFE_PN1P_  (.D(_00347_),
    .SETN(net3660),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\cs_registers_i.mstack_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00348_),
    .RN(net148),
    .CLK(clknet_leaf_610_clk),
    .Q(\cs_registers_i.mstack_epc_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00349_),
    .RN(net148),
    .CLK(clknet_leaf_298_clk),
    .Q(\cs_registers_i.mstack_epc_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00350_),
    .RN(net3660),
    .CLK(clknet_leaf_71_clk),
    .Q(\cs_registers_i.mstack_epc_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00351_),
    .RN(net3660),
    .CLK(clknet_leaf_84_clk),
    .Q(\cs_registers_i.mstack_epc_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00352_),
    .RN(net3660),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00353_),
    .RN(net3660),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00354_),
    .RN(net148),
    .CLK(clknet_leaf_95_clk),
    .Q(\cs_registers_i.mstack_epc_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00355_),
    .RN(net3660),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00356_),
    .RN(net3660),
    .CLK(clknet_leaf_266_clk),
    .Q(\cs_registers_i.mstack_epc_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00357_),
    .RN(net3660),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00358_),
    .RN(net3660),
    .CLK(clknet_leaf_286_clk),
    .Q(\cs_registers_i.mstack_epc_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00359_),
    .RN(net148),
    .CLK(clknet_6_13__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00360_),
    .RN(net148),
    .CLK(clknet_leaf_91_clk),
    .Q(\cs_registers_i.mstack_epc_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00361_),
    .RN(net3660),
    .CLK(clknet_leaf_288_clk),
    .Q(\cs_registers_i.mstack_epc_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00362_),
    .RN(net3660),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00363_),
    .RN(net3660),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00364_),
    .RN(net3660),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00365_),
    .RN(net3660),
    .CLK(clknet_leaf_229_clk),
    .Q(\cs_registers_i.mstack_epc_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00366_),
    .RN(net3660),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00367_),
    .RN(net3660),
    .CLK(clknet_leaf_195_clk),
    .Q(\cs_registers_i.mstack_epc_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00368_),
    .RN(net3660),
    .CLK(clknet_leaf_220_clk),
    .Q(\cs_registers_i.mstack_epc_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00369_),
    .RN(net3660),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00370_),
    .RN(net148),
    .CLK(clknet_leaf_38_clk),
    .Q(\cs_registers_i.mstack_epc_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00371_),
    .RN(net3660),
    .CLK(clknet_leaf_296_clk),
    .Q(\cs_registers_i.mstack_epc_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00372_),
    .RN(net148),
    .CLK(clknet_leaf_110_clk),
    .Q(\cs_registers_i.mstack_epc_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00373_),
    .RN(net148),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00374_),
    .RN(net148),
    .CLK(clknet_6_9__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00375_),
    .RN(net3660),
    .CLK(clknet_6_15__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00376_),
    .RN(net148),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00377_),
    .RN(net148),
    .CLK(clknet_leaf_54_clk),
    .Q(\cs_registers_i.mstack_epc_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00378_),
    .RN(net3660),
    .CLK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.mstack_epc_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00379_),
    .RN(net3660),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.mstack_epc_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00380_),
    .RN(net3660),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\cs_registers_i.csr_mstatus_tw_o ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00381_),
    .RN(net3660),
    .CLK(clknet_leaf_85_clk),
    .Q(\cs_registers_i.mstatus_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[2]$_DFFE_PN0N_  (.D(_00382_),
    .RN(net3660),
    .CLK(clknet_leaf_41_clk),
    .Q(\cs_registers_i.mstatus_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[3]$_DFFE_PN0N_  (.D(_00383_),
    .RN(net3660),
    .CLK(clknet_leaf_41_clk),
    .Q(\cs_registers_i.mstatus_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \cs_registers_i.u_mstatus_csr.rd_data_o[4]$_DFFE_PN1N_  (.D(_00384_),
    .SETN(net3660),
    .CLK(clknet_leaf_40_clk),
    .Q(\cs_registers_i.mstatus_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[5]$_DFFE_PN0N_  (.D(_00385_),
    .RN(net3660),
    .CLK(clknet_leaf_40_clk),
    .Q(\cs_registers_i.csr_mstatus_mie_o ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_00386_),
    .RN(net148),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00387_),
    .RN(net148),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.mtval_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00388_),
    .RN(net3660),
    .CLK(clknet_leaf_61_clk),
    .Q(\cs_registers_i.mtval_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00389_),
    .RN(net3660),
    .CLK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.mtval_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00390_),
    .RN(net148),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.mtval_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00391_),
    .RN(net3660),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.mtval_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00392_),
    .RN(net148),
    .CLK(clknet_leaf_293_clk),
    .Q(\cs_registers_i.mtval_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00393_),
    .RN(net3660),
    .CLK(clknet_leaf_88_clk),
    .Q(\cs_registers_i.mtval_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00394_),
    .RN(net3660),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.mtval_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00395_),
    .RN(net148),
    .CLK(clknet_leaf_154_clk),
    .Q(\cs_registers_i.mtval_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00396_),
    .RN(net3660),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\cs_registers_i.mtval_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_00397_),
    .RN(net148),
    .CLK(clknet_leaf_38_clk),
    .Q(\cs_registers_i.mtval_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00398_),
    .RN(net3660),
    .CLK(clknet_leaf_288_clk),
    .Q(\cs_registers_i.mtval_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00399_),
    .RN(net3660),
    .CLK(clknet_leaf_288_clk),
    .Q(\cs_registers_i.mtval_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00400_),
    .RN(net3660),
    .CLK(clknet_leaf_267_clk),
    .Q(\cs_registers_i.mtval_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00401_),
    .RN(net3660),
    .CLK(clknet_leaf_265_clk),
    .Q(\cs_registers_i.mtval_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00402_),
    .RN(net3660),
    .CLK(clknet_leaf_267_clk),
    .Q(\cs_registers_i.mtval_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00403_),
    .RN(net3660),
    .CLK(clknet_leaf_265_clk),
    .Q(\cs_registers_i.mtval_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00404_),
    .RN(net148),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\cs_registers_i.mtval_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00405_),
    .RN(net148),
    .CLK(clknet_leaf_154_clk),
    .Q(\cs_registers_i.mtval_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00406_),
    .RN(net148),
    .CLK(clknet_6_41__leaf_clk),
    .Q(\cs_registers_i.mtval_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00407_),
    .RN(net3660),
    .CLK(clknet_6_44__leaf_clk),
    .Q(\cs_registers_i.mtval_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_00408_),
    .RN(net148),
    .CLK(clknet_leaf_45_clk),
    .Q(\cs_registers_i.mtval_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00409_),
    .RN(net3660),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.mtval_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00410_),
    .RN(net148),
    .CLK(clknet_leaf_104_clk),
    .Q(\cs_registers_i.mtval_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_00411_),
    .RN(net148),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.mtval_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_00412_),
    .RN(net148),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.mtval_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_00413_),
    .RN(net148),
    .CLK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.mtval_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_00414_),
    .RN(net148),
    .CLK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.mtval_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_00415_),
    .RN(net148),
    .CLK(clknet_leaf_53_clk),
    .Q(\cs_registers_i.mtval_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00416_),
    .RN(net148),
    .CLK(clknet_leaf_52_clk),
    .Q(\cs_registers_i.mtval_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00417_),
    .RN(net3660),
    .CLK(clknet_leaf_293_clk),
    .Q(\cs_registers_i.mtval_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_00418_),
    .RN(net3660),
    .CLK(clknet_leaf_58_clk),
    .Q(\cs_registers_i.csr_mtvec_o[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_00419_),
    .RN(net3660),
    .CLK(clknet_leaf_73_clk),
    .Q(\cs_registers_i.csr_mtvec_o[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_00420_),
    .RN(net3660),
    .CLK(clknet_leaf_72_clk),
    .Q(\cs_registers_i.csr_mtvec_o[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_00421_),
    .RN(net3660),
    .CLK(clknet_6_36__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_00422_),
    .RN(net3660),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_00423_),
    .RN(net148),
    .CLK(clknet_leaf_93_clk),
    .Q(\cs_registers_i.csr_mtvec_o[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_00424_),
    .RN(net3660),
    .CLK(clknet_leaf_209_clk),
    .Q(\cs_registers_i.csr_mtvec_o[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_00425_),
    .RN(net3660),
    .CLK(clknet_leaf_272_clk),
    .Q(\cs_registers_i.csr_mtvec_o[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_00426_),
    .RN(net3660),
    .CLK(clknet_leaf_191_clk),
    .Q(\cs_registers_i.csr_mtvec_o[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_00427_),
    .RN(net3660),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_00428_),
    .RN(net148),
    .CLK(clknet_6_35__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_00429_),
    .RN(net3660),
    .CLK(clknet_6_38__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_00430_),
    .RN(net3660),
    .CLK(clknet_leaf_218_clk),
    .Q(\cs_registers_i.csr_mtvec_o[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_00431_),
    .RN(net3660),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_00432_),
    .RN(net3660),
    .CLK(clknet_leaf_191_clk),
    .Q(\cs_registers_i.csr_mtvec_o[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_00433_),
    .RN(net3660),
    .CLK(clknet_leaf_218_clk),
    .Q(\cs_registers_i.csr_mtvec_o[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_00434_),
    .RN(net3660),
    .CLK(clknet_6_43__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_00435_),
    .RN(net3660),
    .CLK(clknet_6_46__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_00436_),
    .RN(net3660),
    .CLK(clknet_leaf_207_clk),
    .Q(\cs_registers_i.csr_mtvec_o[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_00437_),
    .RN(net3660),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_00438_),
    .RN(net3660),
    .CLK(clknet_leaf_277_clk),
    .Q(\cs_registers_i.csr_mtvec_o[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_00439_),
    .RN(net148),
    .CLK(clknet_6_14__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_00440_),
    .RN(net3660),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\cs_registers_i.csr_mtvec_o[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_00441_),
    .RN(net3660),
    .CLK(clknet_leaf_275_clk),
    .Q(\cs_registers_i.csr_mtvec_o[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.D(_00442_),
    .RN(net3660),
    .CLK(clknet_leaf_383_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.D(_00443_),
    .RN(net3660),
    .CLK(clknet_leaf_377_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.D(_00444_),
    .RN(net3660),
    .CLK(clknet_leaf_378_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.D(_00445_),
    .RN(net3660),
    .CLK(clknet_leaf_377_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.D(_00446_),
    .RN(net3660),
    .CLK(clknet_leaf_378_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.D(_00447_),
    .RN(net3660),
    .CLK(clknet_6_62__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.D(_00000_),
    .SETN(net148),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.D(_00001_),
    .RN(net148),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.D(_00002_),
    .RN(net3660),
    .CLK(clknet_6_62__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.D(_00003_),
    .RN(net3660),
    .CLK(clknet_leaf_384_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.D(_00004_),
    .RN(net3660),
    .CLK(clknet_leaf_382_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.D(_00005_),
    .RN(net3660),
    .CLK(clknet_6_62__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.D(_00448_),
    .RN(net3660),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.D(_00449_),
    .RN(net3660),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.D(_00450_),
    .RN(net3660),
    .CLK(clknet_leaf_336_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.D(_00451_),
    .RN(net3660),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.D(_00452_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.D(_00453_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.D(_00454_),
    .RN(net3660),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.D(_00455_),
    .RN(net3660),
    .CLK(clknet_leaf_332_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.D(_00456_),
    .RN(net3660),
    .CLK(clknet_leaf_331_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.D(_00457_),
    .RN(net3660),
    .CLK(clknet_leaf_331_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.D(_00458_),
    .RN(net3660),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.D(_00459_),
    .RN(net3660),
    .CLK(clknet_leaf_332_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.D(_00460_),
    .RN(net3660),
    .CLK(clknet_leaf_335_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.D(_00461_),
    .RN(net3660),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.D(_00462_),
    .RN(net3660),
    .CLK(clknet_leaf_335_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.D(_00463_),
    .RN(net3660),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.D(_00464_),
    .RN(net3660),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.D(_00465_),
    .RN(net3660),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.D(_00466_),
    .RN(net3660),
    .CLK(clknet_leaf_385_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.D(_00467_),
    .RN(net3660),
    .CLK(clknet_leaf_385_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.D(_00468_),
    .RN(net3660),
    .CLK(clknet_leaf_383_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.D(_00469_),
    .RN(net3660),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.D(_00470_),
    .RN(net3660),
    .CLK(clknet_leaf_390_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.D(_00471_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.D(_00472_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.D(_00473_),
    .RN(net3660),
    .CLK(clknet_leaf_390_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.D(_00474_),
    .RN(net3660),
    .CLK(clknet_leaf_328_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.D(_00475_),
    .RN(net3660),
    .CLK(clknet_leaf_328_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.D(_00476_),
    .RN(net3660),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.D(_00477_),
    .RN(net3660),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.D(_00478_),
    .RN(net3660),
    .CLK(clknet_leaf_336_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.D(_00479_),
    .RN(net3660),
    .CLK(clknet_leaf_336_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.D(_00480_),
    .RN(net3660),
    .CLK(clknet_leaf_406_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.D(_00481_),
    .RN(net3660),
    .CLK(clknet_leaf_408_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.D(_00482_),
    .RN(net3660),
    .CLK(clknet_leaf_410_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.D(_00483_),
    .RN(net3660),
    .CLK(clknet_leaf_410_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.D(_00484_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.D(_00485_),
    .RN(net3660),
    .CLK(clknet_leaf_423_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.D(_00486_),
    .RN(net3660),
    .CLK(clknet_leaf_423_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.D(_00487_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.D(_00488_),
    .RN(net3660),
    .CLK(clknet_leaf_407_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.D(_00489_),
    .RN(net3660),
    .CLK(clknet_leaf_420_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.D(_00490_),
    .RN(net3660),
    .CLK(clknet_leaf_420_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.D(_00491_),
    .RN(net3660),
    .CLK(clknet_leaf_407_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.D(_00492_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.D(_00493_),
    .RN(net3660),
    .CLK(clknet_leaf_420_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.D(_00494_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.D(_00495_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.D(_00496_),
    .RN(net3660),
    .CLK(clknet_leaf_413_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.D(_00497_),
    .RN(net3660),
    .CLK(clknet_leaf_413_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.D(_00498_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.D(_00499_),
    .RN(net3660),
    .CLK(clknet_leaf_426_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.D(_00500_),
    .RN(net3660),
    .CLK(clknet_leaf_413_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.D(_00501_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.D(_00502_),
    .RN(net3660),
    .CLK(clknet_leaf_409_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.D(_00503_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.D(_00504_),
    .RN(net3660),
    .CLK(clknet_6_62__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.D(_00505_),
    .RN(net3660),
    .CLK(clknet_leaf_403_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.D(_00506_),
    .RN(net3660),
    .CLK(clknet_leaf_406_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.D(_00507_),
    .RN(net3660),
    .CLK(clknet_leaf_409_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.D(_00508_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.D(_00509_),
    .RN(net3660),
    .CLK(clknet_leaf_403_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.D(_00510_),
    .RN(net3660),
    .CLK(clknet_leaf_407_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.D(_00511_),
    .RN(net3660),
    .CLK(clknet_leaf_408_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \fetch_enable_q$_DFFE_PN0P_  (.D(_00512_),
    .RN(net148),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(fetch_enable_q));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1000]$_DFFE_PN0P_  (.D(_00513_),
    .RN(net3661),
    .CLK(clknet_6_17__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1000] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1001]$_DFFE_PN0P_  (.D(_00514_),
    .RN(net3661),
    .CLK(clknet_leaf_561_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1001] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1002]$_DFFE_PN0P_  (.D(_00515_),
    .RN(net3661),
    .CLK(clknet_leaf_563_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1002] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1003]$_DFFE_PN0P_  (.D(_00516_),
    .RN(net3663),
    .CLK(clknet_6_37__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1003] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1004]$_DFFE_PN0P_  (.D(_00517_),
    .RN(net3663),
    .CLK(clknet_6_47__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1004] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1005]$_DFFE_PN0P_  (.D(_00518_),
    .RN(net3663),
    .CLK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1005] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1006]$_DFFE_PN0P_  (.D(_00519_),
    .RN(net3661),
    .CLK(clknet_leaf_407_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1006] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1007]$_DFFE_PN0P_  (.D(_00520_),
    .RN(net3662),
    .CLK(clknet_leaf_389_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1007] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1008]$_DFFE_PN0P_  (.D(_00521_),
    .RN(net3662),
    .CLK(clknet_6_11__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1008] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1009]$_DFFE_PN0P_  (.D(_00522_),
    .RN(net3662),
    .CLK(clknet_6_7__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1009] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[100]$_DFFE_PN0P_  (.D(_00523_),
    .RN(net3662),
    .CLK(clknet_leaf_215_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[100] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1010]$_DFFE_PN0P_  (.D(_00524_),
    .RN(net3663),
    .CLK(clknet_6_59__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1010] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1011]$_DFFE_PN0P_  (.D(_00525_),
    .RN(net3662),
    .CLK(clknet_leaf_280_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1011] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1012]$_DFFE_PN0P_  (.D(_00526_),
    .RN(net3664),
    .CLK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1012] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1013]$_DFFE_PN0P_  (.D(_00527_),
    .RN(net3663),
    .CLK(clknet_leaf_197_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1013] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1014]$_DFFE_PN0P_  (.D(_00528_),
    .RN(net3662),
    .CLK(clknet_leaf_325_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1014] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1015]$_DFFE_PN0P_  (.D(_00529_),
    .RN(net3661),
    .CLK(clknet_leaf_403_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1015] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1016]$_DFFE_PN0P_  (.D(_00530_),
    .RN(net3662),
    .CLK(clknet_leaf_343_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1016] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1017]$_DFFE_PN0P_  (.D(_00531_),
    .RN(net3663),
    .CLK(clknet_leaf_182_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1017] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1018]$_DFFE_PN0P_  (.D(_00532_),
    .RN(net3663),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1018] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1019]$_DFFE_PN0P_  (.D(_00533_),
    .RN(net3663),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1019] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[101]$_DFFE_PN0P_  (.D(_00534_),
    .RN(net3662),
    .CLK(clknet_6_4__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[101] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1020]$_DFFE_PN0P_  (.D(_00535_),
    .RN(net3663),
    .CLK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1020] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1021]$_DFFE_PN0P_  (.D(_00536_),
    .RN(net3663),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1021] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1022]$_DFFE_PN0P_  (.D(_00537_),
    .RN(net3663),
    .CLK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1022] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1023]$_DFFE_PN0P_  (.D(_00538_),
    .RN(net3662),
    .CLK(clknet_leaf_252_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1023] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[102]$_DFFE_PN0P_  (.D(_00539_),
    .RN(net3662),
    .CLK(clknet_leaf_468_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[102] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[103]$_DFFE_PN0P_  (.D(_00540_),
    .RN(net3661),
    .CLK(clknet_6_28__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[103] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[104]$_DFFE_PN0P_  (.D(_00541_),
    .RN(net3661),
    .CLK(clknet_leaf_531_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[104] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[105]$_DFFE_PN0P_  (.D(_00542_),
    .RN(net3661),
    .CLK(clknet_leaf_526_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[105] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[106]$_DFFE_PN0P_  (.D(_00543_),
    .RN(net3661),
    .CLK(clknet_leaf_488_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[106] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[107]$_DFFE_PN0P_  (.D(_00544_),
    .RN(net3663),
    .CLK(clknet_leaf_469_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[107] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[108]$_DFFE_PN0P_  (.D(_00545_),
    .RN(net3663),
    .CLK(clknet_leaf_167_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[108] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[109]$_DFFE_PN0P_  (.D(_00546_),
    .RN(net3663),
    .CLK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[109] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[110]$_DFFE_PN0P_  (.D(_00547_),
    .RN(net3662),
    .CLK(clknet_leaf_426_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[110] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[111]$_DFFE_PN0P_  (.D(_00548_),
    .RN(net3662),
    .CLK(clknet_leaf_428_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[111] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[112]$_DFFE_PN0P_  (.D(_00549_),
    .RN(net3662),
    .CLK(clknet_leaf_320_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[112] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[113]$_DFFE_PN0P_  (.D(_00550_),
    .RN(net3662),
    .CLK(clknet_leaf_443_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[113] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[114]$_DFFE_PN0P_  (.D(_00551_),
    .RN(net3663),
    .CLK(clknet_6_59__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[114] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[115]$_DFFE_PN0P_  (.D(_00552_),
    .RN(net3663),
    .CLK(clknet_leaf_147_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[115] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[116]$_DFFE_PN0P_  (.D(_00553_),
    .RN(net3664),
    .CLK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[116] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[117]$_DFFE_PN0P_  (.D(_00554_),
    .RN(net3662),
    .CLK(clknet_leaf_266_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[117] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[118]$_DFFE_PN0P_  (.D(_00555_),
    .RN(net3662),
    .CLK(clknet_leaf_317_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[118] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[119]$_DFFE_PN0P_  (.D(_00556_),
    .RN(net3661),
    .CLK(clknet_6_4__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[119] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[120]$_DFFE_PN0P_  (.D(_00557_),
    .RN(net3662),
    .CLK(clknet_6_9__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[120] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[121]$_DFFE_PN0P_  (.D(_00558_),
    .RN(net3663),
    .CLK(clknet_6_35__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[121] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[122]$_DFFE_PN0P_  (.D(_00559_),
    .RN(net3663),
    .CLK(clknet_leaf_202_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[122] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[123]$_DFFE_PN0P_  (.D(_00560_),
    .RN(net3663),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[123] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[124]$_DFFE_PN0P_  (.D(_00561_),
    .RN(net3663),
    .CLK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[124] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[125]$_DFFE_PN0P_  (.D(_00562_),
    .RN(net3663),
    .CLK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[125] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[126]$_DFFE_PN0P_  (.D(_00563_),
    .RN(net3663),
    .CLK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[126] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[127]$_DFFE_PN0P_  (.D(_00564_),
    .RN(net3662),
    .CLK(clknet_leaf_237_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[127] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[128]$_DFFE_PN0P_  (.D(_00565_),
    .RN(net3662),
    .CLK(clknet_leaf_312_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[128] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[129]$_DFFE_PN0P_  (.D(_00566_),
    .RN(net3661),
    .CLK(clknet_leaf_535_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[129] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[130]$_DFFE_PN0P_  (.D(_00567_),
    .RN(net3662),
    .CLK(clknet_6_40__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[130] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[131]$_DFFE_PN0P_  (.D(_00568_),
    .RN(net3662),
    .CLK(clknet_leaf_307_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[131] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[132]$_DFFE_PN0P_  (.D(_00569_),
    .RN(net3662),
    .CLK(clknet_6_33__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[132] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[133]$_DFFE_PN0P_  (.D(_00570_),
    .RN(net3661),
    .CLK(clknet_leaf_420_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[133] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[134]$_DFFE_PN0P_  (.D(_00571_),
    .RN(net3662),
    .CLK(clknet_6_30__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[134] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[135]$_DFFE_PN0P_  (.D(_00572_),
    .RN(net3661),
    .CLK(clknet_leaf_486_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[135] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[136]$_DFFE_PN0P_  (.D(_00573_),
    .RN(net3661),
    .CLK(clknet_leaf_533_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[136] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[137]$_DFFE_PN0P_  (.D(_00574_),
    .RN(net3661),
    .CLK(clknet_leaf_528_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[137] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[138]$_DFFE_PN0P_  (.D(_00575_),
    .RN(net3661),
    .CLK(clknet_leaf_493_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[138] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[139]$_DFFE_PN0P_  (.D(_00576_),
    .RN(net3663),
    .CLK(clknet_leaf_214_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[139] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[140]$_DFFE_PN0P_  (.D(_00577_),
    .RN(net3663),
    .CLK(clknet_leaf_136_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[140] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[141]$_DFFE_PN0P_  (.D(_00578_),
    .RN(net3663),
    .CLK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[141] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[142]$_DFFE_PN0P_  (.D(_00579_),
    .RN(net3662),
    .CLK(clknet_leaf_430_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[142] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[143]$_DFFE_PN0P_  (.D(_00580_),
    .RN(net3662),
    .CLK(clknet_leaf_428_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[143] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[144]$_DFFE_PN0P_  (.D(_00581_),
    .RN(net3662),
    .CLK(clknet_leaf_322_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[144] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[145]$_DFFE_PN0P_  (.D(_00582_),
    .RN(net3662),
    .CLK(clknet_6_5__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[145] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[146]$_DFFE_PN0P_  (.D(_00583_),
    .RN(net3664),
    .CLK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[146] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[147]$_DFFE_PN0P_  (.D(_00584_),
    .RN(net3662),
    .CLK(clknet_leaf_280_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[147] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[148]$_DFFE_PN0P_  (.D(_00585_),
    .RN(net3664),
    .CLK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[148] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[149]$_DFFE_PN0P_  (.D(_00586_),
    .RN(net3663),
    .CLK(clknet_leaf_158_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[149] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[150]$_DFFE_PN0P_  (.D(_00587_),
    .RN(net3662),
    .CLK(clknet_leaf_325_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[150] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[151]$_DFFE_PN0P_  (.D(_00588_),
    .RN(net3661),
    .CLK(clknet_6_1__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[151] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[152]$_DFFE_PN0P_  (.D(_00589_),
    .RN(net3662),
    .CLK(clknet_leaf_368_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[152] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[153]$_DFFE_PN0P_  (.D(_00590_),
    .RN(net3663),
    .CLK(clknet_leaf_174_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[153] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[154]$_DFFE_PN0P_  (.D(_00591_),
    .RN(net3663),
    .CLK(clknet_leaf_188_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[154] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[155]$_DFFE_PN0P_  (.D(_00592_),
    .RN(net3663),
    .CLK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[155] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[156]$_DFFE_PN0P_  (.D(_00593_),
    .RN(net3663),
    .CLK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[156] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[157]$_DFFE_PN0P_  (.D(_00594_),
    .RN(net3663),
    .CLK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[157] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[158]$_DFFE_PN0P_  (.D(_00595_),
    .RN(net3663),
    .CLK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[158] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[159]$_DFFE_PN0P_  (.D(_00596_),
    .RN(net3662),
    .CLK(clknet_leaf_252_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[159] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[160]$_DFFE_PN0P_  (.D(_00597_),
    .RN(net3662),
    .CLK(clknet_leaf_312_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[160] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[161]$_DFFE_PN0P_  (.D(_00598_),
    .RN(net3661),
    .CLK(clknet_leaf_536_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[161] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[162]$_DFFE_PN0P_  (.D(_00599_),
    .RN(net3662),
    .CLK(clknet_leaf_276_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[162] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[163]$_DFFE_PN0P_  (.D(_00600_),
    .RN(net3662),
    .CLK(clknet_6_40__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[163] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[164]$_DFFE_PN0P_  (.D(_00601_),
    .RN(net3662),
    .CLK(clknet_6_38__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[164] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[165]$_DFFE_PN0P_  (.D(_00602_),
    .RN(net3661),
    .CLK(clknet_6_27__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[165] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[166]$_DFFE_PN0P_  (.D(_00603_),
    .RN(net3662),
    .CLK(clknet_6_30__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[166] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[167]$_DFFE_PN0P_  (.D(_00604_),
    .RN(net3661),
    .CLK(clknet_6_26__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[167] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[168]$_DFFE_PN0P_  (.D(_00605_),
    .RN(net3661),
    .CLK(clknet_leaf_533_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[168] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[169]$_DFFE_PN0P_  (.D(_00606_),
    .RN(net3661),
    .CLK(clknet_leaf_528_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[169] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[170]$_DFFE_PN0P_  (.D(_00607_),
    .RN(net3661),
    .CLK(clknet_leaf_493_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[170] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[171]$_DFFE_PN0P_  (.D(_00608_),
    .RN(net3663),
    .CLK(clknet_leaf_214_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[171] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[172]$_DFFE_PN0P_  (.D(_00609_),
    .RN(net3663),
    .CLK(clknet_6_58__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[172] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[173]$_DFFE_PN0P_  (.D(_00610_),
    .RN(net3663),
    .CLK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[173] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[174]$_DFFE_PN0P_  (.D(_00611_),
    .RN(net3662),
    .CLK(clknet_leaf_423_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[174] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[175]$_DFFE_PN0P_  (.D(_00612_),
    .RN(net3662),
    .CLK(clknet_leaf_427_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[175] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[176]$_DFFE_PN0P_  (.D(_00613_),
    .RN(net3662),
    .CLK(clknet_leaf_334_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[176] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[177]$_DFFE_PN0P_  (.D(_00614_),
    .RN(net3662),
    .CLK(clknet_leaf_446_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[177] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[178]$_DFFE_PN0P_  (.D(_00615_),
    .RN(net3664),
    .CLK(clknet_6_62__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[178] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[179]$_DFFE_PN0P_  (.D(_00616_),
    .RN(net3662),
    .CLK(clknet_6_46__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[179] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[180]$_DFFE_PN0P_  (.D(_00617_),
    .RN(net3664),
    .CLK(clknet_leaf_80_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[180] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[181]$_DFFE_PN0P_  (.D(_00618_),
    .RN(net3663),
    .CLK(clknet_6_44__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[181] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[182]$_DFFE_PN0P_  (.D(_00619_),
    .RN(net3662),
    .CLK(clknet_leaf_324_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[182] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[183]$_DFFE_PN0P_  (.D(_00620_),
    .RN(net3661),
    .CLK(clknet_leaf_405_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[183] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[184]$_DFFE_PN0P_  (.D(_00621_),
    .RN(net3662),
    .CLK(clknet_leaf_376_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[184] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[185]$_DFFE_PN0P_  (.D(_00622_),
    .RN(net3663),
    .CLK(clknet_leaf_174_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[185] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[186]$_DFFE_PN0P_  (.D(_00623_),
    .RN(net3663),
    .CLK(clknet_leaf_188_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[186] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[187]$_DFFE_PN0P_  (.D(_00624_),
    .RN(net3663),
    .CLK(clknet_leaf_38_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[187] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[188]$_DFFE_PN0P_  (.D(_00625_),
    .RN(net3663),
    .CLK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[188] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[189]$_DFFE_PN0P_  (.D(_00626_),
    .RN(net3663),
    .CLK(clknet_leaf_43_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[189] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[190]$_DFFE_PN0P_  (.D(_00627_),
    .RN(net3663),
    .CLK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[190] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[191]$_DFFE_PN0P_  (.D(_00628_),
    .RN(net3662),
    .CLK(clknet_6_32__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[191] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[192]$_DFFE_PN0P_  (.D(_00629_),
    .RN(net3662),
    .CLK(clknet_6_12__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[192] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[193]$_DFFE_PN0P_  (.D(_00630_),
    .RN(net3661),
    .CLK(clknet_leaf_536_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[193] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[194]$_DFFE_PN0P_  (.D(_00631_),
    .RN(net3662),
    .CLK(clknet_6_41__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[194] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[195]$_DFFE_PN0P_  (.D(_00632_),
    .RN(net3662),
    .CLK(clknet_leaf_308_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[195] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[196]$_DFFE_PN0P_  (.D(_00633_),
    .RN(net3662),
    .CLK(clknet_leaf_226_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[196] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[197]$_DFFE_PN0P_  (.D(_00634_),
    .RN(net3661),
    .CLK(clknet_6_27__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[197] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[198]$_DFFE_PN0P_  (.D(_00635_),
    .RN(net3661),
    .CLK(clknet_leaf_484_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[198] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[199]$_DFFE_PN0P_  (.D(_00636_),
    .RN(net3661),
    .CLK(clknet_leaf_488_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[199] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[200]$_DFFE_PN0P_  (.D(_00637_),
    .RN(net3661),
    .CLK(clknet_leaf_533_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[200] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[201]$_DFFE_PN0P_  (.D(_00638_),
    .RN(net3661),
    .CLK(clknet_leaf_528_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[201] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[202]$_DFFE_PN0P_  (.D(_00639_),
    .RN(net3661),
    .CLK(clknet_leaf_492_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[202] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[203]$_DFFE_PN0P_  (.D(_00640_),
    .RN(net3663),
    .CLK(clknet_leaf_211_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[203] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[204]$_DFFE_PN0P_  (.D(_00641_),
    .RN(net3663),
    .CLK(clknet_leaf_151_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[204] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[205]$_DFFE_PN0P_  (.D(_00642_),
    .RN(net3663),
    .CLK(clknet_leaf_113_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[205] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[206]$_DFFE_PN0P_  (.D(_00643_),
    .RN(net3661),
    .CLK(clknet_leaf_424_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[206] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[207]$_DFFE_PN0P_  (.D(_00644_),
    .RN(net3662),
    .CLK(clknet_leaf_427_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[207] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[208]$_DFFE_PN0P_  (.D(_00645_),
    .RN(net3662),
    .CLK(clknet_leaf_352_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[208] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[209]$_DFFE_PN0P_  (.D(_00646_),
    .RN(net3662),
    .CLK(clknet_leaf_446_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[209] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[210]$_DFFE_PN0P_  (.D(_00647_),
    .RN(net3664),
    .CLK(clknet_6_62__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[210] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[211]$_DFFE_PN0P_  (.D(_00648_),
    .RN(net3662),
    .CLK(clknet_leaf_278_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[211] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[212]$_DFFE_PN0P_  (.D(_00649_),
    .RN(net3664),
    .CLK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[212] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[213]$_DFFE_PN0P_  (.D(_00650_),
    .RN(net3663),
    .CLK(clknet_leaf_158_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[213] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[214]$_DFFE_PN0P_  (.D(_00651_),
    .RN(net3662),
    .CLK(clknet_leaf_317_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[214] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[215]$_DFFE_PN0P_  (.D(_00652_),
    .RN(net3661),
    .CLK(clknet_6_26__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[215] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[216]$_DFFE_PN0P_  (.D(_00653_),
    .RN(net3662),
    .CLK(clknet_6_3__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[216] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[217]$_DFFE_PN0P_  (.D(_00654_),
    .RN(net3663),
    .CLK(clknet_leaf_166_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[217] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[218]$_DFFE_PN0P_  (.D(_00655_),
    .RN(net3663),
    .CLK(clknet_6_48__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[218] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[219]$_DFFE_PN0P_  (.D(_00656_),
    .RN(net3663),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[219] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[220]$_DFFE_PN0P_  (.D(_00657_),
    .RN(net3663),
    .CLK(clknet_6_54__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[220] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[221]$_DFFE_PN0P_  (.D(_00658_),
    .RN(net3663),
    .CLK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[221] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[222]$_DFFE_PN0P_  (.D(_00659_),
    .RN(net3663),
    .CLK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[222] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[223]$_DFFE_PN0P_  (.D(_00660_),
    .RN(net3662),
    .CLK(clknet_leaf_238_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[223] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[224]$_DFFE_PN0P_  (.D(_00661_),
    .RN(net3662),
    .CLK(clknet_leaf_248_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[224] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[225]$_DFFE_PN0P_  (.D(_00662_),
    .RN(net3661),
    .CLK(clknet_leaf_536_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[225] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[226]$_DFFE_PN0P_  (.D(_00663_),
    .RN(net3662),
    .CLK(clknet_leaf_255_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[226] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[227]$_DFFE_PN0P_  (.D(_00664_),
    .RN(net3662),
    .CLK(clknet_leaf_307_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[227] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[228]$_DFFE_PN0P_  (.D(_00665_),
    .RN(net3662),
    .CLK(clknet_6_33__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[228] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[229]$_DFFE_PN0P_  (.D(_00666_),
    .RN(net3661),
    .CLK(clknet_6_27__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[229] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[230]$_DFFE_PN0P_  (.D(_00667_),
    .RN(net3662),
    .CLK(clknet_leaf_484_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[230] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[231]$_DFFE_PN0P_  (.D(_00668_),
    .RN(net3661),
    .CLK(clknet_leaf_488_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[231] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[232]$_DFFE_PN0P_  (.D(_00669_),
    .RN(net3661),
    .CLK(clknet_leaf_533_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[232] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[233]$_DFFE_PN0P_  (.D(_00670_),
    .RN(net3661),
    .CLK(clknet_6_24__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[233] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[234]$_DFFE_PN0P_  (.D(_00671_),
    .RN(net3661),
    .CLK(clknet_leaf_492_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[234] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[235]$_DFFE_PN0P_  (.D(_00672_),
    .RN(net3663),
    .CLK(clknet_leaf_211_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[235] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[236]$_DFFE_PN0P_  (.D(_00673_),
    .RN(net3663),
    .CLK(clknet_leaf_151_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[236] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[237]$_DFFE_PN0P_  (.D(_00674_),
    .RN(net3663),
    .CLK(clknet_6_58__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[237] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[238]$_DFFE_PN0P_  (.D(_00675_),
    .RN(net3661),
    .CLK(clknet_leaf_423_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[238] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[239]$_DFFE_PN0P_  (.D(_00676_),
    .RN(net3662),
    .CLK(clknet_leaf_427_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[239] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[240]$_DFFE_PN0P_  (.D(_00677_),
    .RN(net3662),
    .CLK(clknet_leaf_334_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[240] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[241]$_DFFE_PN0P_  (.D(_00678_),
    .RN(net3662),
    .CLK(clknet_leaf_446_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[241] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[242]$_DFFE_PN0P_  (.D(_00679_),
    .RN(net3664),
    .CLK(clknet_leaf_90_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[242] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[243]$_DFFE_PN0P_  (.D(_00680_),
    .RN(net3662),
    .CLK(clknet_leaf_278_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[243] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[244]$_DFFE_PN0P_  (.D(_00681_),
    .RN(net3664),
    .CLK(clknet_leaf_79_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[244] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[245]$_DFFE_PN0P_  (.D(_00682_),
    .RN(net3663),
    .CLK(clknet_6_35__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[245] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[246]$_DFFE_PN0P_  (.D(_00683_),
    .RN(net3662),
    .CLK(clknet_leaf_317_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[246] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[247]$_DFFE_PN0P_  (.D(_00684_),
    .RN(net3661),
    .CLK(clknet_6_27__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[247] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[248]$_DFFE_PN0P_  (.D(_00685_),
    .RN(net3662),
    .CLK(clknet_leaf_368_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[248] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[249]$_DFFE_PN0P_  (.D(_00686_),
    .RN(net3663),
    .CLK(clknet_leaf_166_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[249] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[250]$_DFFE_PN0P_  (.D(_00687_),
    .RN(net3663),
    .CLK(clknet_leaf_202_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[250] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[251]$_DFFE_PN0P_  (.D(_00688_),
    .RN(net3663),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[251] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[252]$_DFFE_PN0P_  (.D(_00689_),
    .RN(net3663),
    .CLK(clknet_leaf_102_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[252] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[253]$_DFFE_PN0P_  (.D(_00690_),
    .RN(net3663),
    .CLK(clknet_6_55__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[253] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[254]$_DFFE_PN0P_  (.D(_00691_),
    .RN(net3663),
    .CLK(clknet_leaf_47_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[254] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[255]$_DFFE_PN0P_  (.D(_00692_),
    .RN(net3662),
    .CLK(clknet_leaf_238_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[255] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[256]$_DFFE_PN0P_  (.D(_00693_),
    .RN(net3662),
    .CLK(clknet_leaf_361_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[256] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[257]$_DFFE_PN0P_  (.D(_00694_),
    .RN(net3661),
    .CLK(clknet_leaf_525_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[257] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[258]$_DFFE_PN0P_  (.D(_00695_),
    .RN(net3662),
    .CLK(clknet_6_40__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[258] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[259]$_DFFE_PN0P_  (.D(_00696_),
    .RN(net3662),
    .CLK(clknet_leaf_250_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[259] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[260]$_DFFE_PN0P_  (.D(_00697_),
    .RN(net3662),
    .CLK(clknet_leaf_219_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[260] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[261]$_DFFE_PN0P_  (.D(_00698_),
    .RN(net3662),
    .CLK(clknet_leaf_447_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[261] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[262]$_DFFE_PN0P_  (.D(_00699_),
    .RN(net3663),
    .CLK(clknet_leaf_476_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[262] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[263]$_DFFE_PN0P_  (.D(_00700_),
    .RN(net3661),
    .CLK(clknet_leaf_483_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[263] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[264]$_DFFE_PN0P_  (.D(_00701_),
    .RN(net3661),
    .CLK(clknet_leaf_516_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[264] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[265]$_DFFE_PN0P_  (.D(_00702_),
    .RN(net3661),
    .CLK(clknet_6_19__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[265] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[266]$_DFFE_PN0P_  (.D(_00703_),
    .RN(net3661),
    .CLK(clknet_leaf_513_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[266] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[267]$_DFFE_PN0P_  (.D(_00704_),
    .RN(net3663),
    .CLK(clknet_leaf_469_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[267] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[268]$_DFFE_PN0P_  (.D(_00705_),
    .RN(net3663),
    .CLK(clknet_6_45__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[268] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[269]$_DFFE_PN0P_  (.D(_00706_),
    .RN(net3663),
    .CLK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[269] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[270]$_DFFE_PN0P_  (.D(_00707_),
    .RN(net3662),
    .CLK(clknet_leaf_422_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[270] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[271]$_DFFE_PN0P_  (.D(_00708_),
    .RN(net3662),
    .CLK(clknet_leaf_371_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[271] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[272]$_DFFE_PN0P_  (.D(_00709_),
    .RN(net3662),
    .CLK(clknet_leaf_338_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[272] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[273]$_DFFE_PN0P_  (.D(_00710_),
    .RN(net3662),
    .CLK(clknet_6_6__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[273] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[274]$_DFFE_PN0P_  (.D(_00711_),
    .RN(net3663),
    .CLK(clknet_6_59__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[274] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[275]$_DFFE_PN0P_  (.D(_00712_),
    .RN(net3663),
    .CLK(clknet_6_44__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[275] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[276]$_DFFE_PN0P_  (.D(_00713_),
    .RN(net3663),
    .CLK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[276] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[277]$_DFFE_PN0P_  (.D(_00714_),
    .RN(net3663),
    .CLK(clknet_leaf_162_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[277] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[278]$_DFFE_PN0P_  (.D(_00715_),
    .RN(net3662),
    .CLK(clknet_leaf_301_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[278] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[279]$_DFFE_PN0P_  (.D(_00716_),
    .RN(net3661),
    .CLK(clknet_leaf_412_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[279] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[280]$_DFFE_PN0P_  (.D(_00717_),
    .RN(net3662),
    .CLK(clknet_leaf_347_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[280] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[281]$_DFFE_PN0P_  (.D(_00718_),
    .RN(net3663),
    .CLK(clknet_leaf_166_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[281] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[282]$_DFFE_PN0P_  (.D(_00719_),
    .RN(net3663),
    .CLK(clknet_leaf_198_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[282] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[283]$_DFFE_PN0P_  (.D(_00720_),
    .RN(net3663),
    .CLK(clknet_6_51__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[283] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[284]$_DFFE_PN0P_  (.D(_00721_),
    .RN(net3663),
    .CLK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[284] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[285]$_DFFE_PN0P_  (.D(_00722_),
    .RN(net3663),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[285] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[286]$_DFFE_PN0P_  (.D(_00723_),
    .RN(net3663),
    .CLK(clknet_6_60__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[286] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[287]$_DFFE_PN0P_  (.D(_00724_),
    .RN(net3662),
    .CLK(clknet_leaf_234_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[287] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[288]$_DFFE_PN0P_  (.D(_00725_),
    .RN(net3662),
    .CLK(clknet_leaf_360_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[288] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[289]$_DFFE_PN0P_  (.D(_00726_),
    .RN(net3661),
    .CLK(clknet_leaf_525_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[289] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[290]$_DFFE_PN0P_  (.D(_00727_),
    .RN(net3662),
    .CLK(clknet_leaf_256_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[290] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[291]$_DFFE_PN0P_  (.D(_00728_),
    .RN(net3662),
    .CLK(clknet_6_40__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[291] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[292]$_DFFE_PN0P_  (.D(_00729_),
    .RN(net3662),
    .CLK(clknet_6_38__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[292] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[293]$_DFFE_PN0P_  (.D(_00730_),
    .RN(net3662),
    .CLK(clknet_6_5__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[293] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[294]$_DFFE_PN0P_  (.D(_00731_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[294] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[295]$_DFFE_PN0P_  (.D(_00732_),
    .RN(net3661),
    .CLK(clknet_leaf_484_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[295] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[296]$_DFFE_PN0P_  (.D(_00733_),
    .RN(net3661),
    .CLK(clknet_leaf_416_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[296] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[297]$_DFFE_PN0P_  (.D(_00734_),
    .RN(net3661),
    .CLK(clknet_leaf_523_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[297] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[298]$_DFFE_PN0P_  (.D(_00735_),
    .RN(net3661),
    .CLK(clknet_leaf_513_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[298] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[299]$_DFFE_PN0P_  (.D(_00736_),
    .RN(net3663),
    .CLK(clknet_leaf_470_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[299] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[300]$_DFFE_PN0P_  (.D(_00737_),
    .RN(net3663),
    .CLK(clknet_leaf_149_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[300] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[301]$_DFFE_PN0P_  (.D(_00738_),
    .RN(net3663),
    .CLK(clknet_leaf_110_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[301] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[302]$_DFFE_PN0P_  (.D(_00739_),
    .RN(net3662),
    .CLK(clknet_leaf_422_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[302] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[303]$_DFFE_PN0P_  (.D(_00740_),
    .RN(net3662),
    .CLK(clknet_leaf_371_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[303] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[304]$_DFFE_PN0P_  (.D(_00741_),
    .RN(net3662),
    .CLK(clknet_leaf_339_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[304] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[305]$_DFFE_PN0P_  (.D(_00742_),
    .RN(net3662),
    .CLK(clknet_leaf_430_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[305] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[306]$_DFFE_PN0P_  (.D(_00743_),
    .RN(net3663),
    .CLK(clknet_6_57__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[306] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[307]$_DFFE_PN0P_  (.D(_00744_),
    .RN(net3663),
    .CLK(clknet_leaf_156_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[307] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[308]$_DFFE_PN0P_  (.D(_00745_),
    .RN(net3663),
    .CLK(clknet_6_61__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[308] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[309]$_DFFE_PN0P_  (.D(_00746_),
    .RN(net3663),
    .CLK(clknet_leaf_162_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[309] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[310]$_DFFE_PN0P_  (.D(_00747_),
    .RN(net3662),
    .CLK(clknet_leaf_301_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[310] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[311]$_DFFE_PN0P_  (.D(_00748_),
    .RN(net3661),
    .CLK(clknet_leaf_404_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[311] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[312]$_DFFE_PN0P_  (.D(_00749_),
    .RN(net3662),
    .CLK(clknet_leaf_347_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[312] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[313]$_DFFE_PN0P_  (.D(_00750_),
    .RN(net3663),
    .CLK(clknet_leaf_165_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[313] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[314]$_DFFE_PN0P_  (.D(_00751_),
    .RN(net3663),
    .CLK(clknet_leaf_198_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[314] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[315]$_DFFE_PN0P_  (.D(_00752_),
    .RN(net3663),
    .CLK(clknet_leaf_179_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[315] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[316]$_DFFE_PN0P_  (.D(_00753_),
    .RN(net3663),
    .CLK(clknet_6_54__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[316] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[317]$_DFFE_PN0P_  (.D(_00754_),
    .RN(net3663),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[317] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[318]$_DFFE_PN0P_  (.D(_00755_),
    .RN(net3663),
    .CLK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[318] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[319]$_DFFE_PN0P_  (.D(_00756_),
    .RN(net3662),
    .CLK(clknet_leaf_234_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[319] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[320]$_DFFE_PN0P_  (.D(_00757_),
    .RN(net3662),
    .CLK(clknet_6_9__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[320] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[321]$_DFFE_PN0P_  (.D(_00758_),
    .RN(net3661),
    .CLK(clknet_leaf_525_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[321] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[322]$_DFFE_PN0P_  (.D(_00759_),
    .RN(net3662),
    .CLK(clknet_6_41__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[322] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[323]$_DFFE_PN0P_  (.D(_00760_),
    .RN(net3662),
    .CLK(clknet_leaf_250_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[323] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[324]$_DFFE_PN0P_  (.D(_00761_),
    .RN(net3662),
    .CLK(clknet_leaf_217_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[324] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[325]$_DFFE_PN0P_  (.D(_00762_),
    .RN(net3662),
    .CLK(clknet_6_4__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[325] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[326]$_DFFE_PN0P_  (.D(_00763_),
    .RN(net3661),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[326] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[327]$_DFFE_PN0P_  (.D(_00764_),
    .RN(net3661),
    .CLK(clknet_leaf_480_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[327] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[328]$_DFFE_PN0P_  (.D(_00765_),
    .RN(net3661),
    .CLK(clknet_leaf_514_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[328] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[329]$_DFFE_PN0P_  (.D(_00766_),
    .RN(net3661),
    .CLK(clknet_6_19__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[329] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[32]$_DFFE_PN0P_  (.D(_00767_),
    .RN(net3662),
    .CLK(clknet_leaf_248_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[330]$_DFFE_PN0P_  (.D(_00768_),
    .RN(net3661),
    .CLK(clknet_leaf_510_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[330] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[331]$_DFFE_PN0P_  (.D(_00769_),
    .RN(net3663),
    .CLK(clknet_leaf_473_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[331] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[332]$_DFFE_PN0P_  (.D(_00770_),
    .RN(net3663),
    .CLK(clknet_leaf_154_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[332] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[333]$_DFFE_PN0P_  (.D(_00771_),
    .RN(net3663),
    .CLK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[333] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[334]$_DFFE_PN0P_  (.D(_00772_),
    .RN(net3662),
    .CLK(clknet_leaf_420_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[334] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[335]$_DFFE_PN0P_  (.D(_00773_),
    .RN(net3662),
    .CLK(clknet_6_3__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[335] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[336]$_DFFE_PN0P_  (.D(_00774_),
    .RN(net3662),
    .CLK(clknet_leaf_339_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[336] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[337]$_DFFE_PN0P_  (.D(_00775_),
    .RN(net3662),
    .CLK(clknet_leaf_431_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[337] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[338]$_DFFE_PN0P_  (.D(_00776_),
    .RN(net3663),
    .CLK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[338] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[339]$_DFFE_PN0P_  (.D(_00777_),
    .RN(net3663),
    .CLK(clknet_6_44__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[339] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[33]$_DFFE_PN0P_  (.D(_00778_),
    .RN(net3661),
    .CLK(clknet_leaf_535_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[340]$_DFFE_PN0P_  (.D(_00779_),
    .RN(net3663),
    .CLK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[340] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[341]$_DFFE_PN0P_  (.D(_00780_),
    .RN(net3663),
    .CLK(clknet_leaf_160_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[341] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[342]$_DFFE_PN0P_  (.D(_00781_),
    .RN(net3662),
    .CLK(clknet_leaf_309_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[342] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[343]$_DFFE_PN0P_  (.D(_00782_),
    .RN(net3661),
    .CLK(clknet_leaf_416_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[343] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[344]$_DFFE_PN0P_  (.D(_00783_),
    .RN(net3662),
    .CLK(clknet_6_8__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[344] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[345]$_DFFE_PN0P_  (.D(_00784_),
    .RN(net3663),
    .CLK(clknet_leaf_191_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[345] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[346]$_DFFE_PN0P_  (.D(_00785_),
    .RN(net3663),
    .CLK(clknet_6_36__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[346] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[347]$_DFFE_PN0P_  (.D(_00786_),
    .RN(net3663),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[347] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[348]$_DFFE_PN0P_  (.D(_00787_),
    .RN(net3663),
    .CLK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[348] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[349]$_DFFE_PN0P_  (.D(_00788_),
    .RN(net3663),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[349] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[34]$_DFFE_PN0P_  (.D(_00789_),
    .RN(net3662),
    .CLK(clknet_6_41__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[350]$_DFFE_PN0P_  (.D(_00790_),
    .RN(net3663),
    .CLK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[350] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[351]$_DFFE_PN0P_  (.D(_00791_),
    .RN(net3662),
    .CLK(clknet_leaf_229_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[351] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[352]$_DFFE_PN0P_  (.D(_00792_),
    .RN(net3662),
    .CLK(clknet_leaf_360_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[352] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[353]$_DFFE_PN0P_  (.D(_00793_),
    .RN(net3661),
    .CLK(clknet_6_19__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[353] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[354]$_DFFE_PN0P_  (.D(_00794_),
    .RN(net3662),
    .CLK(clknet_leaf_256_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[354] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[355]$_DFFE_PN0P_  (.D(_00795_),
    .RN(net3662),
    .CLK(clknet_leaf_250_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[355] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[356]$_DFFE_PN0P_  (.D(_00796_),
    .RN(net3662),
    .CLK(clknet_leaf_217_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[356] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[357]$_DFFE_PN0P_  (.D(_00797_),
    .RN(net3662),
    .CLK(clknet_leaf_447_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[357] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[358]$_DFFE_PN0P_  (.D(_00798_),
    .RN(net3661),
    .CLK(clknet_leaf_478_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[358] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[359]$_DFFE_PN0P_  (.D(_00799_),
    .RN(net3661),
    .CLK(clknet_6_28__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[359] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[35]$_DFFE_PN0P_  (.D(_00800_),
    .RN(net3662),
    .CLK(clknet_leaf_254_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[360]$_DFFE_PN0P_  (.D(_00801_),
    .RN(net3661),
    .CLK(clknet_leaf_516_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[360] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[361]$_DFFE_PN0P_  (.D(_00802_),
    .RN(net3661),
    .CLK(clknet_leaf_522_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[361] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[362]$_DFFE_PN0P_  (.D(_00803_),
    .RN(net3661),
    .CLK(clknet_leaf_513_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[362] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[363]$_DFFE_PN0P_  (.D(_00804_),
    .RN(net3663),
    .CLK(clknet_leaf_473_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[363] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[364]$_DFFE_PN0P_  (.D(_00805_),
    .RN(net3663),
    .CLK(clknet_6_45__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[364] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[365]$_DFFE_PN0P_  (.D(_00806_),
    .RN(net3663),
    .CLK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[365] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[366]$_DFFE_PN0P_  (.D(_00807_),
    .RN(net3662),
    .CLK(clknet_leaf_420_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[366] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[367]$_DFFE_PN0P_  (.D(_00808_),
    .RN(net3662),
    .CLK(clknet_6_3__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[367] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[368]$_DFFE_PN0P_  (.D(_00809_),
    .RN(net3662),
    .CLK(clknet_leaf_339_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[368] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[369]$_DFFE_PN0P_  (.D(_00810_),
    .RN(net3662),
    .CLK(clknet_leaf_431_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[369] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[36]$_DFFE_PN0P_  (.D(_00811_),
    .RN(net3662),
    .CLK(clknet_leaf_215_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[370]$_DFFE_PN0P_  (.D(_00812_),
    .RN(net3663),
    .CLK(clknet_leaf_109_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[370] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[371]$_DFFE_PN0P_  (.D(_00813_),
    .RN(net3663),
    .CLK(clknet_leaf_156_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[371] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[372]$_DFFE_PN0P_  (.D(_00814_),
    .RN(net3663),
    .CLK(clknet_leaf_63_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[372] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[373]$_DFFE_PN0P_  (.D(_00815_),
    .RN(net3663),
    .CLK(clknet_leaf_160_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[373] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[374]$_DFFE_PN0P_  (.D(_00816_),
    .RN(net3662),
    .CLK(clknet_leaf_310_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[374] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[375]$_DFFE_PN0P_  (.D(_00817_),
    .RN(net3661),
    .CLK(clknet_leaf_518_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[375] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[376]$_DFFE_PN0P_  (.D(_00818_),
    .RN(net3662),
    .CLK(clknet_6_8__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[376] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[377]$_DFFE_PN0P_  (.D(_00819_),
    .RN(net3663),
    .CLK(clknet_leaf_191_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[377] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[378]$_DFFE_PN0P_  (.D(_00820_),
    .RN(net3663),
    .CLK(clknet_leaf_200_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[378] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[379]$_DFFE_PN0P_  (.D(_00821_),
    .RN(net3663),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[379] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[37]$_DFFE_PN0P_  (.D(_00822_),
    .RN(net3662),
    .CLK(clknet_leaf_450_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[380]$_DFFE_PN0P_  (.D(_00823_),
    .RN(net3663),
    .CLK(clknet_leaf_40_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[380] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[381]$_DFFE_PN0P_  (.D(_00824_),
    .RN(net3663),
    .CLK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[381] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[382]$_DFFE_PN0P_  (.D(_00825_),
    .RN(net3663),
    .CLK(clknet_leaf_49_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[382] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[383]$_DFFE_PN0P_  (.D(_00826_),
    .RN(net3662),
    .CLK(clknet_leaf_229_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[383] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[384]$_DFFE_PN0P_  (.D(_00827_),
    .RN(net3662),
    .CLK(clknet_6_9__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[384] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[385]$_DFFE_PN0P_  (.D(_00828_),
    .RN(net3661),
    .CLK(clknet_leaf_537_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[385] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[386]$_DFFE_PN0P_  (.D(_00829_),
    .RN(net3662),
    .CLK(clknet_6_41__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[386] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[387]$_DFFE_PN0P_  (.D(_00830_),
    .RN(net3662),
    .CLK(clknet_leaf_251_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[387] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[388]$_DFFE_PN0P_  (.D(_00831_),
    .RN(net3662),
    .CLK(clknet_leaf_219_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[388] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[389]$_DFFE_PN0P_  (.D(_00832_),
    .RN(net3662),
    .CLK(clknet_leaf_462_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[389] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[38]$_DFFE_PN0P_  (.D(_00833_),
    .RN(net3662),
    .CLK(clknet_leaf_468_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[390]$_DFFE_PN0P_  (.D(_00834_),
    .RN(net3663),
    .CLK(clknet_6_29__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[390] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[391]$_DFFE_PN0P_  (.D(_00835_),
    .RN(net3661),
    .CLK(clknet_leaf_483_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[391] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[392]$_DFFE_PN0P_  (.D(_00836_),
    .RN(net3661),
    .CLK(clknet_6_25__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[392] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[393]$_DFFE_PN0P_  (.D(_00837_),
    .RN(net3661),
    .CLK(clknet_leaf_523_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[393] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[394]$_DFFE_PN0P_  (.D(_00838_),
    .RN(net3661),
    .CLK(clknet_6_21__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[394] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[395]$_DFFE_PN0P_  (.D(_00839_),
    .RN(net3663),
    .CLK(clknet_leaf_470_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[395] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[396]$_DFFE_PN0P_  (.D(_00840_),
    .RN(net3663),
    .CLK(clknet_6_45__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[396] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[397]$_DFFE_PN0P_  (.D(_00841_),
    .RN(net3663),
    .CLK(clknet_leaf_171_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[397] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[398]$_DFFE_PN0P_  (.D(_00842_),
    .RN(net3661),
    .CLK(clknet_leaf_408_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[398] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[399]$_DFFE_PN0P_  (.D(_00843_),
    .RN(net3662),
    .CLK(clknet_leaf_375_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[399] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[39]$_DFFE_PN0P_  (.D(_00844_),
    .RN(net3661),
    .CLK(clknet_6_28__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[400]$_DFFE_PN0P_  (.D(_00845_),
    .RN(net3662),
    .CLK(clknet_leaf_352_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[400] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[401]$_DFFE_PN0P_  (.D(_00846_),
    .RN(net3662),
    .CLK(clknet_leaf_440_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[401] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[402]$_DFFE_PN0P_  (.D(_00847_),
    .RN(net3664),
    .CLK(clknet_6_60__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[402] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[403]$_DFFE_PN0P_  (.D(_00848_),
    .RN(net3662),
    .CLK(clknet_leaf_269_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[403] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[404]$_DFFE_PN0P_  (.D(_00849_),
    .RN(net3663),
    .CLK(clknet_6_60__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[404] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[405]$_DFFE_PN0P_  (.D(_00850_),
    .RN(net3662),
    .CLK(clknet_leaf_265_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[405] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[406]$_DFFE_PN0P_  (.D(_00851_),
    .RN(net3662),
    .CLK(clknet_leaf_310_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[406] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[407]$_DFFE_PN0P_  (.D(_00852_),
    .RN(net3661),
    .CLK(clknet_leaf_412_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[407] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[408]$_DFFE_PN0P_  (.D(_00853_),
    .RN(net3662),
    .CLK(clknet_6_2__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[408] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[409]$_DFFE_PN0P_  (.D(_00854_),
    .RN(net3663),
    .CLK(clknet_leaf_183_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[409] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[40]$_DFFE_PN0P_  (.D(_00855_),
    .RN(net3661),
    .CLK(clknet_leaf_531_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[410]$_DFFE_PN0P_  (.D(_00856_),
    .RN(net3663),
    .CLK(clknet_leaf_198_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[410] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[411]$_DFFE_PN0P_  (.D(_00857_),
    .RN(net3663),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[411] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[412]$_DFFE_PN0P_  (.D(_00858_),
    .RN(net3663),
    .CLK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[412] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[413]$_DFFE_PN0P_  (.D(_00859_),
    .RN(net3663),
    .CLK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[413] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[414]$_DFFE_PN0P_  (.D(_00860_),
    .RN(net3663),
    .CLK(clknet_6_60__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[414] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[415]$_DFFE_PN0P_  (.D(_00861_),
    .RN(net3662),
    .CLK(clknet_leaf_263_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[415] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[416]$_DFFE_PN0P_  (.D(_00862_),
    .RN(net3662),
    .CLK(clknet_leaf_364_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[416] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[417]$_DFFE_PN0P_  (.D(_00863_),
    .RN(net3661),
    .CLK(clknet_leaf_537_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[417] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[418]$_DFFE_PN0P_  (.D(_00864_),
    .RN(net3662),
    .CLK(clknet_leaf_258_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[418] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[419]$_DFFE_PN0P_  (.D(_00865_),
    .RN(net3662),
    .CLK(clknet_leaf_251_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[419] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[41]$_DFFE_PN0P_  (.D(_00866_),
    .RN(net3661),
    .CLK(clknet_6_19__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[420]$_DFFE_PN0P_  (.D(_00867_),
    .RN(net3662),
    .CLK(clknet_6_38__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[420] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[421]$_DFFE_PN0P_  (.D(_00868_),
    .RN(net3662),
    .CLK(clknet_leaf_462_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[421] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[422]$_DFFE_PN0P_  (.D(_00869_),
    .RN(net3661),
    .CLK(clknet_leaf_478_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[422] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[423]$_DFFE_PN0P_  (.D(_00870_),
    .RN(net3661),
    .CLK(clknet_6_28__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[423] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[424]$_DFFE_PN0P_  (.D(_00871_),
    .RN(net3661),
    .CLK(clknet_leaf_514_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[424] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[425]$_DFFE_PN0P_  (.D(_00872_),
    .RN(net3661),
    .CLK(clknet_6_19__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[425] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[426]$_DFFE_PN0P_  (.D(_00873_),
    .RN(net3661),
    .CLK(clknet_leaf_512_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[426] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[427]$_DFFE_PN0P_  (.D(_00874_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[427] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[428]$_DFFE_PN0P_  (.D(_00875_),
    .RN(net3663),
    .CLK(clknet_6_56__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[428] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[429]$_DFFE_PN0P_  (.D(_00876_),
    .RN(net3663),
    .CLK(clknet_6_56__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[429] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[42]$_DFFE_PN0P_  (.D(_00877_),
    .RN(net3661),
    .CLK(clknet_6_26__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[430]$_DFFE_PN0P_  (.D(_00878_),
    .RN(net3661),
    .CLK(clknet_leaf_409_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[430] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[431]$_DFFE_PN0P_  (.D(_00879_),
    .RN(net3662),
    .CLK(clknet_leaf_376_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[431] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[432]$_DFFE_PN0P_  (.D(_00880_),
    .RN(net3662),
    .CLK(clknet_6_10__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[432] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[433]$_DFFE_PN0P_  (.D(_00881_),
    .RN(net3662),
    .CLK(clknet_leaf_440_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[433] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[434]$_DFFE_PN0P_  (.D(_00882_),
    .RN(net3663),
    .CLK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[434] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[435]$_DFFE_PN0P_  (.D(_00883_),
    .RN(net3662),
    .CLK(clknet_leaf_269_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[435] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[436]$_DFFE_PN0P_  (.D(_00884_),
    .RN(net3663),
    .CLK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[436] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[437]$_DFFE_PN0P_  (.D(_00885_),
    .RN(net3662),
    .CLK(clknet_leaf_265_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[437] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[438]$_DFFE_PN0P_  (.D(_00886_),
    .RN(net3662),
    .CLK(clknet_leaf_309_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[438] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[439]$_DFFE_PN0P_  (.D(_00887_),
    .RN(net3661),
    .CLK(clknet_leaf_404_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[439] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[43]$_DFFE_PN0P_  (.D(_00888_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[440]$_DFFE_PN0P_  (.D(_00889_),
    .RN(net3662),
    .CLK(clknet_leaf_378_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[440] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[441]$_DFFE_PN0P_  (.D(_00890_),
    .RN(net3663),
    .CLK(clknet_leaf_183_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[441] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[442]$_DFFE_PN0P_  (.D(_00891_),
    .RN(net3663),
    .CLK(clknet_leaf_200_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[442] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[443]$_DFFE_PN0P_  (.D(_00892_),
    .RN(net3663),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[443] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[444]$_DFFE_PN0P_  (.D(_00893_),
    .RN(net3663),
    .CLK(clknet_6_54__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[444] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[445]$_DFFE_PN0P_  (.D(_00894_),
    .RN(net3663),
    .CLK(clknet_leaf_42_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[445] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[446]$_DFFE_PN0P_  (.D(_00895_),
    .RN(net3663),
    .CLK(clknet_leaf_98_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[446] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[447]$_DFFE_PN0P_  (.D(_00896_),
    .RN(net3662),
    .CLK(clknet_leaf_263_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[447] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[448]$_DFFE_PN0P_  (.D(_00897_),
    .RN(net3662),
    .CLK(clknet_6_9__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[448] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[449]$_DFFE_PN0P_  (.D(_00898_),
    .RN(net3661),
    .CLK(clknet_leaf_537_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[449] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[44]$_DFFE_PN0P_  (.D(_00899_),
    .RN(net3663),
    .CLK(clknet_leaf_154_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[450]$_DFFE_PN0P_  (.D(_00900_),
    .RN(net3662),
    .CLK(clknet_leaf_262_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[450] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[451]$_DFFE_PN0P_  (.D(_00901_),
    .RN(net3662),
    .CLK(clknet_leaf_251_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[451] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[452]$_DFFE_PN0P_  (.D(_00902_),
    .RN(net3662),
    .CLK(clknet_6_31__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[452] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[453]$_DFFE_PN0P_  (.D(_00903_),
    .RN(net3662),
    .CLK(clknet_leaf_453_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[453] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[454]$_DFFE_PN0P_  (.D(_00904_),
    .RN(net3661),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[454] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[455]$_DFFE_PN0P_  (.D(_00905_),
    .RN(net3661),
    .CLK(clknet_leaf_480_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[455] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[456]$_DFFE_PN0P_  (.D(_00906_),
    .RN(net3661),
    .CLK(clknet_leaf_517_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[456] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[457]$_DFFE_PN0P_  (.D(_00907_),
    .RN(net3661),
    .CLK(clknet_leaf_522_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[457] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[458]$_DFFE_PN0P_  (.D(_00908_),
    .RN(net3661),
    .CLK(clknet_leaf_512_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[458] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[459]$_DFFE_PN0P_  (.D(_00909_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[459] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[45]$_DFFE_PN0P_  (.D(_00910_),
    .RN(net3663),
    .CLK(clknet_leaf_112_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[460]$_DFFE_PN0P_  (.D(_00911_),
    .RN(net3663),
    .CLK(clknet_6_45__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[460] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[461]$_DFFE_PN0P_  (.D(_00912_),
    .RN(net3663),
    .CLK(clknet_6_56__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[461] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[462]$_DFFE_PN0P_  (.D(_00913_),
    .RN(net3661),
    .CLK(clknet_leaf_409_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[462] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[463]$_DFFE_PN0P_  (.D(_00914_),
    .RN(net3662),
    .CLK(clknet_leaf_373_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[463] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[464]$_DFFE_PN0P_  (.D(_00915_),
    .RN(net3662),
    .CLK(clknet_leaf_350_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[464] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[465]$_DFFE_PN0P_  (.D(_00916_),
    .RN(net3662),
    .CLK(clknet_leaf_449_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[465] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[466]$_DFFE_PN0P_  (.D(_00917_),
    .RN(net3663),
    .CLK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[466] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[467]$_DFFE_PN0P_  (.D(_00918_),
    .RN(net3662),
    .CLK(clknet_6_41__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[467] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[468]$_DFFE_PN0P_  (.D(_00919_),
    .RN(net3663),
    .CLK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[468] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[469]$_DFFE_PN0P_  (.D(_00920_),
    .RN(net3662),
    .CLK(clknet_leaf_264_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[469] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[46]$_DFFE_PN0P_  (.D(_00921_),
    .RN(net3662),
    .CLK(clknet_6_3__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[470]$_DFFE_PN0P_  (.D(_00922_),
    .RN(net3662),
    .CLK(clknet_leaf_311_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[470] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[471]$_DFFE_PN0P_  (.D(_00923_),
    .RN(net3661),
    .CLK(clknet_leaf_518_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[471] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[472]$_DFFE_PN0P_  (.D(_00924_),
    .RN(net3662),
    .CLK(clknet_leaf_375_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[472] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[473]$_DFFE_PN0P_  (.D(_00925_),
    .RN(net3663),
    .CLK(clknet_leaf_183_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[473] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[474]$_DFFE_PN0P_  (.D(_00926_),
    .RN(net3663),
    .CLK(clknet_leaf_205_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[474] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[475]$_DFFE_PN0P_  (.D(_00927_),
    .RN(net3663),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[475] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[476]$_DFFE_PN0P_  (.D(_00928_),
    .RN(net3663),
    .CLK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[476] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[477]$_DFFE_PN0P_  (.D(_00929_),
    .RN(net3663),
    .CLK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[477] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[478]$_DFFE_PN0P_  (.D(_00930_),
    .RN(net3663),
    .CLK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[478] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[479]$_DFFE_PN0P_  (.D(_00931_),
    .RN(net3662),
    .CLK(clknet_leaf_233_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[479] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[47]$_DFFE_PN0P_  (.D(_00932_),
    .RN(net3662),
    .CLK(clknet_6_3__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[480]$_DFFE_PN0P_  (.D(_00933_),
    .RN(net3662),
    .CLK(clknet_leaf_364_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[480] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[481]$_DFFE_PN0P_  (.D(_00934_),
    .RN(net3661),
    .CLK(clknet_leaf_537_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[481] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[482]$_DFFE_PN0P_  (.D(_00935_),
    .RN(net3662),
    .CLK(clknet_leaf_262_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[482] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[483]$_DFFE_PN0P_  (.D(_00936_),
    .RN(net3662),
    .CLK(clknet_6_13__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[483] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[484]$_DFFE_PN0P_  (.D(_00937_),
    .RN(net3662),
    .CLK(clknet_6_31__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[484] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[485]$_DFFE_PN0P_  (.D(_00938_),
    .RN(net3662),
    .CLK(clknet_leaf_453_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[485] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[486]$_DFFE_PN0P_  (.D(_00939_),
    .RN(net3661),
    .CLK(clknet_6_29__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[486] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[487]$_DFFE_PN0P_  (.D(_00940_),
    .RN(net3661),
    .CLK(clknet_leaf_480_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[487] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[488]$_DFFE_PN0P_  (.D(_00941_),
    .RN(net3661),
    .CLK(clknet_leaf_517_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[488] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[489]$_DFFE_PN0P_  (.D(_00942_),
    .RN(net3661),
    .CLK(clknet_leaf_522_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[489] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[48]$_DFFE_PN0P_  (.D(_00943_),
    .RN(net3662),
    .CLK(clknet_leaf_320_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[490]$_DFFE_PN0P_  (.D(_00944_),
    .RN(net3661),
    .CLK(clknet_leaf_510_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[490] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[491]$_DFFE_PN0P_  (.D(_00945_),
    .RN(net3663),
    .CLK(clknet_leaf_473_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[491] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[492]$_DFFE_PN0P_  (.D(_00946_),
    .RN(net3663),
    .CLK(clknet_leaf_169_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[492] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[493]$_DFFE_PN0P_  (.D(_00947_),
    .RN(net3663),
    .CLK(clknet_leaf_171_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[493] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[494]$_DFFE_PN0P_  (.D(_00948_),
    .RN(net3661),
    .CLK(clknet_leaf_408_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[494] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[495]$_DFFE_PN0P_  (.D(_00949_),
    .RN(net3662),
    .CLK(clknet_leaf_373_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[495] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[496]$_DFFE_PN0P_  (.D(_00950_),
    .RN(net3662),
    .CLK(clknet_leaf_350_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[496] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[497]$_DFFE_PN0P_  (.D(_00951_),
    .RN(net3662),
    .CLK(clknet_leaf_449_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[497] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[498]$_DFFE_PN0P_  (.D(_00952_),
    .RN(net3663),
    .CLK(clknet_leaf_101_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[498] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[499]$_DFFE_PN0P_  (.D(_00953_),
    .RN(net3662),
    .CLK(clknet_6_41__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[499] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[49]$_DFFE_PN0P_  (.D(_00954_),
    .RN(net3662),
    .CLK(clknet_leaf_241_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[500]$_DFFE_PN0P_  (.D(_00955_),
    .RN(net3663),
    .CLK(clknet_leaf_97_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[500] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[501]$_DFFE_PN0P_  (.D(_00956_),
    .RN(net3662),
    .CLK(clknet_leaf_264_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[501] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[502]$_DFFE_PN0P_  (.D(_00957_),
    .RN(net3662),
    .CLK(clknet_leaf_311_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[502] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[503]$_DFFE_PN0P_  (.D(_00958_),
    .RN(net3661),
    .CLK(clknet_6_25__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[503] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[504]$_DFFE_PN0P_  (.D(_00959_),
    .RN(net3662),
    .CLK(clknet_leaf_378_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[504] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[505]$_DFFE_PN0P_  (.D(_00960_),
    .RN(net3663),
    .CLK(clknet_6_50__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[505] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[506]$_DFFE_PN0P_  (.D(_00961_),
    .RN(net3663),
    .CLK(clknet_6_39__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[506] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[507]$_DFFE_PN0P_  (.D(_00962_),
    .RN(net3663),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[507] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[508]$_DFFE_PN0P_  (.D(_00963_),
    .RN(net3663),
    .CLK(clknet_leaf_104_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[508] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[509]$_DFFE_PN0P_  (.D(_00964_),
    .RN(net3663),
    .CLK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[509] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[50]$_DFFE_PN0P_  (.D(_00965_),
    .RN(net3663),
    .CLK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[510]$_DFFE_PN0P_  (.D(_00966_),
    .RN(net3663),
    .CLK(clknet_leaf_44_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[510] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[511]$_DFFE_PN0P_  (.D(_00967_),
    .RN(net3662),
    .CLK(clknet_leaf_233_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[511] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[512]$_DFFE_PN0P_  (.D(_00968_),
    .RN(net3662),
    .CLK(clknet_leaf_356_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[512] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[513]$_DFFE_PN0P_  (.D(_00969_),
    .RN(net3661),
    .CLK(clknet_6_18__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[513] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[514]$_DFFE_PN0P_  (.D(_00970_),
    .RN(net3662),
    .CLK(clknet_leaf_294_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[514] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[515]$_DFFE_PN0P_  (.D(_00971_),
    .RN(net3662),
    .CLK(clknet_leaf_295_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[515] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[516]$_DFFE_PN0P_  (.D(_00972_),
    .RN(net3662),
    .CLK(clknet_6_33__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[516] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[517]$_DFFE_PN0P_  (.D(_00973_),
    .RN(net3661),
    .CLK(clknet_leaf_419_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[517] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[518]$_DFFE_PN0P_  (.D(_00974_),
    .RN(net3661),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[518] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[519]$_DFFE_PN0P_  (.D(_00975_),
    .RN(net3661),
    .CLK(clknet_leaf_494_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[519] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[51]$_DFFE_PN0P_  (.D(_00976_),
    .RN(net3663),
    .CLK(clknet_leaf_147_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[520]$_DFFE_PN0P_  (.D(_00977_),
    .RN(net3661),
    .CLK(clknet_6_17__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[520] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[521]$_DFFE_PN0P_  (.D(_00978_),
    .RN(net3661),
    .CLK(clknet_6_19__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[521] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[522]$_DFFE_PN0P_  (.D(_00979_),
    .RN(net3661),
    .CLK(clknet_leaf_512_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[522] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[523]$_DFFE_PN0P_  (.D(_00980_),
    .RN(net3663),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[523] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[524]$_DFFE_PN0P_  (.D(_00981_),
    .RN(net3663),
    .CLK(clknet_leaf_143_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[524] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[525]$_DFFE_PN0P_  (.D(_00982_),
    .RN(net3663),
    .CLK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[525] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[526]$_DFFE_PN0P_  (.D(_00983_),
    .RN(net3661),
    .CLK(clknet_leaf_397_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[526] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[527]$_DFFE_PN0P_  (.D(_00984_),
    .RN(net3662),
    .CLK(clknet_leaf_385_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[527] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[528]$_DFFE_PN0P_  (.D(_00985_),
    .RN(net3662),
    .CLK(clknet_6_11__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[528] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[529]$_DFFE_PN0P_  (.D(_00986_),
    .RN(net3662),
    .CLK(clknet_leaf_436_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[529] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[52]$_DFFE_PN0P_  (.D(_00987_),
    .RN(net3664),
    .CLK(clknet_leaf_95_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[530]$_DFFE_PN0P_  (.D(_00988_),
    .RN(net3664),
    .CLK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[530] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[531]$_DFFE_PN0P_  (.D(_00989_),
    .RN(net3662),
    .CLK(clknet_leaf_283_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[531] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[532]$_DFFE_PN0P_  (.D(_00990_),
    .RN(net3664),
    .CLK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[532] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[533]$_DFFE_PN0P_  (.D(_00991_),
    .RN(net3663),
    .CLK(clknet_6_34__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[533] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[534]$_DFFE_PN0P_  (.D(_00992_),
    .RN(net3662),
    .CLK(clknet_6_14__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[534] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[535]$_DFFE_PN0P_  (.D(_00993_),
    .RN(net3661),
    .CLK(clknet_leaf_400_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[535] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[536]$_DFFE_PN0P_  (.D(_00994_),
    .RN(net3662),
    .CLK(clknet_leaf_348_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[536] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[537]$_DFFE_PN0P_  (.D(_00995_),
    .RN(net3663),
    .CLK(clknet_leaf_178_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[537] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[538]$_DFFE_PN0P_  (.D(_00996_),
    .RN(net3663),
    .CLK(clknet_6_50__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[538] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[539]$_DFFE_PN0P_  (.D(_00997_),
    .RN(net3663),
    .CLK(clknet_leaf_34_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[539] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[53]$_DFFE_PN0P_  (.D(_00998_),
    .RN(net3662),
    .CLK(clknet_leaf_266_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[540]$_DFFE_PN0P_  (.D(_00999_),
    .RN(net3663),
    .CLK(clknet_6_61__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[540] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[541]$_DFFE_PN0P_  (.D(_01000_),
    .RN(net3663),
    .CLK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[541] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[542]$_DFFE_PN0P_  (.D(_01001_),
    .RN(net3663),
    .CLK(clknet_6_63__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[542] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[543]$_DFFE_PN0P_  (.D(_01002_),
    .RN(net3662),
    .CLK(clknet_leaf_244_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[543] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[544]$_DFFE_PN0P_  (.D(_01003_),
    .RN(net3662),
    .CLK(clknet_6_9__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[544] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[545]$_DFFE_PN0P_  (.D(_01004_),
    .RN(net3661),
    .CLK(clknet_leaf_543_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[545] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[546]$_DFFE_PN0P_  (.D(_01005_),
    .RN(net3662),
    .CLK(clknet_leaf_287_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[546] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[547]$_DFFE_PN0P_  (.D(_01006_),
    .RN(net3662),
    .CLK(clknet_leaf_295_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[547] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[548]$_DFFE_PN0P_  (.D(_01007_),
    .RN(net3662),
    .CLK(clknet_leaf_237_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[548] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[549]$_DFFE_PN0P_  (.D(_01008_),
    .RN(net3661),
    .CLK(clknet_leaf_417_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[549] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[54]$_DFFE_PN0P_  (.D(_01009_),
    .RN(net3662),
    .CLK(clknet_6_12__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[550]$_DFFE_PN0P_  (.D(_01010_),
    .RN(net3661),
    .CLK(clknet_6_29__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[550] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[551]$_DFFE_PN0P_  (.D(_01011_),
    .RN(net3661),
    .CLK(clknet_leaf_495_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[551] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[552]$_DFFE_PN0P_  (.D(_01012_),
    .RN(net3661),
    .CLK(clknet_6_16__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[552] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[553]$_DFFE_PN0P_  (.D(_01013_),
    .RN(net3661),
    .CLK(clknet_leaf_507_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[553] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[554]$_DFFE_PN0P_  (.D(_01014_),
    .RN(net3661),
    .CLK(clknet_6_21__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[554] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[555]$_DFFE_PN0P_  (.D(_01015_),
    .RN(net3663),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[555] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[556]$_DFFE_PN0P_  (.D(_01016_),
    .RN(net3663),
    .CLK(clknet_leaf_143_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[556] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[557]$_DFFE_PN0P_  (.D(_01017_),
    .RN(net3663),
    .CLK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[557] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[558]$_DFFE_PN0P_  (.D(_01018_),
    .RN(net3661),
    .CLK(clknet_leaf_397_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[558] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[559]$_DFFE_PN0P_  (.D(_01019_),
    .RN(net3662),
    .CLK(clknet_leaf_384_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[559] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[55]$_DFFE_PN0P_  (.D(_01020_),
    .RN(net3661),
    .CLK(clknet_6_1__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[560]$_DFFE_PN0P_  (.D(_01021_),
    .RN(net3662),
    .CLK(clknet_leaf_330_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[560] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[561]$_DFFE_PN0P_  (.D(_01022_),
    .RN(net3662),
    .CLK(clknet_leaf_435_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[561] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[562]$_DFFE_PN0P_  (.D(_01023_),
    .RN(net3664),
    .CLK(clknet_leaf_125_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[562] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[563]$_DFFE_PN0P_  (.D(_01024_),
    .RN(net3662),
    .CLK(clknet_6_46__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[563] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[564]$_DFFE_PN0P_  (.D(_01025_),
    .RN(net3664),
    .CLK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[564] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[565]$_DFFE_PN0P_  (.D(_01026_),
    .RN(net3663),
    .CLK(clknet_leaf_231_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[565] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[566]$_DFFE_PN0P_  (.D(_01027_),
    .RN(net3662),
    .CLK(clknet_6_14__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[566] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[567]$_DFFE_PN0P_  (.D(_01028_),
    .RN(net3661),
    .CLK(clknet_leaf_400_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[567] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[568]$_DFFE_PN0P_  (.D(_01029_),
    .RN(net3662),
    .CLK(clknet_leaf_349_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[568] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[569]$_DFFE_PN0P_  (.D(_01030_),
    .RN(net3663),
    .CLK(clknet_leaf_178_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[569] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[56]$_DFFE_PN0P_  (.D(_01031_),
    .RN(net3662),
    .CLK(clknet_leaf_359_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[570]$_DFFE_PN0P_  (.D(_01032_),
    .RN(net3663),
    .CLK(clknet_6_50__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[570] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[571]$_DFFE_PN0P_  (.D(_01033_),
    .RN(net3663),
    .CLK(clknet_leaf_35_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[571] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[572]$_DFFE_PN0P_  (.D(_01034_),
    .RN(net3663),
    .CLK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[572] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[573]$_DFFE_PN0P_  (.D(_01035_),
    .RN(net3663),
    .CLK(clknet_6_55__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[573] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[574]$_DFFE_PN0P_  (.D(_01036_),
    .RN(net3663),
    .CLK(clknet_6_63__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[574] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[575]$_DFFE_PN0P_  (.D(_01037_),
    .RN(net3662),
    .CLK(clknet_leaf_244_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[575] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[576]$_DFFE_PN0P_  (.D(_01038_),
    .RN(net3662),
    .CLK(clknet_leaf_359_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[576] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[577]$_DFFE_PN0P_  (.D(_01039_),
    .RN(net3661),
    .CLK(clknet_leaf_543_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[577] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[578]$_DFFE_PN0P_  (.D(_01040_),
    .RN(net3662),
    .CLK(clknet_leaf_288_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[578] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[579]$_DFFE_PN0P_  (.D(_01041_),
    .RN(net3662),
    .CLK(clknet_leaf_302_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[579] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[57]$_DFFE_PN0P_  (.D(_01042_),
    .RN(net3663),
    .CLK(clknet_6_50__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[580]$_DFFE_PN0P_  (.D(_01043_),
    .RN(net3662),
    .CLK(clknet_leaf_222_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[580] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[581]$_DFFE_PN0P_  (.D(_01044_),
    .RN(net3661),
    .CLK(clknet_leaf_418_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[581] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[582]$_DFFE_PN0P_  (.D(_01045_),
    .RN(net3661),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[582] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[583]$_DFFE_PN0P_  (.D(_01046_),
    .RN(net3661),
    .CLK(clknet_leaf_494_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[583] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[584]$_DFFE_PN0P_  (.D(_01047_),
    .RN(net3661),
    .CLK(clknet_leaf_556_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[584] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[585]$_DFFE_PN0P_  (.D(_01048_),
    .RN(net3661),
    .CLK(clknet_leaf_557_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[585] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[586]$_DFFE_PN0P_  (.D(_01049_),
    .RN(net3661),
    .CLK(clknet_6_22__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[586] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[587]$_DFFE_PN0P_  (.D(_01050_),
    .RN(net3663),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[587] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[588]$_DFFE_PN0P_  (.D(_01051_),
    .RN(net3663),
    .CLK(clknet_leaf_142_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[588] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[589]$_DFFE_PN0P_  (.D(_01052_),
    .RN(net3663),
    .CLK(clknet_leaf_127_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[589] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[58]$_DFFE_PN0P_  (.D(_01053_),
    .RN(net3663),
    .CLK(clknet_leaf_201_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[590]$_DFFE_PN0P_  (.D(_01054_),
    .RN(net3661),
    .CLK(clknet_leaf_397_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[590] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[591]$_DFFE_PN0P_  (.D(_01055_),
    .RN(net3662),
    .CLK(clknet_leaf_384_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[591] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[592]$_DFFE_PN0P_  (.D(_01056_),
    .RN(net3662),
    .CLK(clknet_leaf_335_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[592] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[593]$_DFFE_PN0P_  (.D(_01057_),
    .RN(net3662),
    .CLK(clknet_6_6__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[593] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[594]$_DFFE_PN0P_  (.D(_01058_),
    .RN(net3664),
    .CLK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[594] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[595]$_DFFE_PN0P_  (.D(_01059_),
    .RN(net3663),
    .CLK(clknet_leaf_282_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[595] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[596]$_DFFE_PN0P_  (.D(_01060_),
    .RN(net3664),
    .CLK(clknet_6_62__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[596] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[597]$_DFFE_PN0P_  (.D(_01061_),
    .RN(net3663),
    .CLK(clknet_leaf_230_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[597] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[598]$_DFFE_PN0P_  (.D(_01062_),
    .RN(net3662),
    .CLK(clknet_leaf_327_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[598] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[599]$_DFFE_PN0P_  (.D(_01063_),
    .RN(net3661),
    .CLK(clknet_leaf_532_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[599] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[59]$_DFFE_PN0P_  (.D(_01064_),
    .RN(net3663),
    .CLK(clknet_6_51__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[600]$_DFFE_PN0P_  (.D(_01065_),
    .RN(net3662),
    .CLK(clknet_6_8__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[600] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[601]$_DFFE_PN0P_  (.D(_01066_),
    .RN(net3663),
    .CLK(clknet_leaf_179_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[601] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[602]$_DFFE_PN0P_  (.D(_01067_),
    .RN(net3663),
    .CLK(clknet_leaf_186_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[602] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[603]$_DFFE_PN0P_  (.D(_01068_),
    .RN(net3663),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[603] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[604]$_DFFE_PN0P_  (.D(_01069_),
    .RN(net3663),
    .CLK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[604] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[605]$_DFFE_PN0P_  (.D(_01070_),
    .RN(net3663),
    .CLK(clknet_6_53__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[605] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[606]$_DFFE_PN0P_  (.D(_01071_),
    .RN(net3663),
    .CLK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[606] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[607]$_DFFE_PN0P_  (.D(_01072_),
    .RN(net3662),
    .CLK(clknet_6_13__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[607] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[608]$_DFFE_PN0P_  (.D(_01073_),
    .RN(net3662),
    .CLK(clknet_6_9__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[608] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[609]$_DFFE_PN0P_  (.D(_01074_),
    .RN(net3661),
    .CLK(clknet_leaf_544_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[609] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[60]$_DFFE_PN0P_  (.D(_01075_),
    .RN(net3663),
    .CLK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[610]$_DFFE_PN0P_  (.D(_01076_),
    .RN(net3662),
    .CLK(clknet_leaf_294_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[610] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[611]$_DFFE_PN0P_  (.D(_01077_),
    .RN(net3662),
    .CLK(clknet_6_15__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[611] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[612]$_DFFE_PN0P_  (.D(_01078_),
    .RN(net3662),
    .CLK(clknet_leaf_222_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[612] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[613]$_DFFE_PN0P_  (.D(_01079_),
    .RN(net3661),
    .CLK(clknet_6_26__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[613] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[614]$_DFFE_PN0P_  (.D(_01080_),
    .RN(net3661),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[614] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[615]$_DFFE_PN0P_  (.D(_01081_),
    .RN(net3661),
    .CLK(clknet_leaf_495_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[615] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[616]$_DFFE_PN0P_  (.D(_01082_),
    .RN(net3661),
    .CLK(clknet_leaf_556_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[616] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[617]$_DFFE_PN0P_  (.D(_01083_),
    .RN(net3661),
    .CLK(clknet_leaf_507_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[617] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[618]$_DFFE_PN0P_  (.D(_01084_),
    .RN(net3661),
    .CLK(clknet_6_21__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[618] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[619]$_DFFE_PN0P_  (.D(_01085_),
    .RN(net3663),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[619] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[61]$_DFFE_PN0P_  (.D(_01086_),
    .RN(net3663),
    .CLK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[620]$_DFFE_PN0P_  (.D(_01087_),
    .RN(net3663),
    .CLK(clknet_leaf_142_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[620] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[621]$_DFFE_PN0P_  (.D(_01088_),
    .RN(net3663),
    .CLK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[621] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[622]$_DFFE_PN0P_  (.D(_01089_),
    .RN(net3661),
    .CLK(clknet_leaf_398_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[622] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[623]$_DFFE_PN0P_  (.D(_01090_),
    .RN(net3662),
    .CLK(clknet_leaf_381_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[623] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[624]$_DFFE_PN0P_  (.D(_01091_),
    .RN(net3662),
    .CLK(clknet_leaf_330_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[624] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[625]$_DFFE_PN0P_  (.D(_01092_),
    .RN(net3662),
    .CLK(clknet_leaf_435_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[625] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[626]$_DFFE_PN0P_  (.D(_01093_),
    .RN(net3664),
    .CLK(clknet_leaf_124_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[626] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[627]$_DFFE_PN0P_  (.D(_01094_),
    .RN(net3663),
    .CLK(clknet_leaf_282_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[627] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[628]$_DFFE_PN0P_  (.D(_01095_),
    .RN(net3664),
    .CLK(clknet_leaf_74_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[628] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[629]$_DFFE_PN0P_  (.D(_01096_),
    .RN(net3663),
    .CLK(clknet_leaf_230_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[629] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[62]$_DFFE_PN0P_  (.D(_01097_),
    .RN(net3663),
    .CLK(clknet_6_60__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[630]$_DFFE_PN0P_  (.D(_01098_),
    .RN(net3662),
    .CLK(clknet_leaf_327_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[630] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[631]$_DFFE_PN0P_  (.D(_01099_),
    .RN(net3661),
    .CLK(clknet_leaf_532_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[631] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[632]$_DFFE_PN0P_  (.D(_01100_),
    .RN(net3662),
    .CLK(clknet_leaf_348_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[632] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[633]$_DFFE_PN0P_  (.D(_01101_),
    .RN(net3663),
    .CLK(clknet_leaf_179_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[633] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[634]$_DFFE_PN0P_  (.D(_01102_),
    .RN(net3663),
    .CLK(clknet_leaf_187_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[634] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[635]$_DFFE_PN0P_  (.D(_01103_),
    .RN(net3663),
    .CLK(clknet_6_52__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[635] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[636]$_DFFE_PN0P_  (.D(_01104_),
    .RN(net3663),
    .CLK(clknet_6_61__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[636] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[637]$_DFFE_PN0P_  (.D(_01105_),
    .RN(net3663),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[637] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[638]$_DFFE_PN0P_  (.D(_01106_),
    .RN(net3663),
    .CLK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[638] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[639]$_DFFE_PN0P_  (.D(_01107_),
    .RN(net3662),
    .CLK(clknet_leaf_252_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[639] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[63]$_DFFE_PN0P_  (.D(_01108_),
    .RN(net3662),
    .CLK(clknet_leaf_237_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[640]$_DFFE_PN0P_  (.D(_01109_),
    .RN(net3662),
    .CLK(clknet_6_10__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[640] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[641]$_DFFE_PN0P_  (.D(_01110_),
    .RN(net3661),
    .CLK(clknet_leaf_540_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[641] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[642]$_DFFE_PN0P_  (.D(_01111_),
    .RN(net3662),
    .CLK(clknet_leaf_287_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[642] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[643]$_DFFE_PN0P_  (.D(_01112_),
    .RN(net3662),
    .CLK(clknet_6_42__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[643] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[644]$_DFFE_PN0P_  (.D(_01113_),
    .RN(net3662),
    .CLK(clknet_6_33__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[644] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[645]$_DFFE_PN0P_  (.D(_01114_),
    .RN(net3661),
    .CLK(clknet_6_27__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[645] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[646]$_DFFE_PN0P_  (.D(_01115_),
    .RN(net3661),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[646] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[647]$_DFFE_PN0P_  (.D(_01116_),
    .RN(net3661),
    .CLK(clknet_leaf_497_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[647] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[648]$_DFFE_PN0P_  (.D(_01117_),
    .RN(net3661),
    .CLK(clknet_leaf_540_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[648] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[649]$_DFFE_PN0P_  (.D(_01118_),
    .RN(net3661),
    .CLK(clknet_leaf_507_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[649] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[64]$_DFFE_PN0P_  (.D(_01119_),
    .RN(net3662),
    .CLK(clknet_leaf_436_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[64] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[650]$_DFFE_PN0P_  (.D(_01120_),
    .RN(net3661),
    .CLK(clknet_leaf_497_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[650] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[651]$_DFFE_PN0P_  (.D(_01121_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[651] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[652]$_DFFE_PN0P_  (.D(_01122_),
    .RN(net3663),
    .CLK(clknet_leaf_141_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[652] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[653]$_DFFE_PN0P_  (.D(_01123_),
    .RN(net3663),
    .CLK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[653] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[654]$_DFFE_PN0P_  (.D(_01124_),
    .RN(net3661),
    .CLK(clknet_6_0__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[654] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[655]$_DFFE_PN0P_  (.D(_01125_),
    .RN(net3662),
    .CLK(clknet_6_2__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[655] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[656]$_DFFE_PN0P_  (.D(_01126_),
    .RN(net3662),
    .CLK(clknet_leaf_331_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[656] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[657]$_DFFE_PN0P_  (.D(_01127_),
    .RN(net3662),
    .CLK(clknet_leaf_247_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[657] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[658]$_DFFE_PN0P_  (.D(_01128_),
    .RN(net3664),
    .CLK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[658] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[659]$_DFFE_PN0P_  (.D(_01129_),
    .RN(net3662),
    .CLK(clknet_leaf_283_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[659] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[65]$_DFFE_PN0P_  (.D(_01130_),
    .RN(net3661),
    .CLK(clknet_leaf_535_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[65] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[660]$_DFFE_PN0P_  (.D(_01131_),
    .RN(net3664),
    .CLK(clknet_6_62__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[660] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[661]$_DFFE_PN0P_  (.D(_01132_),
    .RN(net3663),
    .CLK(clknet_leaf_231_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[661] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[662]$_DFFE_PN0P_  (.D(_01133_),
    .RN(net3662),
    .CLK(clknet_leaf_296_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[662] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[663]$_DFFE_PN0P_  (.D(_01134_),
    .RN(net3661),
    .CLK(clknet_leaf_398_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[663] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[664]$_DFFE_PN0P_  (.D(_01135_),
    .RN(net3662),
    .CLK(clknet_leaf_342_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[664] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[665]$_DFFE_PN0P_  (.D(_01136_),
    .RN(net3663),
    .CLK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[665] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[666]$_DFFE_PN0P_  (.D(_01137_),
    .RN(net3663),
    .CLK(clknet_leaf_180_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[666] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[667]$_DFFE_PN0P_  (.D(_01138_),
    .RN(net3663),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[667] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[668]$_DFFE_PN0P_  (.D(_01139_),
    .RN(net3663),
    .CLK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[668] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[669]$_DFFE_PN0P_  (.D(_01140_),
    .RN(net3663),
    .CLK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[669] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[66]$_DFFE_PN0P_  (.D(_01141_),
    .RN(net3662),
    .CLK(clknet_6_40__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[66] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[670]$_DFFE_PN0P_  (.D(_01142_),
    .RN(net3663),
    .CLK(clknet_6_63__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[670] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[671]$_DFFE_PN0P_  (.D(_01143_),
    .RN(net3662),
    .CLK(clknet_6_32__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[671] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[672]$_DFFE_PN0P_  (.D(_01144_),
    .RN(net3662),
    .CLK(clknet_6_10__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[672] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[673]$_DFFE_PN0P_  (.D(_01145_),
    .RN(net3661),
    .CLK(clknet_leaf_544_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[673] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[674]$_DFFE_PN0P_  (.D(_01146_),
    .RN(net3662),
    .CLK(clknet_leaf_287_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[674] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[675]$_DFFE_PN0P_  (.D(_01147_),
    .RN(net3662),
    .CLK(clknet_6_42__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[675] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[676]$_DFFE_PN0P_  (.D(_01148_),
    .RN(net3662),
    .CLK(clknet_6_5__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[676] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[677]$_DFFE_PN0P_  (.D(_01149_),
    .RN(net3661),
    .CLK(clknet_leaf_418_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[677] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[678]$_DFFE_PN0P_  (.D(_01150_),
    .RN(net3661),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[678] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[679]$_DFFE_PN0P_  (.D(_01151_),
    .RN(net3661),
    .CLK(clknet_leaf_498_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[679] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[67]$_DFFE_PN0P_  (.D(_01152_),
    .RN(net3662),
    .CLK(clknet_leaf_308_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[67] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[680]$_DFFE_PN0P_  (.D(_01153_),
    .RN(net3661),
    .CLK(clknet_6_17__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[680] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[681]$_DFFE_PN0P_  (.D(_01154_),
    .RN(net3661),
    .CLK(clknet_leaf_557_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[681] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[682]$_DFFE_PN0P_  (.D(_01155_),
    .RN(net3661),
    .CLK(clknet_leaf_503_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[682] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[683]$_DFFE_PN0P_  (.D(_01156_),
    .RN(net3663),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[683] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[684]$_DFFE_PN0P_  (.D(_01157_),
    .RN(net3663),
    .CLK(clknet_leaf_141_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[684] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[685]$_DFFE_PN0P_  (.D(_01158_),
    .RN(net3663),
    .CLK(clknet_6_58__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[685] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[686]$_DFFE_PN0P_  (.D(_01159_),
    .RN(net3661),
    .CLK(clknet_leaf_396_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[686] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[687]$_DFFE_PN0P_  (.D(_01160_),
    .RN(net3662),
    .CLK(clknet_leaf_381_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[687] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[688]$_DFFE_PN0P_  (.D(_01161_),
    .RN(net3662),
    .CLK(clknet_leaf_331_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[688] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[689]$_DFFE_PN0P_  (.D(_01162_),
    .RN(net3662),
    .CLK(clknet_6_7__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[689] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[68]$_DFFE_PN0P_  (.D(_01163_),
    .RN(net3662),
    .CLK(clknet_leaf_226_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[68] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[690]$_DFFE_PN0P_  (.D(_01164_),
    .RN(net3664),
    .CLK(clknet_leaf_87_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[690] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[691]$_DFFE_PN0P_  (.D(_01165_),
    .RN(net3662),
    .CLK(clknet_leaf_284_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[691] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[692]$_DFFE_PN0P_  (.D(_01166_),
    .RN(net3664),
    .CLK(clknet_leaf_84_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[692] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[693]$_DFFE_PN0P_  (.D(_01167_),
    .RN(net3663),
    .CLK(clknet_6_35__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[693] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[694]$_DFFE_PN0P_  (.D(_01168_),
    .RN(net3662),
    .CLK(clknet_leaf_296_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[694] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[695]$_DFFE_PN0P_  (.D(_01169_),
    .RN(net3661),
    .CLK(clknet_leaf_399_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[695] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[696]$_DFFE_PN0P_  (.D(_01170_),
    .RN(net3662),
    .CLK(clknet_leaf_342_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[696] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[697]$_DFFE_PN0P_  (.D(_01171_),
    .RN(net3663),
    .CLK(clknet_leaf_177_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[697] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[698]$_DFFE_PN0P_  (.D(_01172_),
    .RN(net3663),
    .CLK(clknet_leaf_180_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[698] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[699]$_DFFE_PN0P_  (.D(_01173_),
    .RN(net3663),
    .CLK(clknet_6_53__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[699] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[69]$_DFFE_PN0P_  (.D(_01174_),
    .RN(net3662),
    .CLK(clknet_leaf_450_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[69] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[700]$_DFFE_PN0P_  (.D(_01175_),
    .RN(net3663),
    .CLK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[700] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[701]$_DFFE_PN0P_  (.D(_01176_),
    .RN(net3663),
    .CLK(clknet_leaf_51_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[701] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[702]$_DFFE_PN0P_  (.D(_01177_),
    .RN(net3663),
    .CLK(clknet_leaf_62_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[702] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[703]$_DFFE_PN0P_  (.D(_01178_),
    .RN(net3662),
    .CLK(clknet_leaf_242_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[703] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[704]$_DFFE_PN0P_  (.D(_01179_),
    .RN(net3662),
    .CLK(clknet_leaf_356_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[704] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[705]$_DFFE_PN0P_  (.D(_01180_),
    .RN(net3661),
    .CLK(clknet_6_17__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[705] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[706]$_DFFE_PN0P_  (.D(_01181_),
    .RN(net3662),
    .CLK(clknet_leaf_288_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[706] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[707]$_DFFE_PN0P_  (.D(_01182_),
    .RN(net3662),
    .CLK(clknet_leaf_292_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[707] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[708]$_DFFE_PN0P_  (.D(_01183_),
    .RN(net3662),
    .CLK(clknet_6_5__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[708] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[709]$_DFFE_PN0P_  (.D(_01184_),
    .RN(net3661),
    .CLK(clknet_leaf_417_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[709] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[70]$_DFFE_PN0P_  (.D(_01185_),
    .RN(net3662),
    .CLK(clknet_leaf_476_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[70] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[710]$_DFFE_PN0P_  (.D(_01186_),
    .RN(net3661),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[710] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[711]$_DFFE_PN0P_  (.D(_01187_),
    .RN(net3661),
    .CLK(clknet_6_22__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[711] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[712]$_DFFE_PN0P_  (.D(_01188_),
    .RN(net3661),
    .CLK(clknet_leaf_556_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[712] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[713]$_DFFE_PN0P_  (.D(_01189_),
    .RN(net3661),
    .CLK(clknet_leaf_558_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[713] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[714]$_DFFE_PN0P_  (.D(_01190_),
    .RN(net3661),
    .CLK(clknet_leaf_503_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[714] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[715]$_DFFE_PN0P_  (.D(_01191_),
    .RN(net3663),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[715] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[716]$_DFFE_PN0P_  (.D(_01192_),
    .RN(net3663),
    .CLK(clknet_leaf_138_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[716] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[717]$_DFFE_PN0P_  (.D(_01193_),
    .RN(net3663),
    .CLK(clknet_leaf_139_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[717] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[718]$_DFFE_PN0P_  (.D(_01194_),
    .RN(net3661),
    .CLK(clknet_leaf_396_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[718] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[719]$_DFFE_PN0P_  (.D(_01195_),
    .RN(net3662),
    .CLK(clknet_leaf_383_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[719] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[71]$_DFFE_PN0P_  (.D(_01196_),
    .RN(net3661),
    .CLK(clknet_leaf_493_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[71] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[720]$_DFFE_PN0P_  (.D(_01197_),
    .RN(net3662),
    .CLK(clknet_leaf_332_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[720] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[721]$_DFFE_PN0P_  (.D(_01198_),
    .RN(net3662),
    .CLK(clknet_6_7__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[721] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[722]$_DFFE_PN0P_  (.D(_01199_),
    .RN(net3664),
    .CLK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[722] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[723]$_DFFE_PN0P_  (.D(_01200_),
    .RN(net3663),
    .CLK(clknet_leaf_286_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[723] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[724]$_DFFE_PN0P_  (.D(_01201_),
    .RN(net3664),
    .CLK(clknet_6_62__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[724] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[725]$_DFFE_PN0P_  (.D(_01202_),
    .RN(net3663),
    .CLK(clknet_leaf_196_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[725] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[726]$_DFFE_PN0P_  (.D(_01203_),
    .RN(net3662),
    .CLK(clknet_leaf_297_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[726] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[727]$_DFFE_PN0P_  (.D(_01204_),
    .RN(net3661),
    .CLK(clknet_6_24__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[727] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[728]$_DFFE_PN0P_  (.D(_01205_),
    .RN(net3662),
    .CLK(clknet_leaf_380_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[728] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[729]$_DFFE_PN0P_  (.D(_01206_),
    .RN(net3663),
    .CLK(clknet_leaf_178_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[729] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[72]$_DFFE_PN0P_  (.D(_01207_),
    .RN(net3661),
    .CLK(clknet_leaf_531_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[72] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[730]$_DFFE_PN0P_  (.D(_01208_),
    .RN(net3663),
    .CLK(clknet_6_51__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[730] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[731]$_DFFE_PN0P_  (.D(_01209_),
    .RN(net3663),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[731] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[732]$_DFFE_PN0P_  (.D(_01210_),
    .RN(net3663),
    .CLK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[732] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[733]$_DFFE_PN0P_  (.D(_01211_),
    .RN(net3663),
    .CLK(clknet_6_53__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[733] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[734]$_DFFE_PN0P_  (.D(_01212_),
    .RN(net3663),
    .CLK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[734] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[735]$_DFFE_PN0P_  (.D(_01213_),
    .RN(net3662),
    .CLK(clknet_leaf_242_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[735] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[736]$_DFFE_PN0P_  (.D(_01214_),
    .RN(net3662),
    .CLK(clknet_6_10__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[736] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[737]$_DFFE_PN0P_  (.D(_01215_),
    .RN(net3661),
    .CLK(clknet_6_16__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[737] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[738]$_DFFE_PN0P_  (.D(_01216_),
    .RN(net3662),
    .CLK(clknet_leaf_288_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[738] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[739]$_DFFE_PN0P_  (.D(_01217_),
    .RN(net3662),
    .CLK(clknet_leaf_292_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[739] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[73]$_DFFE_PN0P_  (.D(_01218_),
    .RN(net3661),
    .CLK(clknet_leaf_526_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[73] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[740]$_DFFE_PN0P_  (.D(_01219_),
    .RN(net3662),
    .CLK(clknet_6_5__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[740] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[741]$_DFFE_PN0P_  (.D(_01220_),
    .RN(net3661),
    .CLK(clknet_leaf_419_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[741] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[742]$_DFFE_PN0P_  (.D(_01221_),
    .RN(net3661),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[742] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[743]$_DFFE_PN0P_  (.D(_01222_),
    .RN(net3661),
    .CLK(clknet_leaf_498_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[743] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[744]$_DFFE_PN0P_  (.D(_01223_),
    .RN(net3661),
    .CLK(clknet_leaf_556_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[744] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[745]$_DFFE_PN0P_  (.D(_01224_),
    .RN(net3661),
    .CLK(clknet_leaf_558_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[745] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[746]$_DFFE_PN0P_  (.D(_01225_),
    .RN(net3661),
    .CLK(clknet_leaf_503_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[746] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[747]$_DFFE_PN0P_  (.D(_01226_),
    .RN(net3663),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[747] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[748]$_DFFE_PN0P_  (.D(_01227_),
    .RN(net3663),
    .CLK(clknet_leaf_138_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[748] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[749]$_DFFE_PN0P_  (.D(_01228_),
    .RN(net3663),
    .CLK(clknet_leaf_128_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[749] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[74]$_DFFE_PN0P_  (.D(_01229_),
    .RN(net3661),
    .CLK(clknet_6_28__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[74] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[750]$_DFFE_PN0P_  (.D(_01230_),
    .RN(net3661),
    .CLK(clknet_leaf_396_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[750] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[751]$_DFFE_PN0P_  (.D(_01231_),
    .RN(net3662),
    .CLK(clknet_leaf_383_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[751] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[752]$_DFFE_PN0P_  (.D(_01232_),
    .RN(net3662),
    .CLK(clknet_leaf_332_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[752] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[753]$_DFFE_PN0P_  (.D(_01233_),
    .RN(net3662),
    .CLK(clknet_6_7__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[753] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[754]$_DFFE_PN0P_  (.D(_01234_),
    .RN(net3664),
    .CLK(clknet_leaf_89_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[754] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[755]$_DFFE_PN0P_  (.D(_01235_),
    .RN(net3663),
    .CLK(clknet_leaf_284_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[755] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[756]$_DFFE_PN0P_  (.D(_01236_),
    .RN(net3664),
    .CLK(clknet_6_62__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[756] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[757]$_DFFE_PN0P_  (.D(_01237_),
    .RN(net3663),
    .CLK(clknet_leaf_196_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[757] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[758]$_DFFE_PN0P_  (.D(_01238_),
    .RN(net3662),
    .CLK(clknet_leaf_297_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[758] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[759]$_DFFE_PN0P_  (.D(_01239_),
    .RN(net3661),
    .CLK(clknet_leaf_399_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[759] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[75]$_DFFE_PN0P_  (.D(_01240_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[75] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[760]$_DFFE_PN0P_  (.D(_01241_),
    .RN(net3662),
    .CLK(clknet_leaf_380_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[760] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[761]$_DFFE_PN0P_  (.D(_01242_),
    .RN(net3663),
    .CLK(clknet_leaf_106_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[761] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[762]$_DFFE_PN0P_  (.D(_01243_),
    .RN(net3663),
    .CLK(clknet_leaf_185_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[762] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[763]$_DFFE_PN0P_  (.D(_01244_),
    .RN(net3663),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[763] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[764]$_DFFE_PN0P_  (.D(_01245_),
    .RN(net3663),
    .CLK(clknet_leaf_48_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[764] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[765]$_DFFE_PN0P_  (.D(_01246_),
    .RN(net3663),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[765] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[766]$_DFFE_PN0P_  (.D(_01247_),
    .RN(net3664),
    .CLK(clknet_leaf_65_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[766] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[767]$_DFFE_PN0P_  (.D(_01248_),
    .RN(net3662),
    .CLK(clknet_leaf_241_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[767] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[768]$_DFFE_PN0P_  (.D(_01249_),
    .RN(net3662),
    .CLK(clknet_leaf_319_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[768] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[769]$_DFFE_PN0P_  (.D(_01250_),
    .RN(net3661),
    .CLK(clknet_leaf_546_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[769] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[76]$_DFFE_PN0P_  (.D(_01251_),
    .RN(net3663),
    .CLK(clknet_leaf_167_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[76] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[770]$_DFFE_PN0P_  (.D(_01252_),
    .RN(net3662),
    .CLK(clknet_leaf_286_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[770] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[771]$_DFFE_PN0P_  (.D(_01253_),
    .RN(net3662),
    .CLK(clknet_leaf_302_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[771] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[772]$_DFFE_PN0P_  (.D(_01254_),
    .RN(net3662),
    .CLK(clknet_leaf_465_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[772] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[773]$_DFFE_PN0P_  (.D(_01255_),
    .RN(net3661),
    .CLK(clknet_6_27__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[773] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[774]$_DFFE_PN0P_  (.D(_01256_),
    .RN(net3661),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[774] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[775]$_DFFE_PN0P_  (.D(_01257_),
    .RN(net3661),
    .CLK(clknet_6_23__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[775] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[776]$_DFFE_PN0P_  (.D(_01258_),
    .RN(net3661),
    .CLK(clknet_leaf_549_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[776] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[777]$_DFFE_PN0P_  (.D(_01259_),
    .RN(net3661),
    .CLK(clknet_leaf_559_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[777] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[778]$_DFFE_PN0P_  (.D(_01260_),
    .RN(net3661),
    .CLK(clknet_6_20__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[778] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[779]$_DFFE_PN0P_  (.D(_01261_),
    .RN(net3663),
    .CLK(clknet_leaf_205_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[779] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[77]$_DFFE_PN0P_  (.D(_01262_),
    .RN(net3663),
    .CLK(clknet_leaf_134_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[77] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[780]$_DFFE_PN0P_  (.D(_01263_),
    .RN(net3663),
    .CLK(clknet_leaf_142_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[780] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[781]$_DFFE_PN0P_  (.D(_01264_),
    .RN(net3663),
    .CLK(clknet_leaf_129_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[781] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[782]$_DFFE_PN0P_  (.D(_01265_),
    .RN(net3661),
    .CLK(clknet_6_0__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[782] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[783]$_DFFE_PN0P_  (.D(_01266_),
    .RN(net3662),
    .CLK(clknet_6_2__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[783] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[784]$_DFFE_PN0P_  (.D(_01267_),
    .RN(net3662),
    .CLK(clknet_6_11__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[784] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[785]$_DFFE_PN0P_  (.D(_01268_),
    .RN(net3662),
    .CLK(clknet_6_6__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[785] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[786]$_DFFE_PN0P_  (.D(_01269_),
    .RN(net3663),
    .CLK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[786] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[787]$_DFFE_PN0P_  (.D(_01270_),
    .RN(net3662),
    .CLK(clknet_leaf_285_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[787] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[788]$_DFFE_PN0P_  (.D(_01271_),
    .RN(net3664),
    .CLK(clknet_6_62__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[788] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[789]$_DFFE_PN0P_  (.D(_01272_),
    .RN(net3663),
    .CLK(clknet_6_35__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[789] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[78]$_DFFE_PN0P_  (.D(_01273_),
    .RN(net3662),
    .CLK(clknet_leaf_426_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[78] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[790]$_DFFE_PN0P_  (.D(_01274_),
    .RN(net3662),
    .CLK(clknet_leaf_297_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[790] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[791]$_DFFE_PN0P_  (.D(_01275_),
    .RN(net3661),
    .CLK(clknet_6_1__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[791] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[792]$_DFFE_PN0P_  (.D(_01276_),
    .RN(net3662),
    .CLK(clknet_leaf_343_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[792] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[793]$_DFFE_PN0P_  (.D(_01277_),
    .RN(net3663),
    .CLK(clknet_leaf_111_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[793] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[794]$_DFFE_PN0P_  (.D(_01278_),
    .RN(net3663),
    .CLK(clknet_leaf_187_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[794] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[795]$_DFFE_PN0P_  (.D(_01279_),
    .RN(net3663),
    .CLK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[795] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[796]$_DFFE_PN0P_  (.D(_01280_),
    .RN(net3663),
    .CLK(clknet_leaf_58_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[796] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[797]$_DFFE_PN0P_  (.D(_01281_),
    .RN(net3663),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[797] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[798]$_DFFE_PN0P_  (.D(_01282_),
    .RN(net3663),
    .CLK(clknet_leaf_71_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[798] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[799]$_DFFE_PN0P_  (.D(_01283_),
    .RN(net3662),
    .CLK(clknet_6_32__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[799] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[79]$_DFFE_PN0P_  (.D(_01284_),
    .RN(net3662),
    .CLK(clknet_leaf_365_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[79] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[800]$_DFFE_PN0P_  (.D(_01285_),
    .RN(net3662),
    .CLK(clknet_leaf_319_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[800] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[801]$_DFFE_PN0P_  (.D(_01286_),
    .RN(net3661),
    .CLK(clknet_leaf_547_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[801] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[802]$_DFFE_PN0P_  (.D(_01287_),
    .RN(net3662),
    .CLK(clknet_leaf_277_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[802] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[803]$_DFFE_PN0P_  (.D(_01288_),
    .RN(net3662),
    .CLK(clknet_leaf_302_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[803] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[804]$_DFFE_PN0P_  (.D(_01289_),
    .RN(net3662),
    .CLK(clknet_6_5__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[804] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[805]$_DFFE_PN0P_  (.D(_01290_),
    .RN(net3661),
    .CLK(clknet_leaf_456_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[805] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[806]$_DFFE_PN0P_  (.D(_01291_),
    .RN(net3661),
    .CLK(clknet_6_29__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[806] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[807]$_DFFE_PN0P_  (.D(_01292_),
    .RN(net3661),
    .CLK(clknet_6_23__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[807] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[808]$_DFFE_PN0P_  (.D(_01293_),
    .RN(net3661),
    .CLK(clknet_6_17__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[808] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[809]$_DFFE_PN0P_  (.D(_01294_),
    .RN(net3661),
    .CLK(clknet_leaf_559_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[809] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[80]$_DFFE_PN0P_  (.D(_01295_),
    .RN(net3662),
    .CLK(clknet_leaf_320_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[80] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[810]$_DFFE_PN0P_  (.D(_01296_),
    .RN(net3661),
    .CLK(clknet_6_20__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[810] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[811]$_DFFE_PN0P_  (.D(_01297_),
    .RN(net3663),
    .CLK(clknet_6_36__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[811] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[812]$_DFFE_PN0P_  (.D(_01298_),
    .RN(net3663),
    .CLK(clknet_leaf_145_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[812] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[813]$_DFFE_PN0P_  (.D(_01299_),
    .RN(net3663),
    .CLK(clknet_6_59__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[813] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[814]$_DFFE_PN0P_  (.D(_01300_),
    .RN(net3661),
    .CLK(clknet_6_0__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[814] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[815]$_DFFE_PN0P_  (.D(_01301_),
    .RN(net3662),
    .CLK(clknet_leaf_385_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[815] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[816]$_DFFE_PN0P_  (.D(_01302_),
    .RN(net3662),
    .CLK(clknet_leaf_335_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[816] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[817]$_DFFE_PN0P_  (.D(_01303_),
    .RN(net3662),
    .CLK(clknet_leaf_433_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[817] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[818]$_DFFE_PN0P_  (.D(_01304_),
    .RN(net3663),
    .CLK(clknet_leaf_126_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[818] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[819]$_DFFE_PN0P_  (.D(_01305_),
    .RN(net3662),
    .CLK(clknet_leaf_285_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[819] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[81]$_DFFE_PN0P_  (.D(_01306_),
    .RN(net3662),
    .CLK(clknet_leaf_443_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[81] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[820]$_DFFE_PN0P_  (.D(_01307_),
    .RN(net3664),
    .CLK(clknet_6_63__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[820] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[821]$_DFFE_PN0P_  (.D(_01308_),
    .RN(net3663),
    .CLK(clknet_leaf_165_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[821] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[822]$_DFFE_PN0P_  (.D(_01309_),
    .RN(net3662),
    .CLK(clknet_leaf_299_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[822] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[823]$_DFFE_PN0P_  (.D(_01310_),
    .RN(net3661),
    .CLK(clknet_leaf_407_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[823] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[824]$_DFFE_PN0P_  (.D(_01311_),
    .RN(net3662),
    .CLK(clknet_6_8__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[824] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[825]$_DFFE_PN0P_  (.D(_01312_),
    .RN(net3663),
    .CLK(clknet_6_57__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[825] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[826]$_DFFE_PN0P_  (.D(_01313_),
    .RN(net3663),
    .CLK(clknet_leaf_186_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[826] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[827]$_DFFE_PN0P_  (.D(_01314_),
    .RN(net3663),
    .CLK(clknet_leaf_36_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[827] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[828]$_DFFE_PN0P_  (.D(_01315_),
    .RN(net3663),
    .CLK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[828] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[829]$_DFFE_PN0P_  (.D(_01316_),
    .RN(net3663),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[829] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[82]$_DFFE_PN0P_  (.D(_01317_),
    .RN(net3663),
    .CLK(clknet_leaf_119_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[82] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[830]$_DFFE_PN0P_  (.D(_01318_),
    .RN(net3663),
    .CLK(clknet_6_63__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[830] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[831]$_DFFE_PN0P_  (.D(_01319_),
    .RN(net3662),
    .CLK(clknet_leaf_260_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[831] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[832]$_DFFE_PN0P_  (.D(_01320_),
    .RN(net3662),
    .CLK(clknet_6_9__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[832] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[833]$_DFFE_PN0P_  (.D(_01321_),
    .RN(net3661),
    .CLK(clknet_leaf_547_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[833] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[834]$_DFFE_PN0P_  (.D(_01322_),
    .RN(net3662),
    .CLK(clknet_leaf_276_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[834] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[835]$_DFFE_PN0P_  (.D(_01323_),
    .RN(net3662),
    .CLK(clknet_leaf_303_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[835] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[836]$_DFFE_PN0P_  (.D(_01324_),
    .RN(net3662),
    .CLK(clknet_leaf_467_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[836] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[837]$_DFFE_PN0P_  (.D(_01325_),
    .RN(net3661),
    .CLK(clknet_leaf_486_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[837] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[838]$_DFFE_PN0P_  (.D(_01326_),
    .RN(net3661),
    .CLK(clknet_6_23__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[838] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[839]$_DFFE_PN0P_  (.D(_01327_),
    .RN(net3661),
    .CLK(clknet_leaf_566_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[839] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[83]$_DFFE_PN0P_  (.D(_01328_),
    .RN(net3663),
    .CLK(clknet_leaf_147_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[83] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[840]$_DFFE_PN0P_  (.D(_01329_),
    .RN(net3661),
    .CLK(clknet_leaf_551_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[840] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[841]$_DFFE_PN0P_  (.D(_01330_),
    .RN(net3661),
    .CLK(clknet_leaf_560_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[841] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[842]$_DFFE_PN0P_  (.D(_01331_),
    .RN(net3661),
    .CLK(clknet_leaf_501_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[842] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[843]$_DFFE_PN0P_  (.D(_01332_),
    .RN(net3663),
    .CLK(clknet_leaf_207_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[843] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[844]$_DFFE_PN0P_  (.D(_01333_),
    .RN(net3663),
    .CLK(clknet_leaf_149_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[844] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[845]$_DFFE_PN0P_  (.D(_01334_),
    .RN(net3663),
    .CLK(clknet_6_58__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[845] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[846]$_DFFE_PN0P_  (.D(_01335_),
    .RN(net3661),
    .CLK(clknet_leaf_393_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[846] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[847]$_DFFE_PN0P_  (.D(_01336_),
    .RN(net3662),
    .CLK(clknet_leaf_386_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[847] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[848]$_DFFE_PN0P_  (.D(_01337_),
    .RN(net3662),
    .CLK(clknet_leaf_338_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[848] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[849]$_DFFE_PN0P_  (.D(_01338_),
    .RN(net3662),
    .CLK(clknet_leaf_433_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[849] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[84]$_DFFE_PN0P_  (.D(_01339_),
    .RN(net3664),
    .CLK(clknet_6_62__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[84] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[850]$_DFFE_PN0P_  (.D(_01340_),
    .RN(net3663),
    .CLK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[850] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[851]$_DFFE_PN0P_  (.D(_01341_),
    .RN(net3662),
    .CLK(clknet_leaf_281_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[851] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[852]$_DFFE_PN0P_  (.D(_01342_),
    .RN(net3664),
    .CLK(clknet_6_63__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[852] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[853]$_DFFE_PN0P_  (.D(_01343_),
    .RN(net3663),
    .CLK(clknet_leaf_193_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[853] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[854]$_DFFE_PN0P_  (.D(_01344_),
    .RN(net3662),
    .CLK(clknet_6_14__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[854] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[855]$_DFFE_PN0P_  (.D(_01345_),
    .RN(net3661),
    .CLK(clknet_leaf_402_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[855] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[856]$_DFFE_PN0P_  (.D(_01346_),
    .RN(net3662),
    .CLK(clknet_leaf_379_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[856] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[857]$_DFFE_PN0P_  (.D(_01347_),
    .RN(net3663),
    .CLK(clknet_6_56__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[857] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[858]$_DFFE_PN0P_  (.D(_01348_),
    .RN(net3663),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[858] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[859]$_DFFE_PN0P_  (.D(_01349_),
    .RN(net3663),
    .CLK(clknet_6_52__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[859] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[85]$_DFFE_PN0P_  (.D(_01350_),
    .RN(net3662),
    .CLK(clknet_leaf_266_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[85] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[860]$_DFFE_PN0P_  (.D(_01351_),
    .RN(net3663),
    .CLK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[860] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[861]$_DFFE_PN0P_  (.D(_01352_),
    .RN(net3663),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[861] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[862]$_DFFE_PN0P_  (.D(_01353_),
    .RN(net3663),
    .CLK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[862] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[863]$_DFFE_PN0P_  (.D(_01354_),
    .RN(net3662),
    .CLK(clknet_leaf_235_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[863] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[864]$_DFFE_PN0P_  (.D(_01355_),
    .RN(net3662),
    .CLK(clknet_6_12__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[864] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[865]$_DFFE_PN0P_  (.D(_01356_),
    .RN(net3661),
    .CLK(clknet_leaf_546_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[865] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[866]$_DFFE_PN0P_  (.D(_01357_),
    .RN(net3662),
    .CLK(clknet_leaf_276_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[866] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[867]$_DFFE_PN0P_  (.D(_01358_),
    .RN(net3662),
    .CLK(clknet_leaf_303_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[867] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[868]$_DFFE_PN0P_  (.D(_01359_),
    .RN(net3662),
    .CLK(clknet_leaf_466_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[868] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[869]$_DFFE_PN0P_  (.D(_01360_),
    .RN(net3661),
    .CLK(clknet_leaf_456_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[869] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[86]$_DFFE_PN0P_  (.D(_01361_),
    .RN(net3662),
    .CLK(clknet_leaf_317_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[86] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[870]$_DFFE_PN0P_  (.D(_01362_),
    .RN(net3661),
    .CLK(clknet_6_23__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[870] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[871]$_DFFE_PN0P_  (.D(_01363_),
    .RN(net3661),
    .CLK(clknet_leaf_566_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[871] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[872]$_DFFE_PN0P_  (.D(_01364_),
    .RN(net3661),
    .CLK(clknet_leaf_549_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[872] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[873]$_DFFE_PN0P_  (.D(_01365_),
    .RN(net3661),
    .CLK(clknet_leaf_561_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[873] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[874]$_DFFE_PN0P_  (.D(_01366_),
    .RN(net3661),
    .CLK(clknet_leaf_501_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[874] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[875]$_DFFE_PN0P_  (.D(_01367_),
    .RN(net3663),
    .CLK(clknet_leaf_207_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[875] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[876]$_DFFE_PN0P_  (.D(_01368_),
    .RN(net3663),
    .CLK(clknet_6_46__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[876] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[877]$_DFFE_PN0P_  (.D(_01369_),
    .RN(net3663),
    .CLK(clknet_6_58__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[877] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[878]$_DFFE_PN0P_  (.D(_01370_),
    .RN(net3661),
    .CLK(clknet_leaf_393_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[878] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[879]$_DFFE_PN0P_  (.D(_01371_),
    .RN(net3662),
    .CLK(clknet_leaf_386_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[879] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[87]$_DFFE_PN0P_  (.D(_01372_),
    .RN(net3661),
    .CLK(clknet_leaf_424_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[87] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[880]$_DFFE_PN0P_  (.D(_01373_),
    .RN(net3662),
    .CLK(clknet_leaf_338_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[880] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[881]$_DFFE_PN0P_  (.D(_01374_),
    .RN(net3662),
    .CLK(clknet_6_6__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[881] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[882]$_DFFE_PN0P_  (.D(_01375_),
    .RN(net3663),
    .CLK(clknet_leaf_122_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[882] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[883]$_DFFE_PN0P_  (.D(_01376_),
    .RN(net3662),
    .CLK(clknet_leaf_281_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[883] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[884]$_DFFE_PN0P_  (.D(_01377_),
    .RN(net3664),
    .CLK(clknet_leaf_77_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[884] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[885]$_DFFE_PN0P_  (.D(_01378_),
    .RN(net3663),
    .CLK(clknet_leaf_193_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[885] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[886]$_DFFE_PN0P_  (.D(_01379_),
    .RN(net3662),
    .CLK(clknet_leaf_299_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[886] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[887]$_DFFE_PN0P_  (.D(_01380_),
    .RN(net3661),
    .CLK(clknet_leaf_402_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[887] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[888]$_DFFE_PN0P_  (.D(_01381_),
    .RN(net3662),
    .CLK(clknet_leaf_379_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[888] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[889]$_DFFE_PN0P_  (.D(_01382_),
    .RN(net3663),
    .CLK(clknet_leaf_177_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[889] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[88]$_DFFE_PN0P_  (.D(_01383_),
    .RN(net3662),
    .CLK(clknet_leaf_365_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[88] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[890]$_DFFE_PN0P_  (.D(_01384_),
    .RN(net3663),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[890] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[891]$_DFFE_PN0P_  (.D(_01385_),
    .RN(net3663),
    .CLK(clknet_6_52__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[891] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[892]$_DFFE_PN0P_  (.D(_01386_),
    .RN(net3663),
    .CLK(clknet_leaf_57_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[892] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[893]$_DFFE_PN0P_  (.D(_01387_),
    .RN(net3663),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[893] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[894]$_DFFE_PN0P_  (.D(_01388_),
    .RN(net3663),
    .CLK(clknet_leaf_68_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[894] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[895]$_DFFE_PN0P_  (.D(_01389_),
    .RN(net3662),
    .CLK(clknet_leaf_235_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[895] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[896]$_DFFE_PN0P_  (.D(_01390_),
    .RN(net3662),
    .CLK(clknet_6_9__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[896] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[897]$_DFFE_PN0P_  (.D(_01391_),
    .RN(net3661),
    .CLK(clknet_leaf_550_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[897] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[898]$_DFFE_PN0P_  (.D(_01392_),
    .RN(net3662),
    .CLK(clknet_6_42__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[898] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[899]$_DFFE_PN0P_  (.D(_01393_),
    .RN(net3662),
    .CLK(clknet_leaf_306_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[899] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[89]$_DFFE_PN0P_  (.D(_01394_),
    .RN(net3663),
    .CLK(clknet_leaf_169_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[89] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[900]$_DFFE_PN0P_  (.D(_01395_),
    .RN(net3662),
    .CLK(clknet_leaf_465_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[900] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[901]$_DFFE_PN0P_  (.D(_01396_),
    .RN(net3661),
    .CLK(clknet_leaf_462_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[901] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[902]$_DFFE_PN0P_  (.D(_01397_),
    .RN(net3661),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[902] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[903]$_DFFE_PN0P_  (.D(_01398_),
    .RN(net3661),
    .CLK(clknet_leaf_566_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[903] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[904]$_DFFE_PN0P_  (.D(_01399_),
    .RN(net3661),
    .CLK(clknet_leaf_551_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[904] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[905]$_DFFE_PN0P_  (.D(_01400_),
    .RN(net3661),
    .CLK(clknet_6_20__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[905] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[906]$_DFFE_PN0P_  (.D(_01401_),
    .RN(net3661),
    .CLK(clknet_6_20__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[906] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[907]$_DFFE_PN0P_  (.D(_01402_),
    .RN(net3663),
    .CLK(clknet_leaf_208_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[907] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[908]$_DFFE_PN0P_  (.D(_01403_),
    .RN(net3663),
    .CLK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[908] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[909]$_DFFE_PN0P_  (.D(_01404_),
    .RN(net3663),
    .CLK(clknet_leaf_139_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[909] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[90]$_DFFE_PN0P_  (.D(_01405_),
    .RN(net3663),
    .CLK(clknet_leaf_201_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[90] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[910]$_DFFE_PN0P_  (.D(_01406_),
    .RN(net3661),
    .CLK(clknet_leaf_391_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[910] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[911]$_DFFE_PN0P_  (.D(_01407_),
    .RN(net3662),
    .CLK(clknet_leaf_389_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[911] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[912]$_DFFE_PN0P_  (.D(_01408_),
    .RN(net3662),
    .CLK(clknet_leaf_332_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[912] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[913]$_DFFE_PN0P_  (.D(_01409_),
    .RN(net3662),
    .CLK(clknet_leaf_442_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[913] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[914]$_DFFE_PN0P_  (.D(_01410_),
    .RN(net3663),
    .CLK(clknet_6_59__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[914] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[915]$_DFFE_PN0P_  (.D(_01411_),
    .RN(net3662),
    .CLK(clknet_leaf_145_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[915] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[916]$_DFFE_PN0P_  (.D(_01412_),
    .RN(net3664),
    .CLK(clknet_6_63__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[916] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[917]$_DFFE_PN0P_  (.D(_01413_),
    .RN(net3663),
    .CLK(clknet_6_35__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[917] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[918]$_DFFE_PN0P_  (.D(_01414_),
    .RN(net3662),
    .CLK(clknet_6_14__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[918] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[919]$_DFFE_PN0P_  (.D(_01415_),
    .RN(net3661),
    .CLK(clknet_leaf_405_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[919] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[91]$_DFFE_PN0P_  (.D(_01416_),
    .RN(net3663),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[91] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[920]$_DFFE_PN0P_  (.D(_01417_),
    .RN(net3662),
    .CLK(clknet_6_10__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[920] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[921]$_DFFE_PN0P_  (.D(_01418_),
    .RN(net3663),
    .CLK(clknet_6_50__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[921] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[922]$_DFFE_PN0P_  (.D(_01419_),
    .RN(net3663),
    .CLK(clknet_leaf_185_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[922] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[923]$_DFFE_PN0P_  (.D(_01420_),
    .RN(net3663),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[923] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[924]$_DFFE_PN0P_  (.D(_01421_),
    .RN(net3663),
    .CLK(clknet_leaf_53_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[924] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[925]$_DFFE_PN0P_  (.D(_01422_),
    .RN(net3663),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[925] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[926]$_DFFE_PN0P_  (.D(_01423_),
    .RN(net3663),
    .CLK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[926] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[927]$_DFFE_PN0P_  (.D(_01424_),
    .RN(net3662),
    .CLK(clknet_leaf_252_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[927] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[928]$_DFFE_PN0P_  (.D(_01425_),
    .RN(net3662),
    .CLK(clknet_leaf_312_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[928] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[929]$_DFFE_PN0P_  (.D(_01426_),
    .RN(net3661),
    .CLK(clknet_leaf_548_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[929] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[92]$_DFFE_PN0P_  (.D(_01427_),
    .RN(net3663),
    .CLK(clknet_leaf_108_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[92] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[930]$_DFFE_PN0P_  (.D(_01428_),
    .RN(net3662),
    .CLK(clknet_leaf_289_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[930] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[931]$_DFFE_PN0P_  (.D(_01429_),
    .RN(net3662),
    .CLK(clknet_leaf_306_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[931] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[932]$_DFFE_PN0P_  (.D(_01430_),
    .RN(net3662),
    .CLK(clknet_leaf_466_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[932] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[933]$_DFFE_PN0P_  (.D(_01431_),
    .RN(net3661),
    .CLK(clknet_6_30__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[933] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[934]$_DFFE_PN0P_  (.D(_01432_),
    .RN(net3661),
    .CLK(clknet_leaf_571_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[934] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[935]$_DFFE_PN0P_  (.D(_01433_),
    .RN(net3661),
    .CLK(clknet_leaf_566_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[935] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[936]$_DFFE_PN0P_  (.D(_01434_),
    .RN(net3661),
    .CLK(clknet_leaf_551_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[936] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[937]$_DFFE_PN0P_  (.D(_01435_),
    .RN(net3661),
    .CLK(clknet_leaf_561_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[937] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[938]$_DFFE_PN0P_  (.D(_01436_),
    .RN(net3661),
    .CLK(clknet_leaf_563_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[938] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[939]$_DFFE_PN0P_  (.D(_01437_),
    .RN(net3663),
    .CLK(clknet_leaf_208_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[939] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[93]$_DFFE_PN0P_  (.D(_01438_),
    .RN(net3663),
    .CLK(clknet_leaf_39_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[93] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[940]$_DFFE_PN0P_  (.D(_01439_),
    .RN(net3663),
    .CLK(clknet_leaf_137_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[940] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[941]$_DFFE_PN0P_  (.D(_01440_),
    .RN(net3663),
    .CLK(clknet_6_58__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[941] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[942]$_DFFE_PN0P_  (.D(_01441_),
    .RN(net3661),
    .CLK(clknet_leaf_391_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[942] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[943]$_DFFE_PN0P_  (.D(_01442_),
    .RN(net3662),
    .CLK(clknet_6_2__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[943] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[944]$_DFFE_PN0P_  (.D(_01443_),
    .RN(net3662),
    .CLK(clknet_6_11__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[944] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[945]$_DFFE_PN0P_  (.D(_01444_),
    .RN(net3662),
    .CLK(clknet_leaf_247_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[945] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[946]$_DFFE_PN0P_  (.D(_01445_),
    .RN(net3663),
    .CLK(clknet_6_59__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[946] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[947]$_DFFE_PN0P_  (.D(_01446_),
    .RN(net3662),
    .CLK(clknet_leaf_277_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[947] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[948]$_DFFE_PN0P_  (.D(_01447_),
    .RN(net3664),
    .CLK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[948] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[949]$_DFFE_PN0P_  (.D(_01448_),
    .RN(net3663),
    .CLK(clknet_6_35__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[949] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[94]$_DFFE_PN0P_  (.D(_01449_),
    .RN(net3663),
    .CLK(clknet_leaf_100_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[94] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[950]$_DFFE_PN0P_  (.D(_01450_),
    .RN(net3662),
    .CLK(clknet_6_14__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[950] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[951]$_DFFE_PN0P_  (.D(_01451_),
    .RN(net3661),
    .CLK(clknet_leaf_403_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[951] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[952]$_DFFE_PN0P_  (.D(_01452_),
    .RN(net3662),
    .CLK(clknet_leaf_349_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[952] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[953]$_DFFE_PN0P_  (.D(_01453_),
    .RN(net3663),
    .CLK(clknet_leaf_182_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[953] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[954]$_DFFE_PN0P_  (.D(_01454_),
    .RN(net3663),
    .CLK(clknet_6_49__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[954] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[955]$_DFFE_PN0P_  (.D(_01455_),
    .RN(net3663),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[955] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[956]$_DFFE_PN0P_  (.D(_01456_),
    .RN(net3663),
    .CLK(clknet_leaf_54_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[956] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[957]$_DFFE_PN0P_  (.D(_01457_),
    .RN(net3663),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[957] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[958]$_DFFE_PN0P_  (.D(_01458_),
    .RN(net3663),
    .CLK(clknet_leaf_67_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[958] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[959]$_DFFE_PN0P_  (.D(_01459_),
    .RN(net3662),
    .CLK(clknet_leaf_260_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[959] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[95]$_DFFE_PN0P_  (.D(_01460_),
    .RN(net3662),
    .CLK(clknet_leaf_237_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[95] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[960]$_DFFE_PN0P_  (.D(_01461_),
    .RN(net3662),
    .CLK(clknet_leaf_361_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[960] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[961]$_DFFE_PN0P_  (.D(_01462_),
    .RN(net3661),
    .CLK(clknet_leaf_548_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[961] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[962]$_DFFE_PN0P_  (.D(_01463_),
    .RN(net3662),
    .CLK(clknet_leaf_289_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[962] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[963]$_DFFE_PN0P_  (.D(_01464_),
    .RN(net3662),
    .CLK(clknet_leaf_304_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[963] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[964]$_DFFE_PN0P_  (.D(_01465_),
    .RN(net3662),
    .CLK(clknet_leaf_467_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[964] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[965]$_DFFE_PN0P_  (.D(_01466_),
    .RN(net3661),
    .CLK(clknet_6_30__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[965] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[966]$_DFFE_PN0P_  (.D(_01467_),
    .RN(net3661),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[966] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[967]$_DFFE_PN0P_  (.D(_01468_),
    .RN(net3661),
    .CLK(clknet_leaf_565_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[967] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[968]$_DFFE_PN0P_  (.D(_01469_),
    .RN(net3661),
    .CLK(clknet_leaf_551_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[968] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[969]$_DFFE_PN0P_  (.D(_01470_),
    .RN(net3661),
    .CLK(clknet_leaf_560_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[969] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[96]$_DFFE_PN0P_  (.D(_01471_),
    .RN(net3662),
    .CLK(clknet_leaf_248_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[96] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[970]$_DFFE_PN0P_  (.D(_01472_),
    .RN(net3661),
    .CLK(clknet_leaf_563_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[970] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[971]$_DFFE_PN0P_  (.D(_01473_),
    .RN(net3663),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[971] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[972]$_DFFE_PN0P_  (.D(_01474_),
    .RN(net3663),
    .CLK(clknet_leaf_149_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[972] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[973]$_DFFE_PN0P_  (.D(_01475_),
    .RN(net3663),
    .CLK(clknet_6_58__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[973] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[974]$_DFFE_PN0P_  (.D(_01476_),
    .RN(net3661),
    .CLK(clknet_leaf_407_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[974] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[975]$_DFFE_PN0P_  (.D(_01477_),
    .RN(net3662),
    .CLK(clknet_leaf_389_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[975] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[976]$_DFFE_PN0P_  (.D(_01478_),
    .RN(net3662),
    .CLK(clknet_leaf_322_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[976] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[977]$_DFFE_PN0P_  (.D(_01479_),
    .RN(net3662),
    .CLK(clknet_leaf_442_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[977] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[978]$_DFFE_PN0P_  (.D(_01480_),
    .RN(net3663),
    .CLK(clknet_6_59__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[978] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[979]$_DFFE_PN0P_  (.D(_01481_),
    .RN(net3662),
    .CLK(clknet_leaf_280_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[979] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[97]$_DFFE_PN0P_  (.D(_01482_),
    .RN(net3661),
    .CLK(clknet_6_18__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[97] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[980]$_DFFE_PN0P_  (.D(_01483_),
    .RN(net3664),
    .CLK(clknet_leaf_75_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[980] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[981]$_DFFE_PN0P_  (.D(_01484_),
    .RN(net3663),
    .CLK(clknet_leaf_197_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[981] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[982]$_DFFE_PN0P_  (.D(_01485_),
    .RN(net3662),
    .CLK(clknet_leaf_324_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[982] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[983]$_DFFE_PN0P_  (.D(_01486_),
    .RN(net3661),
    .CLK(clknet_6_24__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[983] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[984]$_DFFE_PN0P_  (.D(_01487_),
    .RN(net3662),
    .CLK(clknet_6_8__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[984] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[985]$_DFFE_PN0P_  (.D(_01488_),
    .RN(net3663),
    .CLK(clknet_leaf_182_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[985] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[986]$_DFFE_PN0P_  (.D(_01489_),
    .RN(net3663),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[986] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[987]$_DFFE_PN0P_  (.D(_01490_),
    .RN(net3663),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[987] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[988]$_DFFE_PN0P_  (.D(_01491_),
    .RN(net3663),
    .CLK(clknet_leaf_56_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[988] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[989]$_DFFE_PN0P_  (.D(_01492_),
    .RN(net3663),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[989] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[98]$_DFFE_PN0P_  (.D(_01493_),
    .RN(net3662),
    .CLK(clknet_leaf_255_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[98] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[990]$_DFFE_PN0P_  (.D(_01494_),
    .RN(net3663),
    .CLK(clknet_leaf_60_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[990] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[991]$_DFFE_PN0P_  (.D(_01495_),
    .RN(net3662),
    .CLK(clknet_leaf_258_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[991] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[992]$_DFFE_PN0P_  (.D(_01496_),
    .RN(net3662),
    .CLK(clknet_leaf_361_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[992] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[993]$_DFFE_PN0P_  (.D(_01497_),
    .RN(net3661),
    .CLK(clknet_leaf_550_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[993] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[994]$_DFFE_PN0P_  (.D(_01498_),
    .RN(net3662),
    .CLK(clknet_leaf_289_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[994] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[995]$_DFFE_PN0P_  (.D(_01499_),
    .RN(net3662),
    .CLK(clknet_leaf_304_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[995] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[996]$_DFFE_PN0P_  (.D(_01500_),
    .RN(net3662),
    .CLK(clknet_6_5__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[996] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[997]$_DFFE_PN0P_  (.D(_01501_),
    .RN(net3661),
    .CLK(clknet_6_30__leaf_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[997] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[998]$_DFFE_PN0P_  (.D(_01502_),
    .RN(net3661),
    .CLK(clknet_leaf_571_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[998] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[999]$_DFFE_PN0P_  (.D(_01503_),
    .RN(net3661),
    .CLK(clknet_leaf_565_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[999] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[99]$_DFFE_PN0P_  (.D(_01504_),
    .RN(net3662),
    .CLK(clknet_leaf_254_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[99] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.branch_set$_DFF_PN0_  (.D(\id_stage_i.branch_set_d ),
    .RN(net3661),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\id_stage_i.branch_set ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.D(_01505_),
    .RN(net148),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.D(_01506_),
    .RN(net3661),
    .CLK(clknet_leaf_27_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.D(_01507_),
    .RN(net148),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.D(_01508_),
    .RN(net3661),
    .CLK(clknet_leaf_27_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.debug_mode_o$_DFFE_PN0P_  (.D(_01509_),
    .RN(net3661),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\cs_registers_i.debug_mode_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.exc_req_d ),
    .RN(net3661),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\id_stage_i.controller_i.exc_req_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.illegal_insn_d ),
    .RN(net3661),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\id_stage_i.controller_i.illegal_insn_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.load_err_i ),
    .RN(net3661),
    .CLK(clknet_leaf_522_clk),
    .Q(\id_stage_i.controller_i.load_err_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.nmi_mode_o$_DFFE_PN0P_  (.D(_01510_),
    .RN(net148),
    .CLK(clknet_leaf_25_clk),
    .Q(\cs_registers_i.nmi_mode_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.store_err_i ),
    .RN(net3661),
    .CLK(clknet_leaf_522_clk),
    .Q(\id_stage_i.controller_i.store_err_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.D(_01511_),
    .RN(net3661),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\id_stage_i.id_fsm_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[0]$_DFFE_PN0P_  (.D(_01512_),
    .RN(net148),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[10]$_DFFE_PN0P_  (.D(_01513_),
    .RN(net148),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[11]$_DFFE_PN0P_  (.D(_01514_),
    .RN(net148),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[12]$_DFFE_PN0P_  (.D(_01515_),
    .RN(net148),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[13]$_DFFE_PN0P_  (.D(_01516_),
    .RN(net148),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[14]$_DFFE_PN0P_  (.D(_01517_),
    .RN(net148),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[15]$_DFFE_PN0P_  (.D(_01518_),
    .RN(net148),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[16]$_DFFE_PN0P_  (.D(_01519_),
    .RN(net148),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[17]$_DFFE_PN0P_  (.D(_01520_),
    .RN(net148),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[18]$_DFFE_PN0P_  (.D(_01521_),
    .RN(net148),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[19]$_DFFE_PN0P_  (.D(_01522_),
    .RN(net148),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[1]$_DFFE_PN0P_  (.D(_01523_),
    .RN(net148),
    .CLK(clknet_leaf_468_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[20]$_DFFE_PN0P_  (.D(_01524_),
    .RN(net3660),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[21]$_DFFE_PN0P_  (.D(_01525_),
    .RN(net3660),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[22]$_DFFE_PN0P_  (.D(_01526_),
    .RN(net148),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[23]$_DFFE_PN0P_  (.D(_01527_),
    .RN(net148),
    .CLK(clknet_leaf_452_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[24]$_DFFE_PN0P_  (.D(_01528_),
    .RN(net148),
    .CLK(clknet_6_55__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[25]$_DFFE_PN0P_  (.D(_01529_),
    .RN(net148),
    .CLK(clknet_leaf_455_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[26]$_DFFE_PN0P_  (.D(_01530_),
    .RN(net148),
    .CLK(clknet_leaf_452_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[27]$_DFFE_PN0P_  (.D(_01531_),
    .RN(net148),
    .CLK(clknet_leaf_459_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[28]$_DFFE_PN0P_  (.D(_01532_),
    .RN(net148),
    .CLK(clknet_leaf_459_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[29]$_DFFE_PN0P_  (.D(_01533_),
    .RN(net148),
    .CLK(clknet_leaf_455_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[2]$_DFFE_PN0P_  (.D(_01534_),
    .RN(net148),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[30]$_DFFE_PN0P_  (.D(_01535_),
    .RN(net148),
    .CLK(clknet_6_53__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[31]$_DFFE_PN0P_  (.D(_01536_),
    .RN(net3660),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[34]$_DFFE_PN0P_  (.D(_01537_),
    .RN(net3660),
    .CLK(clknet_leaf_398_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[35]$_DFFE_PN0P_  (.D(_01538_),
    .RN(net3660),
    .CLK(clknet_leaf_398_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[36]$_DFFE_PN0P_  (.D(_01539_),
    .RN(net3660),
    .CLK(clknet_leaf_440_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[37]$_DFFE_PN0P_  (.D(_01540_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[38]$_DFFE_PN0P_  (.D(_01541_),
    .RN(net3660),
    .CLK(clknet_6_54__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[39]$_DFFE_PN0P_  (.D(_01542_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[3]$_DFFE_PN0P_  (.D(_01543_),
    .RN(net148),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[40]$_DFFE_PN0P_  (.D(_01544_),
    .RN(net3660),
    .CLK(clknet_leaf_401_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[41]$_DFFE_PN0P_  (.D(_01545_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[42]$_DFFE_PN0P_  (.D(_01546_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[43]$_DFFE_PN0P_  (.D(_01547_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[44]$_DFFE_PN0P_  (.D(_01548_),
    .RN(net3660),
    .CLK(clknet_6_60__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[45]$_DFFE_PN0P_  (.D(_01549_),
    .RN(net3660),
    .CLK(clknet_leaf_440_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[46]$_DFFE_PN0P_  (.D(_01550_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[47]$_DFFE_PN0P_  (.D(_01551_),
    .RN(net3660),
    .CLK(clknet_leaf_401_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[48]$_DFFE_PN0P_  (.D(_01552_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[49]$_DFFE_PN0P_  (.D(_01553_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[4]$_DFFE_PN0P_  (.D(_01554_),
    .RN(net148),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[50]$_DFFE_PN0P_  (.D(_01555_),
    .RN(net3660),
    .CLK(clknet_leaf_437_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[51]$_DFFE_PN0P_  (.D(_01556_),
    .RN(net3660),
    .CLK(clknet_leaf_437_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[52]$_DFFE_PN0P_  (.D(_01557_),
    .RN(net3660),
    .CLK(clknet_leaf_436_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[53]$_DFFE_PN0P_  (.D(_01558_),
    .RN(net3660),
    .CLK(clknet_leaf_436_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[54]$_DFFE_PN0P_  (.D(_01559_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[55]$_DFFE_PN0P_  (.D(_01560_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[56]$_DFFE_PN0P_  (.D(_01561_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[57]$_DFFE_PN0P_  (.D(_01562_),
    .RN(net3660),
    .CLK(clknet_leaf_428_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[58]$_DFFE_PN0P_  (.D(_01563_),
    .RN(net3660),
    .CLK(clknet_leaf_428_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[59]$_DFFE_PN0P_  (.D(_01564_),
    .RN(net3660),
    .CLK(clknet_leaf_427_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[5]$_DFFE_PN0P_  (.D(_01565_),
    .RN(net148),
    .CLK(clknet_leaf_468_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[60]$_DFFE_PN0P_  (.D(_01566_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[61]$_DFFE_PN0P_  (.D(_01567_),
    .RN(net3660),
    .CLK(clknet_6_61__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[62]$_DFFE_PN0P_  (.D(_01568_),
    .RN(net3660),
    .CLK(clknet_leaf_427_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[63]$_DFFE_PN0P_  (.D(_01569_),
    .RN(net3660),
    .CLK(clknet_leaf_426_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[64]$_DFFE_PN0P_  (.D(_01570_),
    .RN(net3660),
    .CLK(clknet_leaf_426_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[65]$_DFFE_PN0P_  (.D(_01571_),
    .RN(net3660),
    .CLK(clknet_6_63__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[66]$_DFFE_PN0P_  (.D(_01572_),
    .RN(net3660),
    .CLK(clknet_leaf_425_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[67]$_DFFE_PN0P_  (.D(_01573_),
    .RN(net3660),
    .CLK(clknet_leaf_425_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[6]$_DFFE_PN0P_  (.D(_01574_),
    .RN(net148),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[7]$_DFFE_PN0P_  (.D(_01575_),
    .RN(net148),
    .CLK(clknet_6_52__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[8]$_DFFE_PN0P_  (.D(_01576_),
    .RN(net148),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[9]$_DFFE_PN0P_  (.D(_01577_),
    .RN(net148),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .RN(net148),
    .CLK(clknet_leaf_608_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .RN(net148),
    .CLK(clknet_leaf_608_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .RN(net148),
    .CLK(clknet_leaf_609_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.D(_01578_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.D(_01579_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.D(_01580_),
    .CLK(clknet_leaf_228_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.D(_01581_),
    .CLK(clknet_leaf_226_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.D(_01582_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.D(_01583_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.D(_01584_),
    .CLK(clknet_leaf_238_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.D(_01585_),
    .CLK(clknet_leaf_242_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.D(_01586_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.D(_01587_),
    .CLK(clknet_leaf_240_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.D(_01588_),
    .CLK(clknet_leaf_375_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.D(_01589_),
    .CLK(clknet_leaf_376_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.D(_01590_),
    .CLK(clknet_6_57__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.D(_01591_),
    .CLK(clknet_leaf_375_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.D(_01592_),
    .CLK(clknet_6_58__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.D(_01593_),
    .CLK(clknet_6_58__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.D(_01594_),
    .CLK(clknet_leaf_360_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.D(_01595_),
    .CLK(clknet_leaf_361_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.D(_01596_),
    .CLK(clknet_leaf_360_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.D(_01597_),
    .CLK(clknet_leaf_361_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.D(_01598_),
    .CLK(clknet_leaf_242_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.D(_01599_),
    .CLK(clknet_leaf_364_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.D(_01600_),
    .CLK(clknet_leaf_364_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.D(_01601_),
    .CLK(clknet_leaf_354_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.D(_01602_),
    .CLK(clknet_6_59__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.D(_01603_),
    .CLK(clknet_leaf_352_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.D(_01604_),
    .CLK(clknet_leaf_372_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.D(_01605_),
    .CLK(clknet_leaf_375_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.D(_01606_),
    .CLK(clknet_6_58__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.D(_01607_),
    .CLK(clknet_leaf_228_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.D(_01608_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.D(_01609_),
    .CLK(clknet_leaf_530_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.D(_01610_),
    .CLK(clknet_leaf_530_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.D(_01611_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.D(_01612_),
    .CLK(clknet_leaf_248_clk),
    .Q(\cs_registers_i.pc_if_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.D(_01613_),
    .CLK(clknet_leaf_250_clk),
    .Q(\cs_registers_i.pc_if_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.D(_01614_),
    .CLK(clknet_leaf_248_clk),
    .Q(\cs_registers_i.pc_if_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.D(_01615_),
    .CLK(clknet_6_45__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.D(_01616_),
    .CLK(clknet_leaf_250_clk),
    .Q(\cs_registers_i.pc_if_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.D(_01617_),
    .CLK(clknet_leaf_252_clk),
    .Q(\cs_registers_i.pc_if_i[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.D(_01618_),
    .CLK(clknet_leaf_253_clk),
    .Q(\cs_registers_i.pc_if_i[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.D(_01619_),
    .CLK(clknet_leaf_244_clk),
    .Q(\cs_registers_i.pc_if_i[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.D(_01620_),
    .CLK(clknet_leaf_253_clk),
    .Q(\cs_registers_i.pc_if_i[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.D(_01621_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.D(_01622_),
    .CLK(clknet_6_18__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.D(_01623_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.D(_01624_),
    .CLK(clknet_leaf_351_clk),
    .Q(\cs_registers_i.pc_if_i[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.D(_01625_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.D(_01626_),
    .CLK(clknet_leaf_358_clk),
    .Q(\cs_registers_i.pc_if_i[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.D(_01627_),
    .CLK(clknet_leaf_243_clk),
    .Q(\cs_registers_i.pc_if_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.D(_01628_),
    .CLK(clknet_leaf_354_clk),
    .Q(\cs_registers_i.pc_if_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.D(_01629_),
    .CLK(clknet_leaf_358_clk),
    .Q(\cs_registers_i.pc_if_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.D(_01630_),
    .CLK(clknet_leaf_353_clk),
    .Q(\cs_registers_i.pc_if_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.D(_01631_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.D(_01632_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.D(_01633_),
    .CLK(clknet_leaf_255_clk),
    .Q(\cs_registers_i.pc_if_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.D(_01634_),
    .CLK(clknet_leaf_345_clk),
    .Q(\cs_registers_i.pc_if_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.D(_01635_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.D(_01636_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_if_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.D(_01637_),
    .CLK(clknet_leaf_344_clk),
    .Q(\cs_registers_i.pc_if_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.D(_01638_),
    .CLK(clknet_leaf_255_clk),
    .Q(\cs_registers_i.pc_if_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.D(_01639_),
    .CLK(clknet_leaf_344_clk),
    .Q(\cs_registers_i.pc_if_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.D(_01640_),
    .CLK(clknet_leaf_247_clk),
    .Q(\cs_registers_i.pc_if_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.D(_01641_),
    .CLK(clknet_leaf_247_clk),
    .Q(\cs_registers_i.pc_if_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.D(_01642_),
    .CLK(clknet_leaf_531_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.D(_01643_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.D(_01644_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.D(_01645_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.D(_01646_),
    .CLK(clknet_leaf_559_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.D(_01647_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.D(_01648_),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.D(_01649_),
    .CLK(clknet_leaf_601_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.D(_01650_),
    .CLK(clknet_leaf_601_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.D(_01651_),
    .CLK(clknet_leaf_587_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.D(_01652_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.D(_01653_),
    .CLK(clknet_leaf_531_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.D(_01654_),
    .CLK(clknet_6_1__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.D(_01655_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.D(_01656_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.D(_01657_),
    .CLK(clknet_leaf_571_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.D(_01658_),
    .CLK(clknet_leaf_587_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.D(_01659_),
    .CLK(clknet_6_0__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.D(_01660_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.D(_01661_),
    .CLK(clknet_leaf_572_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.D(_01662_),
    .CLK(clknet_leaf_573_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.D(_01663_),
    .CLK(clknet_leaf_571_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.D(_01664_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.D(_01665_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.D(_01666_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.D(_01667_),
    .CLK(clknet_leaf_533_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.D(_01668_),
    .CLK(clknet_leaf_532_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.D(_01669_),
    .CLK(clknet_leaf_546_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.D(_01670_),
    .CLK(clknet_leaf_580_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.D(_01671_),
    .CLK(clknet_leaf_549_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.D(_01672_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.D(_01673_),
    .CLK(clknet_leaf_553_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.D(_01674_),
    .CLK(clknet_leaf_555_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.D(_01675_),
    .CLK(clknet_leaf_580_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.D(_01676_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.D(_01677_),
    .CLK(clknet_leaf_569_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.D(_01678_),
    .CLK(clknet_leaf_567_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.D(_01679_),
    .CLK(clknet_leaf_552_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.D(_01680_),
    .CLK(clknet_leaf_575_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.D(_01681_),
    .CLK(clknet_leaf_559_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.D(_01682_),
    .CLK(clknet_leaf_560_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.D(_01683_),
    .CLK(clknet_leaf_564_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.D(_01684_),
    .CLK(clknet_leaf_593_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.D(_01685_),
    .CLK(clknet_leaf_592_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.D(_01686_),
    .CLK(clknet_leaf_550_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.D(_01687_),
    .CLK(clknet_leaf_590_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.D(_01688_),
    .CLK(clknet_leaf_584_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.D(_01689_),
    .CLK(clknet_leaf_590_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.D(_01690_),
    .CLK(clknet_leaf_583_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.D(_01691_),
    .CLK(clknet_leaf_583_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.D(_01692_),
    .CLK(clknet_leaf_588_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.D(_01693_),
    .CLK(clknet_leaf_589_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.D(_01694_),
    .CLK(clknet_leaf_594_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.D(_01695_),
    .CLK(clknet_leaf_570_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.D(_01696_),
    .CLK(clknet_leaf_572_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.D(_01697_),
    .CLK(clknet_leaf_550_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.D(_01698_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.D(_01699_),
    .CLK(clknet_6_0__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.D(_01700_),
    .CLK(clknet_leaf_593_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.D(_01701_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.D(_01702_),
    .CLK(clknet_leaf_533_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.D(_01703_),
    .CLK(clknet_leaf_532_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.D(_01704_),
    .CLK(clknet_leaf_546_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.D(_01705_),
    .CLK(clknet_leaf_580_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.D(_01706_),
    .CLK(clknet_leaf_549_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.D(_01707_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.D(_01708_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.D(_01709_),
    .CLK(clknet_leaf_553_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.D(_01710_),
    .CLK(clknet_leaf_555_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.D(_01711_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.D(_01712_),
    .CLK(clknet_leaf_569_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.D(_01713_),
    .CLK(clknet_leaf_567_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.D(_01714_),
    .CLK(clknet_leaf_552_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.D(_01715_),
    .CLK(clknet_leaf_575_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.D(_01716_),
    .CLK(clknet_leaf_559_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.D(_01717_),
    .CLK(clknet_leaf_560_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.D(_01718_),
    .CLK(clknet_leaf_564_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.D(_01719_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.D(_01720_),
    .CLK(clknet_leaf_592_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.D(_01721_),
    .CLK(clknet_leaf_592_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.D(_01722_),
    .CLK(clknet_leaf_589_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.D(_01723_),
    .CLK(clknet_leaf_584_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.D(_01724_),
    .CLK(clknet_leaf_590_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.D(_01725_),
    .CLK(clknet_6_4__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.D(_01726_),
    .CLK(clknet_leaf_580_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.D(_01727_),
    .CLK(clknet_leaf_588_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.D(_01728_),
    .CLK(clknet_leaf_588_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.D(_01729_),
    .CLK(clknet_leaf_594_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.D(_01730_),
    .CLK(clknet_6_5__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.D(_01731_),
    .CLK(clknet_leaf_570_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.D(_01732_),
    .CLK(clknet_leaf_572_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.D(_01733_),
    .CLK(clknet_leaf_573_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.D(_01734_),
    .CLK(clknet_6_0__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.D(_01735_),
    .CLK(clknet_leaf_594_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.D(_01736_),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.D(_01737_),
    .CLK(clknet_6_6__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .RN(net148),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .RN(net148),
    .CLK(clknet_6_7__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .RN(net148),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .RN(net148),
    .CLK(clknet_6_2__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .RN(net148),
    .CLK(clknet_6_3__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.D(_01738_),
    .CLK(clknet_leaf_224_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.D(_01739_),
    .CLK(clknet_leaf_224_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.D(_01740_),
    .CLK(clknet_leaf_226_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.D(_01741_),
    .CLK(clknet_leaf_225_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.D(_01742_),
    .CLK(clknet_leaf_238_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.D(_01743_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.D(_01744_),
    .CLK(clknet_leaf_238_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.D(_01745_),
    .CLK(clknet_leaf_240_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.D(_01746_),
    .CLK(clknet_6_47__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.D(_01747_),
    .CLK(clknet_leaf_240_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.D(_01748_),
    .CLK(clknet_6_59__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.D(_01749_),
    .CLK(clknet_6_59__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.D(_01750_),
    .CLK(clknet_leaf_376_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.D(_01751_),
    .CLK(clknet_leaf_376_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.D(_01752_),
    .CLK(clknet_leaf_241_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.D(_01753_),
    .CLK(clknet_leaf_241_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.D(_01754_),
    .CLK(clknet_leaf_366_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.D(_01755_),
    .CLK(clknet_leaf_365_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.D(_01756_),
    .CLK(clknet_leaf_363_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.D(_01757_),
    .CLK(clknet_leaf_363_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.D(_01758_),
    .CLK(clknet_leaf_242_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.D(_01759_),
    .CLK(clknet_leaf_365_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.D(_01760_),
    .CLK(clknet_leaf_366_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.D(_01761_),
    .CLK(clknet_leaf_372_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.D(_01762_),
    .CLK(clknet_6_59__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.D(_01763_),
    .CLK(clknet_leaf_384_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.D(_01764_),
    .CLK(clknet_6_59__leaf_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.D(_01765_),
    .CLK(clknet_leaf_377_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.D(_01766_),
    .CLK(clknet_leaf_377_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.D(_01767_),
    .CLK(clknet_leaf_225_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .RN(net148),
    .CLK(clknet_leaf_609_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.illegal_c_insn_id_o$_DFFE_PN_  (.D(_01768_),
    .CLK(clknet_leaf_497_clk),
    .Q(\id_stage_i.decoder_i.illegal_c_insn_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_fetch_err_o$_DFFE_PN_  (.D(_01769_),
    .CLK(clknet_leaf_528_clk),
    .Q(\id_stage_i.controller_i.instr_fetch_err_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0N_  (.D(_01770_),
    .CLK(clknet_6_16__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_fetch_err_plus2_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_is_compressed_id_o$_DFFE_PN_  (.D(_01771_),
    .CLK(clknet_leaf_534_clk),
    .Q(\id_stage_i.controller_i.instr_is_compressed_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PN_  (.D(_01772_),
    .CLK(clknet_leaf_540_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PN_  (.D(_01773_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PN_  (.D(_01774_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PN_  (.D(_01775_),
    .CLK(clknet_leaf_543_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PN_  (.D(_01776_),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PN_  (.D(_01777_),
    .CLK(clknet_leaf_503_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PN_  (.D(_01778_),
    .CLK(clknet_leaf_503_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PN_  (.D(_01779_),
    .CLK(clknet_leaf_534_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PN_  (.D(_01780_),
    .CLK(clknet_leaf_514_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PN_  (.D(_01781_),
    .CLK(clknet_leaf_514_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PN_  (.D(_01782_),
    .CLK(clknet_leaf_543_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PN_  (.D(_01783_),
    .CLK(clknet_leaf_539_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PN_  (.D(_01784_),
    .CLK(clknet_leaf_537_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PN_  (.D(_01785_),
    .CLK(clknet_leaf_544_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PN_  (.D(_01786_),
    .CLK(clknet_leaf_544_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PN_  (.D(_01787_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[0]$_DFFE_PN_  (.D(_01788_),
    .CLK(clknet_leaf_540_clk),
    .Q(\id_stage_i.controller_i.instr_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[10]$_DFFE_PN_  (.D(_01789_),
    .CLK(clknet_leaf_537_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[11]$_DFFE_PN_  (.D(_01790_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[12]$_DFFE_PN_  (.D(_01791_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[13]$_DFFE_PN_  (.D(_01792_),
    .CLK(clknet_leaf_497_clk),
    .Q(\id_stage_i.controller_i.instr_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[14]$_DFFE_PN_  (.D(_01793_),
    .CLK(clknet_leaf_499_clk),
    .Q(\id_stage_i.controller_i.instr_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[15]$_DFFE_PN_  (.D(_01794_),
    .CLK(clknet_leaf_502_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[16]$_DFFE_PN_  (.D(_01795_),
    .CLK(clknet_leaf_501_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[17]$_DFFE_PN_  (.D(_01796_),
    .CLK(clknet_leaf_501_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[18]$_DFFE_PN_  (.D(_01797_),
    .CLK(clknet_6_20__leaf_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[19]$_DFFE_PN_  (.D(_01798_),
    .CLK(clknet_6_20__leaf_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[1]$_DFFE_PN_  (.D(_01799_),
    .CLK(clknet_leaf_534_clk),
    .Q(\id_stage_i.controller_i.instr_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[20]$_DFFE_PN_  (.D(_01800_),
    .CLK(clknet_6_21__leaf_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[21]$_DFFE_PN_  (.D(_01801_),
    .CLK(clknet_leaf_497_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[22]$_DFFE_PN_  (.D(_01802_),
    .CLK(clknet_leaf_498_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[23]$_DFFE_PN_  (.D(_01803_),
    .CLK(clknet_leaf_499_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[24]$_DFFE_PN_  (.D(_01804_),
    .CLK(clknet_leaf_499_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[25]$_DFFE_PN_  (.D(_01805_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[26]$_DFFE_PN_  (.D(_01806_),
    .CLK(clknet_leaf_515_clk),
    .Q(\id_stage_i.controller_i.instr_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[27]$_DFFE_PN_  (.D(_01807_),
    .CLK(clknet_leaf_520_clk),
    .Q(\id_stage_i.controller_i.instr_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[28]$_DFFE_PN_  (.D(_01808_),
    .CLK(clknet_leaf_521_clk),
    .Q(\id_stage_i.controller_i.instr_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[29]$_DFFE_PN_  (.D(_01809_),
    .CLK(clknet_leaf_521_clk),
    .Q(\id_stage_i.controller_i.instr_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[2]$_DFFE_PN_  (.D(_01810_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[30]$_DFFE_PN_  (.D(_01811_),
    .CLK(clknet_6_19__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[31]$_DFFE_PN_  (.D(_01812_),
    .CLK(clknet_leaf_520_clk),
    .Q(\id_stage_i.controller_i.instr_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[3]$_DFFE_PN_  (.D(_01813_),
    .CLK(clknet_leaf_515_clk),
    .Q(\id_stage_i.controller_i.instr_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[4]$_DFFE_PN_  (.D(_01814_),
    .CLK(clknet_6_22__leaf_clk),
    .Q(\id_stage_i.controller_i.instr_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[5]$_DFFE_PN_  (.D(_01815_),
    .CLK(clknet_leaf_543_clk),
    .Q(\id_stage_i.controller_i.instr_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[6]$_DFFE_PN_  (.D(_01816_),
    .CLK(clknet_leaf_539_clk),
    .Q(\id_stage_i.controller_i.instr_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[7]$_DFFE_PN_  (.D(_01817_),
    .CLK(clknet_leaf_502_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[8]$_DFFE_PN_  (.D(_01818_),
    .CLK(clknet_leaf_498_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[9]$_DFFE_PN_  (.D(_01819_),
    .CLK(clknet_6_17__leaf_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.instr_valid_id_o$_DFF_PN0_  (.D(\if_stage_i.instr_valid_id_d ),
    .RN(net3661),
    .CLK(clknet_leaf_528_clk),
    .Q(\id_stage_i.controller_i.instr_valid_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[10]$_DFFE_PN_  (.D(_01820_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[11]$_DFFE_PN_  (.D(_01821_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[12]$_DFFE_PN_  (.D(_01822_),
    .CLK(clknet_leaf_297_clk),
    .Q(\cs_registers_i.pc_id_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[13]$_DFFE_PN_  (.D(_01823_),
    .CLK(clknet_leaf_297_clk),
    .Q(\cs_registers_i.pc_id_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[14]$_DFFE_PN_  (.D(_01824_),
    .CLK(clknet_leaf_252_clk),
    .Q(\cs_registers_i.pc_id_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[15]$_DFFE_PN_  (.D(_01825_),
    .CLK(clknet_leaf_293_clk),
    .Q(\cs_registers_i.pc_id_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[16]$_DFFE_PN_  (.D(_01826_),
    .CLK(clknet_leaf_252_clk),
    .Q(\cs_registers_i.pc_id_i[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[17]$_DFFE_PN_  (.D(_01827_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[18]$_DFFE_PN_  (.D(_01828_),
    .CLK(clknet_leaf_244_clk),
    .Q(\cs_registers_i.pc_id_i[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[19]$_DFFE_PN_  (.D(_01829_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[1]$_DFFE_PN_  (.D(_01830_),
    .CLK(clknet_leaf_32_clk),
    .Q(\cs_registers_i.pc_id_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[20]$_DFFE_PN_  (.D(_01831_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[21]$_DFFE_PN_  (.D(_01832_),
    .CLK(clknet_leaf_345_clk),
    .Q(\cs_registers_i.pc_id_i[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[22]$_DFFE_PN_  (.D(_01833_),
    .CLK(clknet_leaf_351_clk),
    .Q(\cs_registers_i.pc_id_i[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[23]$_DFFE_PN_  (.D(_01834_),
    .CLK(clknet_leaf_243_clk),
    .Q(\cs_registers_i.pc_id_i[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[24]$_DFFE_PN_  (.D(_01835_),
    .CLK(clknet_leaf_358_clk),
    .Q(\cs_registers_i.pc_id_i[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[25]$_DFFE_PN_  (.D(_01836_),
    .CLK(clknet_6_58__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[26]$_DFFE_PN_  (.D(_01837_),
    .CLK(clknet_leaf_353_clk),
    .Q(\cs_registers_i.pc_id_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[27]$_DFFE_PN_  (.D(_01838_),
    .CLK(clknet_6_58__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[28]$_DFFE_PN_  (.D(_01839_),
    .CLK(clknet_leaf_352_clk),
    .Q(\cs_registers_i.pc_id_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[29]$_DFFE_PN_  (.D(_01840_),
    .CLK(clknet_6_56__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[2]$_DFFE_PN_  (.D(_01841_),
    .CLK(clknet_leaf_33_clk),
    .Q(\cs_registers_i.pc_id_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[30]$_DFFE_PN_  (.D(_01842_),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[31]$_DFFE_PN_  (.D(_01843_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[3]$_DFFE_PN_  (.D(_01844_),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[4]$_DFFE_PN_  (.D(_01845_),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[5]$_DFFE_PN_  (.D(_01846_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[6]$_DFFE_PN_  (.D(_01847_),
    .CLK(clknet_6_37__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[7]$_DFFE_PN_  (.D(_01848_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[8]$_DFFE_PN_  (.D(_01849_),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[9]$_DFFE_PN_  (.D(_01850_),
    .CLK(clknet_6_39__leaf_clk),
    .Q(\cs_registers_i.pc_id_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[0]$_DFFE_PN0P_  (.D(_01851_),
    .RN(net3661),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[10]$_DFFE_PN0P_  (.D(_01852_),
    .RN(net148),
    .CLK(clknet_leaf_312_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[11]$_DFFE_PN0P_  (.D(_01853_),
    .RN(net148),
    .CLK(clknet_leaf_312_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[12]$_DFFE_PN0P_  (.D(_01854_),
    .RN(net148),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[13]$_DFFE_PN0P_  (.D(_01855_),
    .RN(net148),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[14]$_DFFE_PN0P_  (.D(_01856_),
    .RN(net148),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[15]$_DFFE_PN0P_  (.D(_01857_),
    .RN(net148),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[16]$_DFFE_PN0P_  (.D(_01858_),
    .RN(net148),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[17]$_DFFE_PN0P_  (.D(_01859_),
    .RN(net148),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[18]$_DFFE_PN0P_  (.D(_01860_),
    .RN(net148),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[19]$_DFFE_PN0P_  (.D(_01861_),
    .RN(net3660),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[1]$_DFFE_PN0P_  (.D(_01862_),
    .RN(net3661),
    .CLK(clknet_6_25__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[20]$_DFFE_PN0P_  (.D(_01863_),
    .RN(net3660),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[21]$_DFFE_PN0P_  (.D(_01864_),
    .RN(net3660),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[22]$_DFFE_PN0P_  (.D(_01865_),
    .RN(net3660),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[23]$_DFFE_PN0P_  (.D(_01866_),
    .RN(net3660),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[24]$_DFFE_PN0P_  (.D(_01867_),
    .RN(net3660),
    .CLK(clknet_leaf_344_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[25]$_DFFE_PN0P_  (.D(_01868_),
    .RN(net3660),
    .CLK(clknet_6_50__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[26]$_DFFE_PN0P_  (.D(_01869_),
    .RN(net3660),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[27]$_DFFE_PN0P_  (.D(_01870_),
    .RN(net3660),
    .CLK(clknet_leaf_323_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[28]$_DFFE_PN0P_  (.D(_01871_),
    .RN(net3660),
    .CLK(clknet_6_51__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[29]$_DFFE_PN0P_  (.D(_01872_),
    .RN(net3660),
    .CLK(clknet_leaf_323_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[2]$_DFFE_PN0P_  (.D(_01873_),
    .RN(net148),
    .CLK(clknet_leaf_511_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[30]$_DFFE_PN0P_  (.D(_01874_),
    .RN(net3660),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[31]$_DFFE_PN0P_  (.D(_01875_),
    .RN(net148),
    .CLK(clknet_6_48__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[3]$_DFFE_PN0P_  (.D(_01876_),
    .RN(net148),
    .CLK(clknet_leaf_511_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[4]$_DFFE_PN0P_  (.D(_01877_),
    .RN(net148),
    .CLK(clknet_6_27__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[5]$_DFFE_PN0P_  (.D(_01878_),
    .RN(net148),
    .CLK(clknet_leaf_307_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[6]$_DFFE_PN0P_  (.D(_01879_),
    .RN(net148),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[7]$_DFFE_PN0P_  (.D(_01880_),
    .RN(net148),
    .CLK(clknet_leaf_307_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[8]$_DFFE_PN0P_  (.D(_01881_),
    .RN(net148),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[9]$_DFFE_PN0P_  (.D(_01882_),
    .RN(net148),
    .CLK(clknet_6_49__leaf_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.D(_01883_),
    .RN(net3663),
    .CLK(clknet_leaf_475_clk),
    .Q(\load_store_unit_i.data_sign_ext_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.D(_01884_),
    .RN(net3661),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\load_store_unit_i.data_we_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.D(_01885_),
    .RN(net3661),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\load_store_unit_i.handle_misaligned_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.D(_01886_),
    .RN(net3661),
    .CLK(clknet_leaf_504_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.D(_01887_),
    .RN(net3661),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.D(_01888_),
    .RN(net3661),
    .CLK(clknet_leaf_504_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.D(_01889_),
    .RN(net3661),
    .CLK(clknet_6_23__leaf_clk),
    .Q(\load_store_unit_i.lsu_err_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.D(_01890_),
    .RN(net3663),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\load_store_unit_i.rdata_offset_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.D(_01891_),
    .RN(net3663),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\load_store_unit_i.rdata_offset_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[0]$_DFFE_PN0P_  (.D(_01892_),
    .RN(net3663),
    .CLK(clknet_leaf_495_clk),
    .Q(\load_store_unit_i.rdata_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.D(_01893_),
    .RN(net3663),
    .CLK(clknet_leaf_479_clk),
    .Q(\load_store_unit_i.rdata_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.D(_01894_),
    .RN(net3663),
    .CLK(clknet_leaf_489_clk),
    .Q(\load_store_unit_i.rdata_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.D(_01895_),
    .RN(net3663),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.D(_01896_),
    .RN(net3663),
    .CLK(clknet_leaf_486_clk),
    .Q(\load_store_unit_i.rdata_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.D(_01897_),
    .RN(net3663),
    .CLK(clknet_leaf_485_clk),
    .Q(\load_store_unit_i.rdata_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.D(_01898_),
    .RN(net3663),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.D(_01899_),
    .RN(net3663),
    .CLK(clknet_leaf_476_clk),
    .Q(\load_store_unit_i.rdata_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.D(_01900_),
    .RN(net3663),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.D(_01901_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.D(_01902_),
    .RN(net3663),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[1]$_DFFE_PN0P_  (.D(_01903_),
    .RN(net3663),
    .CLK(clknet_leaf_494_clk),
    .Q(\load_store_unit_i.rdata_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.D(_01904_),
    .RN(net3663),
    .CLK(clknet_6_29__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.D(_01905_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.D(_01906_),
    .RN(net3663),
    .CLK(clknet_6_31__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.D(_01907_),
    .RN(net3663),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[2]$_DFFE_PN0P_  (.D(_01908_),
    .RN(net3663),
    .CLK(clknet_leaf_479_clk),
    .Q(\load_store_unit_i.rdata_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[3]$_DFFE_PN0P_  (.D(_01909_),
    .RN(net3663),
    .CLK(clknet_leaf_489_clk),
    .Q(\load_store_unit_i.rdata_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[4]$_DFFE_PN0P_  (.D(_01910_),
    .RN(net3663),
    .CLK(clknet_6_28__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[5]$_DFFE_PN0P_  (.D(_01911_),
    .RN(net3663),
    .CLK(clknet_leaf_486_clk),
    .Q(\load_store_unit_i.rdata_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[6]$_DFFE_PN0P_  (.D(_01912_),
    .RN(net3663),
    .CLK(clknet_leaf_485_clk),
    .Q(\load_store_unit_i.rdata_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[7]$_DFFE_PN0P_  (.D(_01913_),
    .RN(net3663),
    .CLK(clknet_6_30__leaf_clk),
    .Q(\load_store_unit_i.rdata_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.D(_01914_),
    .RN(net3663),
    .CLK(clknet_leaf_495_clk),
    .Q(\load_store_unit_i.rdata_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.D(_01915_),
    .RN(net3663),
    .CLK(clknet_leaf_494_clk),
    .Q(\load_store_unit_i.rdata_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Right_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Right_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Right_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Right_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Right_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Right_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Right_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Right_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Right_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Right_205 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Right_206 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Right_207 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Right_208 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Right_209 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Right_210 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Right_211 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Right_212 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Right_213 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Right_214 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Right_215 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Right_216 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Right_217 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Right_218 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Right_219 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Right_220 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Right_221 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Right_222 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Right_223 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Right_224 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Right_225 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Right_226 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Right_227 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Right_228 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Right_229 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Right_230 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Right_231 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Right_232 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Right_233 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Right_234 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_235 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_236 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_237 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_238 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_239 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_240 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_241 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_242 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_243 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_244 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_245 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_246 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_247 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_248 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_249 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_250 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_251 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_252 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_253 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_254 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_255 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_256 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_257 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_258 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_259 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_260 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_261 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_262 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_263 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_264 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_265 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_266 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_267 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_268 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_269 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_270 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_271 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_272 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_273 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_274 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_275 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_276 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_277 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_278 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_279 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_280 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_281 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_282 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_283 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_284 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_285 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_286 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_287 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_288 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_289 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_290 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_291 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_292 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_293 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_294 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_295 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_296 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_297 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_298 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_299 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_300 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_301 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_302 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_303 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_304 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_305 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_306 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_307 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_308 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_309 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_310 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_311 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_312 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_313 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_314 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_315 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_316 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_317 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_318 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_319 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_320 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_321 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_322 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_323 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_324 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_325 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_326 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_327 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_328 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_329 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_330 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_331 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_332 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_333 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_334 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_335 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_336 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_337 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_338 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_339 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_340 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_341 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_342 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_343 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_344 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_345 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_346 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_347 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_348 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_349 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_350 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_351 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_352 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_353 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_354 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_355 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_356 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_357 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_358 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_359 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_360 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_361 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_362 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_363 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_364 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_365 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_366 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_367 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_368 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_369 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_370 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_371 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_372 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_373 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_374 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_375 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_376 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_377 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_378 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_379 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_380 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_381 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_382 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_383 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_384 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_385 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_386 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_387 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_388 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_389 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_390 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_391 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_392 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_393 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_394 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_395 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_396 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_397 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_398 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_399 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_400 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_401 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_402 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_403 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_404 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_405 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_406 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_407 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_408 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_409 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_410 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_411 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_412 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_413 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_414 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_415 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_416 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_417 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_418 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_419 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_420 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_421 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_422 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_423 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_424 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_425 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_426 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_427 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_428 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_429 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Left_430 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Left_431 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Left_432 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Left_433 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Left_434 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Left_435 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Left_436 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Left_437 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Left_438 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Left_439 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Left_440 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Left_441 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Left_442 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Left_443 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Left_444 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Left_445 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Left_446 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Left_447 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Left_448 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Left_449 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Left_450 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Left_451 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Left_452 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Left_453 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Left_454 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Left_455 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Left_456 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Left_457 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Left_458 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Left_459 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Left_460 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Left_461 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Left_462 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Left_463 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Left_464 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Left_465 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Left_466 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Left_467 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Left_468 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Left_469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_772 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_773 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_774 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_775 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_776 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_777 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_778 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_779 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_780 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_781 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_782 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_783 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_784 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_785 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_786 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_787 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_788 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_789 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_790 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_791 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_792 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_793 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_794 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_795 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_796 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_797 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_798 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_799 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_800 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_801 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_802 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_803 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_804 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_805 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_806 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_807 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_808 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_809 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_810 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_811 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_812 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_813 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_814 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_815 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_816 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_817 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_818 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_819 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_820 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_821 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_822 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_823 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_824 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_825 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_826 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_827 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_828 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_829 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_830 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_831 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_832 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_833 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_834 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_835 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_836 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_837 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_838 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_839 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_840 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_841 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_842 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_843 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_844 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_845 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_846 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_847 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_848 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_849 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_850 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_851 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_852 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_853 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_854 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_855 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_856 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_857 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_858 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_859 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_860 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_861 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_862 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_863 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_864 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_865 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_866 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_867 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_868 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_869 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_870 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_871 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_872 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_873 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_874 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_875 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_876 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_877 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_878 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_879 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_880 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_881 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_882 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_883 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_884 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_885 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_886 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_887 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_888 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_889 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_890 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_891 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_892 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_893 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_894 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_895 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_896 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_897 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_898 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_899 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_900 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_901 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_902 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_903 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_904 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_905 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_906 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_907 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_908 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_909 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_910 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_911 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_912 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_913 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_914 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_915 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_916 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_917 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_918 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_919 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_920 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_921 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_922 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_923 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_924 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_925 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_926 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_927 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_928 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_929 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_930 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_931 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_932 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_933 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_934 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_935 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_936 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_937 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_938 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_939 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_940 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_941 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_942 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_943 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_944 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_945 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_946 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_947 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_948 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_949 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_950 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_951 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_952 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_953 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_954 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_955 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_956 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_957 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_958 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_959 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_960 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_961 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_962 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_963 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_964 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_965 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_966 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_967 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_968 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_969 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_970 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_971 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_972 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_973 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_974 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_975 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_976 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_977 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_978 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_979 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_980 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_981 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_982 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_983 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_984 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_985 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_986 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_987 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_988 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_989 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_990 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_991 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_992 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_993 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_994 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_995 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_996 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_997 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_998 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_999 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3472 (.I(\load_store_unit_i.ls_fsm_cs[2] ),
    .Z(net3472));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3474 (.I(net355),
    .Z(net3474));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3476 (.I(\id_stage_i.controller_i.instr_i[4] ),
    .Z(net3476));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3488 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .Z(net3488));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3479 (.I(\id_stage_i.controller_i.instr_i[31] ),
    .Z(net3479));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3481 (.I(\id_stage_i.controller_i.instr_i[2] ),
    .Z(net3481));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3482 (.I(\id_stage_i.controller_i.instr_i[29] ),
    .Z(net3482));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3483 (.I(\id_stage_i.controller_i.instr_i[28] ),
    .Z(net3483));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3484 (.I(\id_stage_i.controller_i.instr_i[27] ),
    .Z(net3484));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3485 (.I(\id_stage_i.controller_i.instr_i[26] ),
    .Z(net3485));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3486 (.I(\id_stage_i.controller_i.instr_i[25] ),
    .Z(net3486));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3487 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .Z(net3487));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3490 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(net3490));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3506 (.I(net3505),
    .Z(net3506));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3529 (.I(net3513),
    .Z(net3529));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3560 (.I(net3559),
    .Z(net3560));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3556 (.I(net3553),
    .Z(net3556));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3600 (.I(net3597),
    .Z(net3600));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3603 (.I(net3597),
    .Z(net3603));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3598 (.I(net3597),
    .Z(net3598));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3597 (.I(net3589),
    .Z(net3597));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3607 (.I(net333),
    .Z(net3607));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22913__2 (.ZN(net251));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3611 (.I(net333),
    .Z(net3611));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3606 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .Z(net3606));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3610 (.I(net3609),
    .Z(net3610));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3441 (.I(_06367_),
    .Z(net3441));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3649 (.I(\id_stage_i.controller_i.instr_i[12] ),
    .Z(net3649));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3440 (.I(_06367_),
    .Z(net3440));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3571 (.I(net3569),
    .Z(net3571));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_89_clk_i_regs (.I(clknet_6_62__leaf_clk_i_regs),
    .Z(clknet_leaf_89_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_87_clk_i_regs (.I(clknet_6_62__leaf_clk_i_regs),
    .Z(clknet_leaf_87_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_84_clk_i_regs (.I(clknet_6_62__leaf_clk_i_regs),
    .Z(clknet_leaf_84_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_80_clk_i_regs (.I(clknet_6_62__leaf_clk_i_regs),
    .Z(clknet_leaf_80_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_79_clk_i_regs (.I(clknet_6_62__leaf_clk_i_regs),
    .Z(clknet_leaf_79_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_clk_i_regs (.I(clknet_6_37__leaf_clk_i_regs),
    .Z(clknet_leaf_9_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_60_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_60_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3568 (.I(net3567),
    .Z(net3568));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3609 (.I(net416),
    .Z(net3609));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3583 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .Z(net3583));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3635 (.I(net3634),
    .Z(net3635));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3585 (.I(net3583),
    .Z(net3585));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3582 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .Z(net3582));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3242 (.I(net3240),
    .Z(net3242));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3581 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .Z(net3581));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3439 (.I(_06367_),
    .Z(net3439));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_36_clk_i_regs (.I(clknet_6_52__leaf_clk_i_regs),
    .Z(clknet_leaf_36_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3229 (.I(net3228),
    .Z(net3229));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3438 (.I(net3437),
    .Z(net3438));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_35_clk_i_regs (.I(clknet_6_52__leaf_clk_i_regs),
    .Z(clknet_leaf_35_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22946__5 (.ZN(net254));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3437 (.I(_06367_),
    .Z(net3437));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_34_clk_i_regs (.I(clknet_6_53__leaf_clk_i_regs),
    .Z(clknet_leaf_34_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk_i_regs (.I(clknet_6_48__leaf_clk_i_regs),
    .Z(clknet_leaf_12_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3124 (.I(net3123),
    .Z(net3124));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3122 (.I(_11279_[0]),
    .Z(net3122));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3436 (.I(_06367_),
    .Z(net3436));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3133 (.I(_11348_[0]),
    .Z(net3133));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_31_clk_i_regs (.I(clknet_6_52__leaf_clk_i_regs),
    .Z(clknet_leaf_31_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_29_clk_i_regs (.I(clknet_6_53__leaf_clk_i_regs),
    .Z(clknet_leaf_29_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3132 (.I(_11349_[0]),
    .Z(net3132));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3435 (.I(net3434),
    .Z(net3435));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk_i_regs (.I(clknet_6_48__leaf_clk_i_regs),
    .Z(clknet_leaf_11_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3217 (.I(net3216),
    .Z(net3217));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3538 (.I(net3534),
    .Z(net3538));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_26_clk_i_regs (.I(clknet_6_53__leaf_clk_i_regs),
    .Z(clknet_leaf_26_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3434 (.I(_06367_),
    .Z(net3434));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3622 (.I(net449),
    .Z(net3622));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3130 (.I(_03309_),
    .Z(net3130));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3140 (.I(_11330_[0]),
    .Z(net3140));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_28_clk_i_regs (.I(clknet_6_53__leaf_clk_i_regs),
    .Z(clknet_leaf_28_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3620 (.I(net3619),
    .Z(net3620));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_24_clk_i_regs (.I(clknet_6_53__leaf_clk_i_regs),
    .Z(clknet_leaf_24_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk_i_regs (.I(clknet_6_52__leaf_clk_i_regs),
    .Z(clknet_leaf_18_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3621 (.I(net3619),
    .Z(net3621));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_clk_i_regs (.I(clknet_6_52__leaf_clk_i_regs),
    .Z(clknet_leaf_17_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_23_clk_i_regs (.I(clknet_6_53__leaf_clk_i_regs),
    .Z(clknet_leaf_23_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk_i_regs (.I(clknet_6_52__leaf_clk_i_regs),
    .Z(clknet_leaf_22_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_27_clk_i_regs (.I(clknet_6_53__leaf_clk_i_regs),
    .Z(clknet_leaf_27_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3135 (.I(net3134),
    .Z(net3135));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3282 (.I(net3281),
    .Z(net3282));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3144 (.I(net3143),
    .Z(net3144));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3269 (.I(net3268),
    .Z(net3269));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3260 (.I(net3259),
    .Z(net3260));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk_i_regs (.I(clknet_6_49__leaf_clk_i_regs),
    .Z(clknet_leaf_21_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_clk_i_regs (.I(clknet_6_37__leaf_clk_i_regs),
    .Z(clknet_leaf_10_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk_i_regs (.I(clknet_6_49__leaf_clk_i_regs),
    .Z(clknet_leaf_20_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3246 (.I(net3245),
    .Z(net3246));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3245 (.I(net3244),
    .Z(net3245));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_77_clk_i_regs (.I(clknet_6_63__leaf_clk_i_regs),
    .Z(clknet_leaf_77_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_75_clk_i_regs (.I(clknet_6_63__leaf_clk_i_regs),
    .Z(clknet_leaf_75_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_74_clk_i_regs (.I(clknet_6_63__leaf_clk_i_regs),
    .Z(clknet_leaf_74_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3634 (.I(net3606),
    .Z(net3634));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3633 (.I(net417),
    .Z(net3633));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_71_clk_i_regs (.I(clknet_6_63__leaf_clk_i_regs),
    .Z(clknet_leaf_71_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_68_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_68_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 place3632 (.I(net3631),
    .Z(net3632));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3552 (.I(net433),
    .Z(net3552));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3551 (.I(net3550),
    .Z(net3551));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3550 (.I(net423),
    .Z(net3550));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_102_clk_i_regs (.I(clknet_6_57__leaf_clk_i_regs),
    .Z(clknet_leaf_102_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 place3547 (.I(net528),
    .Z(net3547));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_58_clk_i_regs (.I(clknet_6_61__leaf_clk_i_regs),
    .Z(clknet_leaf_58_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place3546 (.I(net435),
    .Z(net3546));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3540 (.I(net423),
    .Z(net3540));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3647 (.I(net3646),
    .Z(net3647));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3646 (.I(\id_stage_i.controller_i.instr_i[14] ),
    .Z(net3646));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place3549 (.I(net314),
    .Z(net3549));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3569 (.I(net3558),
    .Z(net3569));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3545 (.I(net3543),
    .Z(net3545));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3544 (.I(net3543),
    .Z(net3544));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place3543 (.I(net3541),
    .Z(net3543));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3548 (.I(net423),
    .Z(net3548));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 place3541 (.I(net3513),
    .Z(net3541));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3542 (.I(net3541),
    .Z(net3542));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3659 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Z(net3659));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3567 (.I(net3558),
    .Z(net3567));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place3631 (.I(net418),
    .Z(net3631));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3087 (.I(_03831_),
    .Z(net3087));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3630 (.I(net449),
    .Z(net3630));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3650 (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(net3650));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3629 (.I(net3624),
    .Z(net3629));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3657 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Z(net3657));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3628 (.I(net3624),
    .Z(net3628));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3570 (.I(net3569),
    .Z(net3570));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3627 (.I(net3624),
    .Z(net3627));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22915__4 (.ZN(net253));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3083 (.I(_02019_),
    .Z(net3083));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3099 (.I(_03553_),
    .Z(net3099));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3075 (.I(_03797_),
    .Z(net3075));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3073 (.I(_03941_),
    .Z(net3073));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place3626 (.I(net3624),
    .Z(net3626));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3072 (.I(_05080_),
    .Z(net3072));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3112 (.I(_11301_[0]),
    .Z(net3112));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3575 (.I(net3574),
    .Z(net3575));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3574 (.I(net3558),
    .Z(net3574));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3069 (.I(_05115_),
    .Z(net3069));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3111 (.I(_03453_),
    .Z(net3111));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3061 (.I(_03982_),
    .Z(net3061));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3667 (.I(net142),
    .Z(net3667));
 gf180mcu_fd_sc_mcu9t5v0__tiel ibex_core_1 (.ZN(net250));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3064 (.I(_03760_),
    .Z(net3064));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3078 (.I(_03977_),
    .Z(net3078));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3068 (.I(_05329_),
    .Z(net3068));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3110 (.I(net3109),
    .Z(net3110));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place3063 (.I(_03785_),
    .Z(net3063));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3666 (.I(net143),
    .Z(net3666));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3070 (.I(_05115_),
    .Z(net3070));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place3051 (.I(_03813_),
    .Z(net3051));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3059 (.I(_05101_),
    .Z(net3059));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 place3050 (.I(net460),
    .Z(net3050));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3677 (.I(net131),
    .Z(net3677));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3675 (.I(net133),
    .Z(net3675));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3674 (.I(net134),
    .Z(net3674));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3654 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .Z(net3654));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3661 (.I(net148),
    .Z(net3661));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3656 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Z(net3656));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place3658 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Z(net3658));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place3660 (.I(net148),
    .Z(net3660));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place3573 (.I(net3569),
    .Z(net3573));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3572 (.I(net3569),
    .Z(net3572));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3673 (.I(net136),
    .Z(net3673));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3668 (.I(net141),
    .Z(net3668));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3672 (.I(net137),
    .Z(net3672));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3671 (.I(net138),
    .Z(net3671));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 place3676 (.I(net132),
    .Z(net3676));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_468_clk_i_regs (.I(clknet_6_30__leaf_clk_i_regs),
    .Z(clknet_leaf_468_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_469_clk_i_regs (.I(clknet_6_31__leaf_clk_i_regs),
    .Z(clknet_leaf_469_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_470_clk_i_regs (.I(clknet_6_31__leaf_clk_i_regs),
    .Z(clknet_leaf_470_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_473_clk_i_regs (.I(clknet_6_31__leaf_clk_i_regs),
    .Z(clknet_leaf_473_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_476_clk_i_regs (.I(clknet_6_30__leaf_clk_i_regs),
    .Z(clknet_leaf_476_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_478_clk_i_regs (.I(clknet_6_29__leaf_clk_i_regs),
    .Z(clknet_leaf_478_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_480_clk_i_regs (.I(clknet_6_28__leaf_clk_i_regs),
    .Z(clknet_leaf_480_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_483_clk_i_regs (.I(clknet_6_28__leaf_clk_i_regs),
    .Z(clknet_leaf_483_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_484_clk_i_regs (.I(clknet_6_30__leaf_clk_i_regs),
    .Z(clknet_leaf_484_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_486_clk_i_regs (.I(clknet_6_26__leaf_clk_i_regs),
    .Z(clknet_leaf_486_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_488_clk_i_regs (.I(clknet_6_26__leaf_clk_i_regs),
    .Z(clknet_leaf_488_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_492_clk_i_regs (.I(clknet_6_28__leaf_clk_i_regs),
    .Z(clknet_leaf_492_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_493_clk_i_regs (.I(clknet_6_28__leaf_clk_i_regs),
    .Z(clknet_leaf_493_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_494_clk_i_regs (.I(clknet_6_28__leaf_clk_i_regs),
    .Z(clknet_leaf_494_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_495_clk_i_regs (.I(clknet_6_28__leaf_clk_i_regs),
    .Z(clknet_leaf_495_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_497_clk_i_regs (.I(clknet_6_22__leaf_clk_i_regs),
    .Z(clknet_leaf_497_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_498_clk_i_regs (.I(clknet_6_22__leaf_clk_i_regs),
    .Z(clknet_leaf_498_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_501_clk_i_regs (.I(clknet_6_20__leaf_clk_i_regs),
    .Z(clknet_leaf_501_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_503_clk_i_regs (.I(clknet_6_21__leaf_clk_i_regs),
    .Z(clknet_leaf_503_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_507_clk_i_regs (.I(clknet_6_21__leaf_clk_i_regs),
    .Z(clknet_leaf_507_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_510_clk_i_regs (.I(clknet_6_21__leaf_clk_i_regs),
    .Z(clknet_leaf_510_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_512_clk_i_regs (.I(clknet_6_21__leaf_clk_i_regs),
    .Z(clknet_leaf_512_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_513_clk_i_regs (.I(clknet_6_26__leaf_clk_i_regs),
    .Z(clknet_leaf_513_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_514_clk_i_regs (.I(clknet_6_26__leaf_clk_i_regs),
    .Z(clknet_leaf_514_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_516_clk_i_regs (.I(clknet_6_26__leaf_clk_i_regs),
    .Z(clknet_leaf_516_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_517_clk_i_regs (.I(clknet_6_25__leaf_clk_i_regs),
    .Z(clknet_leaf_517_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_518_clk_i_regs (.I(clknet_6_25__leaf_clk_i_regs),
    .Z(clknet_leaf_518_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_522_clk_i_regs (.I(clknet_6_19__leaf_clk_i_regs),
    .Z(clknet_leaf_522_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_523_clk_i_regs (.I(clknet_6_19__leaf_clk_i_regs),
    .Z(clknet_leaf_523_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_525_clk_i_regs (.I(clknet_6_18__leaf_clk_i_regs),
    .Z(clknet_leaf_525_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_526_clk_i_regs (.I(clknet_6_19__leaf_clk_i_regs),
    .Z(clknet_leaf_526_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_528_clk_i_regs (.I(clknet_6_24__leaf_clk_i_regs),
    .Z(clknet_leaf_528_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_531_clk_i_regs (.I(clknet_6_18__leaf_clk_i_regs),
    .Z(clknet_leaf_531_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_532_clk_i_regs (.I(clknet_6_24__leaf_clk_i_regs),
    .Z(clknet_leaf_532_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_533_clk_i_regs (.I(clknet_6_18__leaf_clk_i_regs),
    .Z(clknet_leaf_533_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_535_clk_i_regs (.I(clknet_6_18__leaf_clk_i_regs),
    .Z(clknet_leaf_535_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_536_clk_i_regs (.I(clknet_6_18__leaf_clk_i_regs),
    .Z(clknet_leaf_536_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_537_clk_i_regs (.I(clknet_6_18__leaf_clk_i_regs),
    .Z(clknet_leaf_537_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_540_clk_i_regs (.I(clknet_6_16__leaf_clk_i_regs),
    .Z(clknet_leaf_540_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_543_clk_i_regs (.I(clknet_6_16__leaf_clk_i_regs),
    .Z(clknet_leaf_543_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_544_clk_i_regs (.I(clknet_6_16__leaf_clk_i_regs),
    .Z(clknet_leaf_544_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_546_clk_i_regs (.I(clknet_6_16__leaf_clk_i_regs),
    .Z(clknet_leaf_546_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_547_clk_i_regs (.I(clknet_6_16__leaf_clk_i_regs),
    .Z(clknet_leaf_547_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_548_clk_i_regs (.I(clknet_6_17__leaf_clk_i_regs),
    .Z(clknet_leaf_548_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_549_clk_i_regs (.I(clknet_6_17__leaf_clk_i_regs),
    .Z(clknet_leaf_549_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_550_clk_i_regs (.I(clknet_6_17__leaf_clk_i_regs),
    .Z(clknet_leaf_550_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_551_clk_i_regs (.I(clknet_6_17__leaf_clk_i_regs),
    .Z(clknet_leaf_551_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_556_clk_i_regs (.I(clknet_6_17__leaf_clk_i_regs),
    .Z(clknet_leaf_556_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_557_clk_i_regs (.I(clknet_6_21__leaf_clk_i_regs),
    .Z(clknet_leaf_557_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_558_clk_i_regs (.I(clknet_6_20__leaf_clk_i_regs),
    .Z(clknet_leaf_558_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_559_clk_i_regs (.I(clknet_6_20__leaf_clk_i_regs),
    .Z(clknet_leaf_559_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_560_clk_i_regs (.I(clknet_6_20__leaf_clk_i_regs),
    .Z(clknet_leaf_560_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_561_clk_i_regs (.I(clknet_6_20__leaf_clk_i_regs),
    .Z(clknet_leaf_561_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_563_clk_i_regs (.I(clknet_6_20__leaf_clk_i_regs),
    .Z(clknet_leaf_563_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_565_clk_i_regs (.I(clknet_6_22__leaf_clk_i_regs),
    .Z(clknet_leaf_565_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_566_clk_i_regs (.I(clknet_6_23__leaf_clk_i_regs),
    .Z(clknet_leaf_566_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_571_clk_i_regs (.I(clknet_6_23__leaf_clk_i_regs),
    .Z(clknet_leaf_571_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk_i_regs (.I(clk_i_regs),
    .Z(clknet_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_0_0_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_3_0_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_1_0_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_3_1_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_2_0_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_3_2_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_3_0_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_3_3_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_4_0_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_3_4_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_5_0_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_3_5_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_6_0_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_3_6_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_7_0_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_3_7_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_0__f_clk_i_regs (.I(clknet_3_0_0_clk_i_regs),
    .Z(clknet_6_0__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_1__f_clk_i_regs (.I(clknet_3_0_0_clk_i_regs),
    .Z(clknet_6_1__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_2__f_clk_i_regs (.I(clknet_3_0_0_clk_i_regs),
    .Z(clknet_6_2__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_3__f_clk_i_regs (.I(clknet_3_0_0_clk_i_regs),
    .Z(clknet_6_3__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_4__f_clk_i_regs (.I(clknet_3_0_0_clk_i_regs),
    .Z(clknet_6_4__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_5__f_clk_i_regs (.I(clknet_3_0_0_clk_i_regs),
    .Z(clknet_6_5__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_6__f_clk_i_regs (.I(clknet_3_0_0_clk_i_regs),
    .Z(clknet_6_6__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_7__f_clk_i_regs (.I(clknet_3_0_0_clk_i_regs),
    .Z(clknet_6_7__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_8__f_clk_i_regs (.I(clknet_3_1_0_clk_i_regs),
    .Z(clknet_6_8__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_9__f_clk_i_regs (.I(clknet_3_1_0_clk_i_regs),
    .Z(clknet_6_9__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_10__f_clk_i_regs (.I(clknet_3_1_0_clk_i_regs),
    .Z(clknet_6_10__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_11__f_clk_i_regs (.I(clknet_3_1_0_clk_i_regs),
    .Z(clknet_6_11__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_12__f_clk_i_regs (.I(clknet_3_1_0_clk_i_regs),
    .Z(clknet_6_12__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_13__f_clk_i_regs (.I(clknet_3_1_0_clk_i_regs),
    .Z(clknet_6_13__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_14__f_clk_i_regs (.I(clknet_3_1_0_clk_i_regs),
    .Z(clknet_6_14__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_15__f_clk_i_regs (.I(clknet_3_1_0_clk_i_regs),
    .Z(clknet_6_15__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_16__f_clk_i_regs (.I(clknet_3_2_0_clk_i_regs),
    .Z(clknet_6_16__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_17__f_clk_i_regs (.I(clknet_3_2_0_clk_i_regs),
    .Z(clknet_6_17__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_18__f_clk_i_regs (.I(clknet_3_2_0_clk_i_regs),
    .Z(clknet_6_18__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_19__f_clk_i_regs (.I(clknet_3_2_0_clk_i_regs),
    .Z(clknet_6_19__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_20__f_clk_i_regs (.I(clknet_3_2_0_clk_i_regs),
    .Z(clknet_6_20__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_21__f_clk_i_regs (.I(clknet_3_2_0_clk_i_regs),
    .Z(clknet_6_21__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_22__f_clk_i_regs (.I(clknet_3_2_0_clk_i_regs),
    .Z(clknet_6_22__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_23__f_clk_i_regs (.I(clknet_3_2_0_clk_i_regs),
    .Z(clknet_6_23__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_24__f_clk_i_regs (.I(clknet_3_3_0_clk_i_regs),
    .Z(clknet_6_24__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_25__f_clk_i_regs (.I(clknet_3_3_0_clk_i_regs),
    .Z(clknet_6_25__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_26__f_clk_i_regs (.I(clknet_3_3_0_clk_i_regs),
    .Z(clknet_6_26__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_27__f_clk_i_regs (.I(clknet_3_3_0_clk_i_regs),
    .Z(clknet_6_27__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_28__f_clk_i_regs (.I(clknet_3_3_0_clk_i_regs),
    .Z(clknet_6_28__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_29__f_clk_i_regs (.I(clknet_3_3_0_clk_i_regs),
    .Z(clknet_6_29__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_30__f_clk_i_regs (.I(clknet_3_3_0_clk_i_regs),
    .Z(clknet_6_30__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_31__f_clk_i_regs (.I(clknet_3_3_0_clk_i_regs),
    .Z(clknet_6_31__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_32__f_clk_i_regs (.I(clknet_3_4_0_clk_i_regs),
    .Z(clknet_6_32__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_33__f_clk_i_regs (.I(clknet_3_4_0_clk_i_regs),
    .Z(clknet_6_33__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_34__f_clk_i_regs (.I(clknet_3_4_0_clk_i_regs),
    .Z(clknet_6_34__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_35__f_clk_i_regs (.I(clknet_3_4_0_clk_i_regs),
    .Z(clknet_6_35__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_36__f_clk_i_regs (.I(clknet_3_4_0_clk_i_regs),
    .Z(clknet_6_36__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_37__f_clk_i_regs (.I(clknet_3_4_0_clk_i_regs),
    .Z(clknet_6_37__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_38__f_clk_i_regs (.I(clknet_3_4_0_clk_i_regs),
    .Z(clknet_6_38__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_39__f_clk_i_regs (.I(clknet_3_4_0_clk_i_regs),
    .Z(clknet_6_39__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_40__f_clk_i_regs (.I(clknet_3_5_0_clk_i_regs),
    .Z(clknet_6_40__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_41__f_clk_i_regs (.I(clknet_3_5_0_clk_i_regs),
    .Z(clknet_6_41__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_42__f_clk_i_regs (.I(clknet_3_5_0_clk_i_regs),
    .Z(clknet_6_42__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_43__f_clk_i_regs (.I(clknet_3_5_0_clk_i_regs),
    .Z(clknet_6_43__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_44__f_clk_i_regs (.I(clknet_3_5_0_clk_i_regs),
    .Z(clknet_6_44__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_45__f_clk_i_regs (.I(clknet_3_5_0_clk_i_regs),
    .Z(clknet_6_45__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_46__f_clk_i_regs (.I(clknet_3_5_0_clk_i_regs),
    .Z(clknet_6_46__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_47__f_clk_i_regs (.I(clknet_3_5_0_clk_i_regs),
    .Z(clknet_6_47__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_48__f_clk_i_regs (.I(clknet_3_6_0_clk_i_regs),
    .Z(clknet_6_48__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_49__f_clk_i_regs (.I(clknet_3_6_0_clk_i_regs),
    .Z(clknet_6_49__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_50__f_clk_i_regs (.I(clknet_3_6_0_clk_i_regs),
    .Z(clknet_6_50__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_51__f_clk_i_regs (.I(clknet_3_6_0_clk_i_regs),
    .Z(clknet_6_51__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_52__f_clk_i_regs (.I(clknet_3_6_0_clk_i_regs),
    .Z(clknet_6_52__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_53__f_clk_i_regs (.I(clknet_3_6_0_clk_i_regs),
    .Z(clknet_6_53__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_54__f_clk_i_regs (.I(clknet_3_6_0_clk_i_regs),
    .Z(clknet_6_54__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_55__f_clk_i_regs (.I(clknet_3_6_0_clk_i_regs),
    .Z(clknet_6_55__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_56__f_clk_i_regs (.I(clknet_3_7_0_clk_i_regs),
    .Z(clknet_6_56__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_57__f_clk_i_regs (.I(clknet_3_7_0_clk_i_regs),
    .Z(clknet_6_57__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_58__f_clk_i_regs (.I(clknet_3_7_0_clk_i_regs),
    .Z(clknet_6_58__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_59__f_clk_i_regs (.I(clknet_3_7_0_clk_i_regs),
    .Z(clknet_6_59__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_60__f_clk_i_regs (.I(clknet_3_7_0_clk_i_regs),
    .Z(clknet_6_60__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_61__f_clk_i_regs (.I(clknet_3_7_0_clk_i_regs),
    .Z(clknet_6_61__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_62__f_clk_i_regs (.I(clknet_3_7_0_clk_i_regs),
    .Z(clknet_6_62__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_63__f_clk_i_regs (.I(clknet_3_7_0_clk_i_regs),
    .Z(clknet_6_63__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload0 (.I(clknet_6_0__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload1 (.I(clknet_6_1__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload2 (.I(clknet_6_3__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload3 (.I(clknet_6_4__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload4 (.I(clknet_6_5__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload5 (.I(clknet_6_6__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload6 (.I(clknet_6_7__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload7 (.I(clknet_6_9__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload8 (.I(clknet_6_10__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload9 (.I(clknet_6_11__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload10 (.I(clknet_6_12__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload11 (.I(clknet_6_13__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload12 (.I(clknet_6_14__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload13 (.I(clknet_6_15__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload14 (.I(clknet_6_16__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload15 (.I(clknet_6_17__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload16 (.I(clknet_6_18__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload17 (.I(clknet_6_19__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload18 (.I(clknet_6_21__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload19 (.I(clknet_6_22__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload20 (.I(clknet_6_23__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload21 (.I(clknet_6_24__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload22 (.I(clknet_6_25__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload23 (.I(clknet_6_27__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload24 (.I(clknet_6_28__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload25 (.I(clknet_6_29__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload26 (.I(clknet_6_30__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload27 (.I(clknet_6_31__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload28 (.I(clknet_6_33__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload29 (.I(clknet_6_34__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload30 (.I(clknet_6_35__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload31 (.I(clknet_6_36__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload32 (.I(clknet_6_37__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload33 (.I(clknet_6_38__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload34 (.I(clknet_6_39__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload35 (.I(clknet_6_40__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload36 (.I(clknet_6_41__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload37 (.I(clknet_6_42__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload38 (.I(clknet_6_44__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload39 (.I(clknet_6_45__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload40 (.I(clknet_6_46__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload41 (.I(clknet_6_47__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload42 (.I(clknet_6_48__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload43 (.I(clknet_6_49__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload44 (.I(clknet_6_50__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload45 (.I(clknet_6_51__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload46 (.I(clknet_6_52__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload47 (.I(clknet_6_54__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload48 (.I(clknet_6_55__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload49 (.I(clknet_6_56__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload50 (.I(clknet_6_57__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload51 (.I(clknet_6_58__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload52 (.I(clknet_6_59__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload53 (.I(clknet_6_60__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 clkload54 (.I(clknet_6_62__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload55 (.I(clknet_6_63__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload56 (.I(clknet_leaf_391_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload57 (.I(clknet_leaf_393_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload58 (.I(clknet_leaf_398_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload59 (.I(clknet_leaf_405_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload60 (.I(clknet_leaf_408_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload61 (.I(clknet_leaf_409_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload62 (.I(clknet_leaf_373_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload63 (.I(clknet_leaf_375_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload64 (.I(clknet_leaf_381_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload65 (.I(clknet_leaf_383_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload66 (.I(clknet_leaf_384_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload67 (.I(clknet_leaf_385_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload68 (.I(clknet_leaf_386_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload69 (.I(clknet_leaf_371_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload70 (.I(clknet_leaf_426_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload71 (.I(clknet_leaf_428_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload72 (.I(clknet_leaf_422_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload73 (.I(clknet_leaf_423_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload74 (.I(clknet_leaf_424_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload75 (.I(clknet_leaf_447_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload76 (.I(clknet_leaf_449_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload77 (.I(clknet_leaf_450_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload78 (.I(clknet_leaf_217_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload79 (.I(clknet_leaf_219_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload80 (.I(clknet_leaf_465_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload81 (.I(clknet_leaf_466_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload82 (.I(clknet_leaf_356_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload83 (.I(clknet_leaf_359_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload84 (.I(clknet_leaf_360_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload85 (.I(clknet_leaf_365_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload86 (.I(clknet_leaf_319_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload87 (.I(clknet_leaf_349_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload88 (.I(clknet_leaf_350_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload89 (.I(clknet_leaf_330_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload90 (.I(clknet_leaf_331_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload91 (.I(clknet_leaf_334_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload92 (.I(clknet_leaf_335_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload93 (.I(clknet_leaf_352_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload94 (.I(clknet_leaf_309_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload95 (.I(clknet_leaf_311_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload96 (.I(clknet_leaf_436_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload97 (.I(clknet_leaf_247_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload98 (.I(clknet_leaf_307_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload99 (.I(clknet_leaf_308_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload100 (.I(clknet_leaf_296_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload101 (.I(clknet_leaf_297_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload102 (.I(clknet_leaf_322_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload103 (.I(clknet_leaf_324_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload104 (.I(clknet_leaf_325_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload105 (.I(clknet_leaf_327_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload106 (.I(clknet_leaf_295_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload107 (.I(clknet_leaf_299_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload108 (.I(clknet_leaf_301_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload109 (.I(clknet_leaf_303_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload110 (.I(clknet_leaf_306_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload111 (.I(clknet_leaf_310_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload112 (.I(clknet_leaf_548_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload113 (.I(clknet_leaf_549_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload114 (.I(clknet_leaf_550_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload115 (.I(clknet_leaf_525_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload116 (.I(clknet_leaf_531_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload117 (.I(clknet_leaf_535_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload118 (.I(clknet_leaf_536_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload119 (.I(clknet_leaf_523_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload120 (.I(clknet_leaf_526_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload121 (.I(clknet_leaf_501_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload122 (.I(clknet_leaf_558_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload123 (.I(clknet_leaf_559_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload124 (.I(clknet_leaf_560_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload125 (.I(clknet_leaf_510_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload126 (.I(clknet_leaf_557_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload127 (.I(clknet_leaf_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload128 (.I(clknet_leaf_571_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload129 (.I(clknet_leaf_399_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload130 (.I(clknet_leaf_400_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload131 (.I(clknet_leaf_402_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload132 (.I(clknet_leaf_403_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload133 (.I(clknet_leaf_404_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload134 (.I(clknet_leaf_532_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload135 (.I(clknet_leaf_416_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload136 (.I(clknet_leaf_417_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload137 (.I(clknet_leaf_418_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload138 (.I(clknet_leaf_486_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload139 (.I(clknet_leaf_514_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload140 (.I(clknet_leaf_516_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload141 (.I(clknet_leaf_483_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload142 (.I(clknet_leaf_492_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload143 (.I(clknet_leaf_494_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload144 (.I(clknet_leaf_495_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload145 (.I(clknet_leaf_1_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload146 (.I(clknet_leaf_4_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload147 (.I(clknet_leaf_478_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload148 (.I(clknet_leaf_467_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload149 (.I(clknet_leaf_468_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload150 (.I(clknet_leaf_476_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload151 (.I(clknet_leaf_211_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload152 (.I(clknet_leaf_469_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload153 (.I(clknet_leaf_470_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload154 (.I(clknet_leaf_233_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload155 (.I(clknet_leaf_235_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload156 (.I(clknet_leaf_241_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload157 (.I(clknet_leaf_242_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload158 (.I(clknet_leaf_244_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload159 (.I(clknet_leaf_260_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload160 (.I(clknet_leaf_229_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload161 (.I(clknet_leaf_234_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload162 (.I(clknet_leaf_238_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload163 (.I(clknet_leaf_10_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload164 (.I(clknet_leaf_208_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload165 (.I(clknet_leaf_222_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload166 (.I(clknet_leaf_226_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload167 (.I(clknet_leaf_292_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload168 (.I(clknet_leaf_294_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload169 (.I(clknet_leaf_277_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload170 (.I(clknet_leaf_278_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload171 (.I(clknet_leaf_281_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload172 (.I(clknet_leaf_284_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload173 (.I(clknet_leaf_285_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload174 (.I(clknet_leaf_286_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload175 (.I(clknet_leaf_156_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload176 (.I(clknet_leaf_158_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload177 (.I(clknet_leaf_269_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload178 (.I(clknet_leaf_145_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload179 (.I(clknet_leaf_282_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload180 (.I(clknet_leaf_283_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload181 (.I(clknet_leaf_137_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload182 (.I(clknet_leaf_138_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload183 (.I(clknet_leaf_141_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload184 (.I(clknet_leaf_143_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkload185 (.I(clknet_leaf_11_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkload186 (.I(clknet_leaf_12_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkload187 (.I(clknet_leaf_186_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload188 (.I(clknet_leaf_191_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload189 (.I(clknet_leaf_13_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload190 (.I(clknet_leaf_15_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload191 (.I(clknet_leaf_180_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload192 (.I(clknet_leaf_17_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload193 (.I(clknet_leaf_18_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload194 (.I(clknet_leaf_22_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload195 (.I(clknet_leaf_36_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload196 (.I(clknet_leaf_23_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload197 (.I(clknet_leaf_27_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload198 (.I(clknet_leaf_28_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload199 (.I(clknet_leaf_29_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload200 (.I(clknet_leaf_34_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload201 (.I(clknet_leaf_38_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload202 (.I(clknet_leaf_40_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload203 (.I(clknet_leaf_102_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload204 (.I(clknet_leaf_108_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload205 (.I(clknet_leaf_109_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload206 (.I(clknet_leaf_110_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload207 (.I(clknet_leaf_113_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload208 (.I(clknet_leaf_177_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload209 (.I(clknet_leaf_128_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload210 (.I(clknet_leaf_129_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload211 (.I(clknet_leaf_134_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload212 (.I(clknet_leaf_136_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload213 (.I(clknet_leaf_139_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload214 (.I(clknet_leaf_47_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload215 (.I(clknet_leaf_49_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload216 (.I(clknet_leaf_97_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload217 (.I(clknet_leaf_98_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload218 (.I(clknet_leaf_100_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload219 (.I(clknet_leaf_48_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload220 (.I(clknet_leaf_57_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload221 (.I(clknet_leaf_60_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload222 (.I(clknet_leaf_65_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload223 (.I(clknet_leaf_67_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload224 (.I(clknet_leaf_68_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload225 (.I(clknet_leaf_74_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload226 (.I(clknet_leaf_77_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_23_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_25_clk (.I(clknet_6_12__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_27_clk (.I(clknet_6_18__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_29_clk (.I(clknet_6_18__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_32_clk (.I(clknet_6_24__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_33_clk (.I(clknet_6_24__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_34_clk (.I(clknet_6_24__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_35_clk (.I(clknet_6_18__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_37_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_38_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_40_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_41_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_42_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_44_clk (.I(clknet_6_13__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_45_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_48_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_52_clk (.I(clknet_6_27__leaf_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_53_clk (.I(clknet_6_25__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_54_clk (.I(clknet_6_27__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_56_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_57_clk (.I(clknet_6_27__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_58_clk (.I(clknet_6_27__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_61_clk (.I(clknet_6_15__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_64_clk (.I(clknet_6_15__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_66_clk (.I(clknet_6_15__leaf_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_71_clk (.I(clknet_6_15__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_72_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_73_clk (.I(clknet_6_15__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_74_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_78_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_84_clk (.I(clknet_6_36__leaf_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_85_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_88_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_91_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_93_clk (.I(clknet_6_33__leaf_clk),
    .Z(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_95_clk (.I(clknet_6_33__leaf_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_98_clk (.I(clknet_6_33__leaf_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_100_clk (.I(clknet_6_14__leaf_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_102_clk (.I(clknet_6_33__leaf_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_104_clk (.I(clknet_6_14__leaf_clk),
    .Z(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_107_clk (.I(clknet_6_14__leaf_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_109_clk (.I(clknet_6_14__leaf_clk),
    .Z(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_110_clk (.I(clknet_6_14__leaf_clk),
    .Z(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_117_clk (.I(clknet_6_11__leaf_clk),
    .Z(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_125_clk (.I(clknet_6_10__leaf_clk),
    .Z(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_127_clk (.I(clknet_6_10__leaf_clk),
    .Z(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_128_clk (.I(clknet_6_10__leaf_clk),
    .Z(clknet_leaf_128_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_129_clk (.I(clknet_6_32__leaf_clk),
    .Z(clknet_leaf_129_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_130_clk (.I(clknet_6_32__leaf_clk),
    .Z(clknet_leaf_130_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_131_clk (.I(clknet_6_32__leaf_clk),
    .Z(clknet_leaf_131_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_132_clk (.I(clknet_6_32__leaf_clk),
    .Z(clknet_leaf_132_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_135_clk (.I(clknet_6_32__leaf_clk),
    .Z(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_138_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_139_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_140_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_140_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_143_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_143_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_146_clk (.I(clknet_6_32__leaf_clk),
    .Z(clknet_leaf_146_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_149_clk (.I(clknet_6_34__leaf_clk),
    .Z(clknet_leaf_149_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_150_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_151_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_151_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_152_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_154_clk (.I(clknet_6_35__leaf_clk),
    .Z(clknet_leaf_154_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_155_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_155_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_156_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_157_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_157_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_160_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_160_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_161_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_161_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_162_clk (.I(clknet_6_40__leaf_clk),
    .Z(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_165_clk (.I(clknet_6_40__leaf_clk),
    .Z(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_167_clk (.I(clknet_6_40__leaf_clk),
    .Z(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_168_clk (.I(clknet_6_40__leaf_clk),
    .Z(clknet_leaf_168_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_173_clk (.I(clknet_6_40__leaf_clk),
    .Z(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_174_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_175_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_178_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_181_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_183_clk (.I(clknet_6_42__leaf_clk),
    .Z(clknet_leaf_183_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_186_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_188_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_188_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_191_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_192_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_192_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_195_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_195_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_197_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_198_clk (.I(clknet_6_43__leaf_clk),
    .Z(clknet_leaf_198_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_199_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_199_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_202_clk (.I(clknet_6_41__leaf_clk),
    .Z(clknet_leaf_202_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_206_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_206_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_207_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_207_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_209_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_211_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_213_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_214_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_215_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_218_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_218_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_220_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_220_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_224_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_225_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_225_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_226_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_228_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_228_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_229_clk (.I(clknet_6_46__leaf_clk),
    .Z(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_233_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_233_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_238_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_238_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_240_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_240_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_241_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_242_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_242_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_243_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_244_clk (.I(clknet_6_56__leaf_clk),
    .Z(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_247_clk (.I(clknet_6_47__leaf_clk),
    .Z(clknet_leaf_247_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_248_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_248_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_250_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_250_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_252_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_252_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_253_clk (.I(clknet_6_56__leaf_clk),
    .Z(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_255_clk (.I(clknet_6_56__leaf_clk),
    .Z(clknet_leaf_255_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_258_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_258_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_264_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_264_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_265_clk (.I(clknet_6_45__leaf_clk),
    .Z(clknet_leaf_265_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_266_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_266_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_267_clk (.I(clknet_6_44__leaf_clk),
    .Z(clknet_leaf_267_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_269_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_269_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_272_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_272_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_275_clk (.I(clknet_6_39__leaf_clk),
    .Z(clknet_leaf_275_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_277_clk (.I(clknet_6_38__leaf_clk),
    .Z(clknet_leaf_277_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_281_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_281_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_284_clk (.I(clknet_6_39__leaf_clk),
    .Z(clknet_leaf_284_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_286_clk (.I(clknet_6_39__leaf_clk),
    .Z(clknet_leaf_286_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_288_clk (.I(clknet_6_39__leaf_clk),
    .Z(clknet_leaf_288_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_293_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_293_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_296_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_296_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_297_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_297_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_298_clk (.I(clknet_6_37__leaf_clk),
    .Z(clknet_leaf_298_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_307_clk (.I(clknet_6_48__leaf_clk),
    .Z(clknet_leaf_307_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_312_clk (.I(clknet_6_48__leaf_clk),
    .Z(clknet_leaf_312_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_323_clk (.I(clknet_6_50__leaf_clk),
    .Z(clknet_leaf_323_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_328_clk (.I(clknet_6_51__leaf_clk),
    .Z(clknet_leaf_328_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_331_clk (.I(clknet_6_51__leaf_clk),
    .Z(clknet_leaf_331_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_332_clk (.I(clknet_6_51__leaf_clk),
    .Z(clknet_leaf_332_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_335_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_335_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_336_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_336_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_344_clk (.I(clknet_6_56__leaf_clk),
    .Z(clknet_leaf_344_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_345_clk (.I(clknet_6_56__leaf_clk),
    .Z(clknet_leaf_345_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_351_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_351_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_352_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_352_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_353_clk (.I(clknet_6_56__leaf_clk),
    .Z(clknet_leaf_353_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_354_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_354_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_358_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_358_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_360_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_360_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_361_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_361_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_363_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_363_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_364_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_364_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_365_clk (.I(clknet_6_58__leaf_clk),
    .Z(clknet_leaf_365_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_366_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_366_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_372_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_372_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_375_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_375_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_376_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_376_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_377_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_377_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_378_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_378_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_382_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_382_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_383_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_383_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_384_clk (.I(clknet_6_59__leaf_clk),
    .Z(clknet_leaf_384_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_385_clk (.I(clknet_6_57__leaf_clk),
    .Z(clknet_leaf_385_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_390_clk (.I(clknet_6_51__leaf_clk),
    .Z(clknet_leaf_390_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_398_clk (.I(clknet_6_54__leaf_clk),
    .Z(clknet_leaf_398_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_401_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_401_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_403_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_403_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_406_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_406_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_407_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_407_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_408_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_408_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_409_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_409_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_410_clk (.I(clknet_6_63__leaf_clk),
    .Z(clknet_leaf_410_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_413_clk (.I(clknet_6_62__leaf_clk),
    .Z(clknet_leaf_413_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_420_clk (.I(clknet_6_63__leaf_clk),
    .Z(clknet_leaf_420_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_423_clk (.I(clknet_6_63__leaf_clk),
    .Z(clknet_leaf_423_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_425_clk (.I(clknet_6_63__leaf_clk),
    .Z(clknet_leaf_425_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_426_clk (.I(clknet_6_63__leaf_clk),
    .Z(clknet_leaf_426_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_427_clk (.I(clknet_6_63__leaf_clk),
    .Z(clknet_leaf_427_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_428_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_428_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_436_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_436_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_437_clk (.I(clknet_6_61__leaf_clk),
    .Z(clknet_leaf_437_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_440_clk (.I(clknet_6_60__leaf_clk),
    .Z(clknet_leaf_440_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_452_clk (.I(clknet_6_53__leaf_clk),
    .Z(clknet_leaf_452_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_455_clk (.I(clknet_6_53__leaf_clk),
    .Z(clknet_leaf_455_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_459_clk (.I(clknet_6_53__leaf_clk),
    .Z(clknet_leaf_459_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_468_clk (.I(clknet_6_52__leaf_clk),
    .Z(clknet_leaf_468_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_475_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_475_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_476_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_476_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_479_clk (.I(clknet_6_31__leaf_clk),
    .Z(clknet_leaf_479_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_485_clk (.I(clknet_6_30__leaf_clk),
    .Z(clknet_leaf_485_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_486_clk (.I(clknet_6_31__leaf_clk),
    .Z(clknet_leaf_486_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_489_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_489_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_494_clk (.I(clknet_6_29__leaf_clk),
    .Z(clknet_leaf_494_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_495_clk (.I(clknet_6_28__leaf_clk),
    .Z(clknet_leaf_495_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_497_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_497_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_498_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_498_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_499_clk (.I(clknet_6_21__leaf_clk),
    .Z(clknet_leaf_499_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_501_clk (.I(clknet_6_21__leaf_clk),
    .Z(clknet_leaf_501_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_502_clk (.I(clknet_6_21__leaf_clk),
    .Z(clknet_leaf_502_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_503_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_503_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_504_clk (.I(clknet_6_23__leaf_clk),
    .Z(clknet_leaf_504_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_511_clk (.I(clknet_6_26__leaf_clk),
    .Z(clknet_leaf_511_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_514_clk (.I(clknet_6_22__leaf_clk),
    .Z(clknet_leaf_514_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_515_clk (.I(clknet_6_19__leaf_clk),
    .Z(clknet_leaf_515_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_520_clk (.I(clknet_6_19__leaf_clk),
    .Z(clknet_leaf_520_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_521_clk (.I(clknet_6_19__leaf_clk),
    .Z(clknet_leaf_521_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_522_clk (.I(clknet_6_19__leaf_clk),
    .Z(clknet_leaf_522_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_528_clk (.I(clknet_6_18__leaf_clk),
    .Z(clknet_leaf_528_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_530_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_530_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_531_clk (.I(clknet_6_16__leaf_clk),
    .Z(clknet_leaf_531_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_532_clk (.I(clknet_6_16__leaf_clk),
    .Z(clknet_leaf_532_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_533_clk (.I(clknet_6_16__leaf_clk),
    .Z(clknet_leaf_533_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_534_clk (.I(clknet_6_17__leaf_clk),
    .Z(clknet_leaf_534_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_537_clk (.I(clknet_6_22__leaf_clk),
    .Z(clknet_leaf_537_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_539_clk (.I(clknet_6_22__leaf_clk),
    .Z(clknet_leaf_539_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_540_clk (.I(clknet_6_22__leaf_clk),
    .Z(clknet_leaf_540_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_543_clk (.I(clknet_6_22__leaf_clk),
    .Z(clknet_leaf_543_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_544_clk (.I(clknet_6_20__leaf_clk),
    .Z(clknet_leaf_544_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_546_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_546_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_549_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_549_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_550_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_550_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_552_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_552_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_553_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_553_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_555_clk (.I(clknet_6_5__leaf_clk),
    .Z(clknet_leaf_555_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_559_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_559_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_560_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_560_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_564_clk (.I(clknet_6_7__leaf_clk),
    .Z(clknet_leaf_564_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_567_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_567_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_569_clk (.I(clknet_6_3__leaf_clk),
    .Z(clknet_leaf_569_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_570_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_570_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_571_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_571_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_572_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_572_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_573_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_573_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_575_clk (.I(clknet_6_6__leaf_clk),
    .Z(clknet_leaf_575_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_580_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_580_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_583_clk (.I(clknet_6_4__leaf_clk),
    .Z(clknet_leaf_583_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_584_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_584_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_587_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_587_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_588_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_588_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_589_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_589_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_590_clk (.I(clknet_6_1__leaf_clk),
    .Z(clknet_leaf_590_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_592_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_592_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_593_clk (.I(clknet_6_3__leaf_clk),
    .Z(clknet_leaf_593_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_594_clk (.I(clknet_6_0__leaf_clk),
    .Z(clknet_leaf_594_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_601_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_601_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_608_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_608_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_609_clk (.I(clknet_6_2__leaf_clk),
    .Z(clknet_leaf_609_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_610_clk (.I(clknet_6_9__leaf_clk),
    .Z(clknet_leaf_610_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_611_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_611_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_612_clk (.I(clknet_6_8__leaf_clk),
    .Z(clknet_leaf_612_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_620_clk (.I(clknet_6_11__leaf_clk),
    .Z(clknet_leaf_620_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_3_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_0__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_6_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_1__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_6_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_2__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_6_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_3__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_6_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_4__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_6_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_5__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_6_5__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_6__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_6_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_7__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_6_7__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_8__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_6_8__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_9__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_6_9__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_10__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_6_10__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_11__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_6_11__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_12__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_6_12__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_13__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_6_13__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_14__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_6_14__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_15__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_6_15__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_16__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_6_16__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_17__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_6_17__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_18__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_6_18__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_19__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_6_19__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_20__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_6_20__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_21__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_6_21__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_22__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_6_22__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_23__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_6_23__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_24__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_6_24__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_25__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_6_25__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_26__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_6_26__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_27__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_6_27__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_28__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_6_28__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_29__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_6_29__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_30__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_6_30__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_31__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_6_31__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_32__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_6_32__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_33__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_6_33__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_34__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_6_34__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_35__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_6_35__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_36__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_6_36__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_37__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_6_37__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_38__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_6_38__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_39__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_6_39__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_40__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_6_40__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_41__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_6_41__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_42__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_6_42__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_43__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_6_43__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_44__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_6_44__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_45__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_6_45__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_46__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_6_46__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_47__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_6_47__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_48__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_6_48__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_49__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_6_49__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_50__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_6_50__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_51__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_6_51__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_52__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_6_52__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_53__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_6_53__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_54__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_6_54__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_55__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_6_55__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_56__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_6_56__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_57__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_6_57__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_58__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_6_58__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_59__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_6_59__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_60__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_6_60__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_61__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_6_61__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_62__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_6_62__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_6_63__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_6_63__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload227 (.I(clknet_6_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_12 clkload228 (.I(clknet_6_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload229 (.I(clknet_6_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload230 (.I(clknet_6_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload231 (.I(clknet_6_4__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload232 (.I(clknet_6_6__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload233 (.I(clknet_6_7__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload234 (.I(clknet_6_8__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload235 (.I(clknet_6_9__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload236 (.I(clknet_6_10__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload237 (.I(clknet_6_11__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload238 (.I(clknet_6_12__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload239 (.I(clknet_6_14__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_16 clkload240 (.I(clknet_6_15__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload241 (.I(clknet_6_16__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload242 (.I(clknet_6_17__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload243 (.I(clknet_6_18__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload244 (.I(clknet_6_19__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload245 (.I(clknet_6_20__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload246 (.I(clknet_6_21__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload247 (.I(clknet_6_23__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload248 (.I(clknet_6_24__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload249 (.I(clknet_6_25__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload250 (.I(clknet_6_26__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload251 (.I(clknet_6_28__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload252 (.I(clknet_6_29__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload253 (.I(clknet_6_30__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload254 (.I(clknet_6_31__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload255 (.I(clknet_6_32__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload256 (.I(clknet_6_33__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload257 (.I(clknet_6_34__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload258 (.I(clknet_6_35__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload259 (.I(clknet_6_36__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload260 (.I(clknet_6_37__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload261 (.I(clknet_6_39__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload262 (.I(clknet_6_40__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 clkload263 (.I(clknet_6_41__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload264 (.I(clknet_6_42__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload265 (.I(clknet_6_43__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload266 (.I(clknet_6_44__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload267 (.I(clknet_6_45__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkload268 (.I(clknet_6_46__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload269 (.I(clknet_6_48__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload270 (.I(clknet_6_49__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload271 (.I(clknet_6_50__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload272 (.I(clknet_6_52__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload273 (.I(clknet_6_53__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload274 (.I(clknet_6_54__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload275 (.I(clknet_6_55__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload276 (.I(clknet_6_56__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload277 (.I(clknet_6_57__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload278 (.I(clknet_6_59__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload279 (.I(clknet_6_60__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload280 (.I(clknet_6_61__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload281 (.I(clknet_6_62__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload282 (.I(clknet_6_63__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload283 (.I(clknet_leaf_571_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload284 (.I(clknet_leaf_584_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload285 (.I(clknet_leaf_587_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload286 (.I(clknet_leaf_589_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload287 (.I(clknet_leaf_601_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload288 (.I(clknet_leaf_608_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload289 (.I(clknet_leaf_609_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload290 (.I(clknet_leaf_572_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload291 (.I(clknet_leaf_573_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload292 (.I(clknet_leaf_583_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload293 (.I(clknet_leaf_567_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload294 (.I(clknet_leaf_570_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload295 (.I(clknet_leaf_575_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload296 (.I(clknet_leaf_611_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload297 (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload298 (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload299 (.I(clknet_leaf_610_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload300 (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload301 (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload302 (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload303 (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload304 (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload305 (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload306 (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload307 (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload308 (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload309 (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload310 (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload311 (.I(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload312 (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload313 (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload314 (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload315 (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload316 (.I(clknet_leaf_528_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload317 (.I(clknet_leaf_515_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload318 (.I(clknet_leaf_520_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload319 (.I(clknet_leaf_521_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload320 (.I(clknet_leaf_498_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload321 (.I(clknet_leaf_503_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload322 (.I(clknet_leaf_544_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload323 (.I(clknet_leaf_501_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload324 (.I(clknet_leaf_502_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload325 (.I(clknet_leaf_514_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload326 (.I(clknet_leaf_537_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload327 (.I(clknet_leaf_539_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload328 (.I(clknet_leaf_540_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload329 (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload330 (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload331 (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload332 (.I(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload333 (.I(clknet_leaf_511_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload334 (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload335 (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload336 (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload337 (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload338 (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload339 (.I(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload340 (.I(clknet_leaf_151_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload341 (.I(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload342 (.I(clknet_leaf_154_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload343 (.I(clknet_leaf_281_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload344 (.I(clknet_leaf_293_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload345 (.I(clknet_leaf_296_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload346 (.I(clknet_leaf_297_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload347 (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload348 (.I(clknet_leaf_266_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload349 (.I(clknet_leaf_269_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload350 (.I(clknet_leaf_272_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload351 (.I(clknet_leaf_277_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload352 (.I(clknet_leaf_275_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload353 (.I(clknet_leaf_284_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload354 (.I(clknet_leaf_286_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload355 (.I(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload356 (.I(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload357 (.I(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload358 (.I(clknet_leaf_168_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload359 (.I(clknet_leaf_155_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload360 (.I(clknet_leaf_157_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload361 (.I(clknet_leaf_161_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload362 (.I(clknet_leaf_199_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload363 (.I(clknet_leaf_202_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload364 (.I(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload365 (.I(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload366 (.I(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload367 (.I(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload368 (.I(clknet_leaf_192_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload369 (.I(clknet_leaf_195_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload370 (.I(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload371 (.I(clknet_leaf_206_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload372 (.I(clknet_leaf_207_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload373 (.I(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload374 (.I(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload375 (.I(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload376 (.I(clknet_leaf_267_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload377 (.I(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload378 (.I(clknet_leaf_248_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload379 (.I(clknet_leaf_250_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload380 (.I(clknet_leaf_252_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload381 (.I(clknet_leaf_258_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload382 (.I(clknet_leaf_188_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload383 (.I(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload384 (.I(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload385 (.I(clknet_leaf_218_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload386 (.I(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload387 (.I(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload388 (.I(clknet_leaf_225_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload389 (.I(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload390 (.I(clknet_leaf_228_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload391 (.I(clknet_leaf_233_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload392 (.I(clknet_leaf_247_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload393 (.I(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload394 (.I(clknet_leaf_253_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload395 (.I(clknet_leaf_255_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload396 (.I(clknet_leaf_345_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload397 (.I(clknet_leaf_353_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload398 (.I(clknet_leaf_335_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload399 (.I(clknet_leaf_351_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload400 (.I(clknet_leaf_352_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload401 (.I(clknet_leaf_383_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload402 (.I(clknet_leaf_385_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload403 (.I(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload404 (.I(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload405 (.I(clknet_leaf_354_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload406 (.I(clknet_leaf_360_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload407 (.I(clknet_leaf_361_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload408 (.I(clknet_leaf_363_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload409 (.I(clknet_leaf_364_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload410 (.I(clknet_leaf_365_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload411 (.I(clknet_leaf_366_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload412 (.I(clknet_leaf_372_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload413 (.I(clknet_leaf_375_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload414 (.I(clknet_leaf_376_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload415 (.I(clknet_leaf_378_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload416 (.I(clknet_leaf_384_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload417 (.I(clknet_leaf_403_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload418 (.I(clknet_leaf_406_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload419 (.I(clknet_leaf_408_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload420 (.I(clknet_leaf_409_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload421 (.I(clknet_leaf_410_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload422 (.I(clknet_leaf_423_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload423 (.I(clknet_leaf_425_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload424 (.I(clknet_leaf_427_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_0_core_clock (.I(delaynet_0_core_clock),
    .Z(delaynet_1_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_1_core_clock (.I(delaynet_1_core_clock),
    .Z(delaynet_2_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_2_core_clock (.I(delaynet_2_core_clock),
    .Z(delaynet_3_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_3_core_clock (.I(delaynet_3_core_clock),
    .Z(clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer1 (.I(net172),
    .Z(net256));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer2 (.I(net172),
    .Z(net257));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer3 (.I(net172),
    .Z(net258));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer4 (.I(_08248_),
    .Z(net259));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer5 (.I(net317),
    .Z(net260));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer6 (.I(_06254_),
    .Z(net261));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer7 (.I(net344),
    .Z(net262));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer8 (.I(_11391_[0]),
    .Z(net263));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer9 (.I(_11391_[0]),
    .Z(net264));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer10 (.I(_06202_),
    .Z(net265));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer11 (.I(net265),
    .Z(net266));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 clone12 (.A1(_07012_),
    .A2(net283),
    .ZN(net267));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer13 (.I(_06198_),
    .Z(net268));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer14 (.I(_06198_),
    .Z(net269));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer15 (.I(net269),
    .Z(net270));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer16 (.I(_11077_[0]),
    .Z(net271));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer17 (.I(_07195_),
    .Z(net272));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer18 (.I(_08253_),
    .Z(net273));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer19 (.I(_06214_),
    .Z(net274));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer20 (.I(\id_stage_i.id_fsm_q ),
    .Z(net275));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 rebuffer21 (.I(_06437_),
    .Z(net276));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer22 (.I(\id_stage_i.controller_i.instr_i[6] ),
    .Z(net277));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer23 (.I(_07195_),
    .Z(net278));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer24 (.I(net3094),
    .Z(net279));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer25 (.I(net3094),
    .Z(net280));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer26 (.I(_11057_[0]),
    .Z(net281));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone27 (.I(net285),
    .Z(net282));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer28 (.I(_07009_),
    .Z(net283));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer29 (.I(_07255_),
    .Z(net284));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer30 (.I(_07013_),
    .Z(net285));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer31 (.I(_07304_),
    .Z(net286));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer32 (.I(_07304_),
    .Z(net287));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer33 (.I(_11041_[0]),
    .Z(net288));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer34 (.I(net166),
    .Z(net289));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer35 (.I(_06997_),
    .Z(net290));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone36 (.A1(net3190),
    .A2(net450),
    .B(_03927_),
    .ZN(net291));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer37 (.I(_11033_[0]),
    .Z(net292));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer38 (.I(_11049_[0]),
    .Z(net293));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer39 (.I(_11049_[0]),
    .Z(net294));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer40 (.I(net173),
    .Z(net295));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer41 (.I(net173),
    .Z(net296));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer42 (.I(_08254_),
    .Z(net297));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer43 (.I(_11007_[0]),
    .Z(net298));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer44 (.I(_06953_),
    .Z(net299));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer45 (.I(_06954_),
    .Z(net300));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer46 (.I(_06387_),
    .Z(net301));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer47 (.I(_06387_),
    .Z(net302));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer48 (.I(\id_stage_i.controller_i.instr_i[13] ),
    .Z(net303));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer49 (.I(\id_stage_i.controller_i.instr_i[13] ),
    .Z(net304));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clone50 (.I(net306),
    .Z(net305));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer51 (.I(net307),
    .Z(net306));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer52 (.I(_07009_),
    .Z(net307));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer53 (.I(_11025_[0]),
    .Z(net308));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer54 (.I(net3195),
    .Z(net309));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer55 (.I(_11045_[0]),
    .Z(net310));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer56 (.I(_11045_[0]),
    .Z(net311));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer57 (.I(_11045_[0]),
    .Z(net312));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer200 (.I(_06440_),
    .Z(net484));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clone59 (.I(net440),
    .Z(net314));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer60 (.I(_11053_[0]),
    .Z(net315));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer61 (.I(_07683_),
    .Z(net316));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer62 (.I(net267),
    .Z(net317));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer63 (.I(_07283_),
    .Z(net318));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer64 (.I(_07283_),
    .Z(net319));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone65 (.I(net356),
    .Z(net320));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer66 (.I(_06212_),
    .Z(net321));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer67 (.I(_06212_),
    .Z(net322));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer68 (.I(_06212_),
    .Z(net323));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer69 (.I(_06780_),
    .Z(net324));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer70 (.I(_06780_),
    .Z(net325));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer71 (.I(_06780_),
    .Z(net326));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer72 (.I(net326),
    .Z(net327));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer73 (.I(_06749_),
    .Z(net328));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer74 (.I(_06439_),
    .Z(net329));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer75 (.I(_06526_),
    .Z(net330));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer76 (.I(_06526_),
    .Z(net331));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer77 (.I(_06996_),
    .Z(net332));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 clone78 (.I(net452),
    .Z(net333));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer79 (.I(_06384_),
    .Z(net334));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer81 (.I(_05038_),
    .Z(net336));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer82 (.I(net170),
    .Z(net337));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer83 (.I(net170),
    .Z(net338));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer84 (.I(net170),
    .Z(net339));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer85 (.I(_05016_),
    .Z(net340));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer86 (.I(_06577_),
    .Z(net341));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer87 (.I(net341),
    .Z(net342));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer91 (.I(_04997_),
    .Z(net346));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer92 (.I(_08078_),
    .Z(net347));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer93 (.I(_11061_[0]),
    .Z(net348));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer94 (.I(_07258_),
    .Z(net349));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer95 (.I(_07197_),
    .Z(net350));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer96 (.I(_07191_),
    .Z(net351));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer97 (.I(_07508_),
    .Z(net352));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer98 (.I(_06966_),
    .Z(net353));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer99 (.I(\id_stage_i.controller_i.instr_i[6] ),
    .Z(net354));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer100 (.I(\id_stage_i.controller_i.instr_i[6] ),
    .Z(net355));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer101 (.I(\id_stage_i.controller_i.instr_i[12] ),
    .Z(net356));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer102 (.I(\id_stage_i.controller_i.instr_i[5] ),
    .Z(net357));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer103 (.I(_04987_),
    .Z(net358));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer104 (.I(_07396_),
    .Z(net359));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer105 (.I(net159),
    .Z(net360));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer106 (.I(net159),
    .Z(net361));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer107 (.I(_04862_),
    .Z(net362));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer108 (.I(_04862_),
    .Z(net363));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer109 (.I(net3097),
    .Z(net364));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer110 (.I(net3097),
    .Z(net365));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer111 (.I(net168),
    .Z(net366));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer112 (.I(net168),
    .Z(net367));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer113 (.I(net168),
    .Z(net368));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer117 (.I(net164),
    .Z(net372));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer118 (.I(net164),
    .Z(net373));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer119 (.I(_07246_),
    .Z(net374));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer120 (.I(_04953_),
    .Z(net375));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer121 (.I(net165),
    .Z(net376));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer122 (.I(net165),
    .Z(net377));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer123 (.I(_07793_),
    .Z(net378));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer124 (.I(_07601_),
    .Z(net379));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer125 (.I(_04962_),
    .Z(net380));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer126 (.I(_04962_),
    .Z(net381));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer127 (.I(_11021_[0]),
    .Z(net382));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer131 (.I(_07797_),
    .Z(net386));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer132 (.I(_08160_),
    .Z(net387));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer136 (.I(_04932_),
    .Z(net391));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer137 (.I(_04931_),
    .Z(net392));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer147 (.I(net157),
    .Z(net402));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer148 (.I(net157),
    .Z(net403));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer149 (.I(net157),
    .Z(net404));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer150 (.I(_04882_),
    .Z(net405));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer151 (.I(_04882_),
    .Z(net406));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer152 (.I(_06714_),
    .Z(net407));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer153 (.I(net407),
    .Z(net408));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 rebuffer154 (.I(_03928_),
    .Z(net409));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer155 (.I(_07732_),
    .Z(net410));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer156 (.I(_07817_),
    .Z(net411));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer157 (.I(_06683_),
    .Z(net412));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer158 (.I(net412),
    .Z(net413));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer159 (.I(_07641_),
    .Z(net414));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer160 (.I(net3606),
    .Z(net415));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 rebuffer161 (.I(net3606),
    .Z(net416));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer162 (.I(net449),
    .Z(net417));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer163 (.I(net3606),
    .Z(net418));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer164 (.I(_08055_),
    .Z(net419));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer165 (.I(_07346_),
    .Z(net420));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer166 (.I(_08543_),
    .Z(net421));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer167 (.I(_08543_),
    .Z(net422));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clone168 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .Z(net423));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer169 (.I(_07389_),
    .Z(net424));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer170 (.I(_06805_),
    .Z(net425));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer171 (.I(_06653_),
    .Z(net426));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer172 (.I(_06653_),
    .Z(net427));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer173 (.I(_08275_),
    .Z(net428));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer174 (.I(_08275_),
    .Z(net429));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer175 (.I(_08231_),
    .Z(net430));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer176 (.I(_08231_),
    .Z(net431));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer177 (.I(net431),
    .Z(net432));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer178 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .Z(net433));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone179 (.I(_03928_),
    .Z(net434));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer180 (.I(net3513),
    .Z(net435));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer181 (.I(_06487_),
    .Z(net436));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer182 (.I(net3280),
    .Z(net437));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer183 (.I(_07641_),
    .Z(net438));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer184 (.I(_07920_),
    .Z(net439));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer185 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .Z(net440));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer186 (.I(_07676_),
    .Z(net441));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer187 (.I(_07776_),
    .Z(net442));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer188 (.I(_07239_),
    .Z(net443));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone189 (.I(net3631),
    .Z(net444));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer190 (.I(_07566_),
    .Z(net445));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer191 (.I(net3272),
    .Z(net446));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer192 (.I(_08544_),
    .Z(net447));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer193 (.I(_06797_),
    .Z(net448));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clone194 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .Z(net449));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer195 (.I(_03925_),
    .Z(net450));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer196 (.I(_08507_),
    .Z(net451));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer197 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .Z(net452));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer198 (.I(net3633),
    .Z(net453));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer199 (.I(net3633),
    .Z(net454));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clone204 (.I(net335),
    .Z(net459));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer205 (.I(_03986_),
    .Z(net460));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 clone209 (.A1(net3190),
    .A2(net450),
    .B(_03927_),
    .ZN(net464));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone211 (.I(_03838_),
    .Z(net466));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone212 (.I(_03838_),
    .Z(net467));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer213 (.I(net276),
    .Z(net468));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer214 (.I(_07859_),
    .Z(net469));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer215 (.I(_07426_),
    .Z(net470));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer221 (.I(_10187_[0]),
    .Z(net476));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer222 (.I(net3115),
    .Z(net477));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer223 (.I(net3307),
    .Z(net478));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer224 (.I(net3276),
    .Z(net479));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone225 (.I(net3606),
    .Z(net480));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer226 (.I(net3307),
    .Z(net481));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer227 (.I(net3307),
    .Z(net482));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer228 (.I(_06511_),
    .Z(net483));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone273 (.I(net435),
    .Z(net528));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer274 (.I(_08496_),
    .Z(net529));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer275 (.I(_08110_),
    .Z(net530));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone292 (.I(net335),
    .Z(net547));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone300 (.I(_03956_),
    .Z(net555));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone301 (.I(_03956_),
    .Z(net556));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer302 (.I(_06457_),
    .Z(net557));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer303 (.I(net3516),
    .Z(net558));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer304 (.I(net3516),
    .Z(net559));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer320 (.I(net3541),
    .Z(net575));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer322 (.I(net3335),
    .Z(net577));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone323 (.I(net487),
    .Z(net578));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone324 (.I(net487),
    .Z(net579));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone325 (.I(_03813_),
    .Z(net580));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone451 (.I(_03760_),
    .Z(net737));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer329 (.I(_03813_),
    .Z(net584));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer330 (.I(_03748_),
    .Z(net585));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer370 (.I(_05008_),
    .Z(net625));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 clone372 (.A1(_03587_),
    .A2(_03571_),
    .ZN(net627));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer377 (.I(_07891_),
    .Z(net632));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer378 (.I(_04942_),
    .Z(net633));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold384 (.I(net640),
    .Z(net639));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold385 (.I(net642),
    .Z(net640));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold386 (.I(net639),
    .Z(net641));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold387 (.I(\core_clock_gate_i.en_latch ),
    .Z(net642));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 rebuffer12 (.I(net460),
    .Z(net335));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer27 (.I(_11097_[0]),
    .Z(net343));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer36 (.I(_06254_),
    .Z(net344));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 rebuffer50 (.I(_08065_),
    .Z(net345));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone80 (.I(net460),
    .Z(net385));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer88 (.I(_07304_),
    .Z(net388));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer89 (.I(_11025_[0]),
    .Z(net389));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer90 (.I(_06202_),
    .Z(net390));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer114 (.I(net3187),
    .Z(net393));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer115 (.I(net3187),
    .Z(net394));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer116 (.I(_08073_),
    .Z(net395));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer128 (.I(_08263_),
    .Z(net396));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer129 (.I(_05028_),
    .Z(net397));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer130 (.I(\id_stage_i.controller_i.instr_i[1] ),
    .Z(net398));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer133 (.I(_07395_),
    .Z(net399));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer134 (.I(_11029_[0]),
    .Z(net400));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer135 (.I(_11037_[0]),
    .Z(net401));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer138 (.I(_11037_[0]),
    .Z(net455));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer141 (.I(_09747_[0]),
    .Z(net458));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer142 (.I(_05018_),
    .Z(net461));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer143 (.I(_11101_[0]),
    .Z(net462));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer144 (.I(_11009_[0]),
    .Z(net463));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer145 (.I(_07002_),
    .Z(net465));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer146 (.I(_07002_),
    .Z(net471));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer168 (.I(_07008_),
    .Z(net472));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer179 (.I(_07008_),
    .Z(net473));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer189 (.I(_11014_[0]),
    .Z(net474));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer194 (.I(_07177_),
    .Z(net475));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer201 (.I(_06440_),
    .Z(net485));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 rebuffer202 (.I(_08154_),
    .Z(net486));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer203 (.I(_03860_),
    .Z(net487));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone452 (.I(_03760_),
    .Z(net738));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_2067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_72_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_2082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_2052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_1872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_2034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_103_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_103_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_103_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_103_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_103_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_103_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_104_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_104_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_104_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_104_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_104_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_104_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_104_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_105_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_105_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_105_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_105_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_105_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_105_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_106_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_106_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_106_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_106_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_106_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_106_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_106_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_107_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_107_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_107_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_107_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_107_2064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_107_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_107_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_108_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_108_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_108_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_108_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_108_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_108_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_108_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_109_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_109_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_109_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_109_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_109_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_109_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_110_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_110_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_110_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_110_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_110_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_110_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_111_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_111_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_111_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_111_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_111_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_111_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_112_1122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_112_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_112_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_112_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_112_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_112_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_112_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_113_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_113_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_113_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_113_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_113_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_113_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_114_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_114_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_114_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_114_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_114_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_114_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_115_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_115_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_115_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_115_2025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_115_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_115_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_115_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_116_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_116_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_116_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_116_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_116_2060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_116_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_116_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_117_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_117_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_117_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_117_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_117_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_117_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_118_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_118_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_118_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_118_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_118_2051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_118_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_118_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_119_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_119_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_119_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_119_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_119_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_119_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_119_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_120_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_120_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_120_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_120_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_120_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_2031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_120_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_120_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_121_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_121_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_121_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_121_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_121_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_121_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_121_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_122_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_122_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_122_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_122_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_122_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_122_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_122_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_123_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_123_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_123_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_123_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_123_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_123_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_123_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_124_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_124_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_124_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_124_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_124_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_124_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_124_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_125_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_125_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_125_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_125_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_125_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_125_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_125_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_126_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_126_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_126_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_126_2032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_126_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_126_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_127_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_127_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_127_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_127_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_127_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_127_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_127_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_128_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_128_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_128_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_128_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_128_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_128_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_128_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_129_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_129_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_129_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_129_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_129_2043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_129_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_129_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_130_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_130_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_130_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_130_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_130_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_130_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_131_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_131_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_131_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_131_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_131_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_131_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_132_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_132_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_132_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_132_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_132_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_132_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_133_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_133_2037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_133_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_133_2047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_133_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_134_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_134_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_134_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_134_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_134_2055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_134_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_135_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_135_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_135_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_135_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_135_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_135_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_135_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_136_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_136_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_136_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_136_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_136_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_136_2054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_136_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_137_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_137_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_137_1990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_137_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_137_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_137_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_137_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_138_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_138_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_138_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_138_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_138_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_138_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_139_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_139_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_139_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_139_2070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_139_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_139_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_139_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_140_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_140_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_140_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_140_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_140_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_140_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_140_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_141_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_141_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_141_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_141_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_141_2078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_141_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_141_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_142_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_142_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_142_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_142_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_142_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_142_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_142_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_143_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_143_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_143_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_143_2045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_143_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_143_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_143_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_144_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_1943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_144_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_144_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_144_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_144_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_144_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_144_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_145_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_145_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_145_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_145_2036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_145_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_145_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_146_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_146_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_146_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_146_2018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_146_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_146_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_146_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_147_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_147_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_147_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_147_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_147_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_147_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_147_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_148_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_148_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_148_1996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_148_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_148_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_148_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_148_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_149_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_149_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_149_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_149_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_149_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_149_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_149_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_150_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_150_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_150_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_150_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_150_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_150_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_150_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_1763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_151_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_151_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_151_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_151_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_151_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_151_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_151_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_152_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_152_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_152_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_152_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_152_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_152_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_152_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_153_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_153_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_153_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_153_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_153_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_153_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_153_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_154_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_154_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_154_1930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_154_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_154_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_154_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_154_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_155_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_155_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_155_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_1937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_155_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_155_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_155_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_155_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_156_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_156_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_156_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_156_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_156_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_156_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_156_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_157_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_157_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_157_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_157_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_157_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_157_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_157_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_158_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_158_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_158_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_158_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_158_2076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_158_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_158_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_159_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_159_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_159_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_159_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_159_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_159_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_159_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_160_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_160_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_160_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_160_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_160_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_160_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_160_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_161_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_161_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_161_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_161_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_161_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_161_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_161_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1043 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_162_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_162_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_162_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_162_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_162_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_162_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_162_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_163_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_163_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_163_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_163_2028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_163_2092 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_163_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_163_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_164_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_164_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_164_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_164_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_164_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_164_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_164_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1032 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_165_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_165_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_165_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_165_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_165_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_165_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_165_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_166_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_166_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_166_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_166_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_166_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_166_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_166_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_167_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_167_2057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_167_2089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_167_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_167_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_167_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_167_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1036 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_168_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_168_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_168_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_168_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_168_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_168_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1052 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_169_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_169_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_169_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_169_2042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_169_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_169_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_169_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_1785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_170_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_170_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_170_2058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_170_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_170_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_170_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_170_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_171_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_171_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_171_1959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_171_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_171_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_171_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_171_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_172_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_172_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_172_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_172_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_172_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_172_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_172_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_173_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_173_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_173_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_173_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_173_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_173_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_173_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_174_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_174_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_174_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_174_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_174_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_174_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_175_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_175_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_175_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_175_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_175_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_175_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_175_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_176_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_176_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_176_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_176_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_176_2016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_176_2080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_176_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_177_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_1926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_177_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_177_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_177_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_177_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_177_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_177_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_361 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_178_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_178_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_1981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_178_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_178_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_178_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_178_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_178_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_179_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_179_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_1841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_179_1888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_179_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_179_2050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_179_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_179_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_180_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_180_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_180_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_180_1975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_180_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_180_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_180_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1034 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_181_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_1986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_181_1997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_181_2061 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_181_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_181_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_181_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_181_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_182_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_182_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_182_1993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_182_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_182_2068 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_182_2100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_182_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_183_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_183_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_1904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_183_2017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_183_2081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_183_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_183_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_183_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_184_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_184_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_184_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_184_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_184_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_184_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_184_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1082 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_185_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_185_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_185_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_185_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_185_2022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_185_2086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_185_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_981 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_1796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_186_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_186_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_186_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_186_2015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_186_2079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_186_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_186_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_187_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_187_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_187_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_187_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_187_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_187_2040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_187_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_188_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_188_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_188_1998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_188_2062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_188_2094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_188_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_188_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_189_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_189_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_189_2029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_189_2093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_189_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_189_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_189_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_190_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_190_1914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_1922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_190_1976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_190_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_190_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_190_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_190_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_191_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_191_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_191_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_191_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_191_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_191_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_191_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_1575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_192_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_192_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_192_2004 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_2014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_192_2021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_192_2085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_192_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_192_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_193_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_193_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_193_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_193_2075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_193_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_193_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_193_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_194_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_194_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1970 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_194_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_194_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_194_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_194_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_194_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1045 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_195_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_1804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_195_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_195_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_195_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_195_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_195_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_195_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_196_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_196_2001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_196_2065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_196_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_196_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_196_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_196_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_197_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_197_1963 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_197_1979 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_197_1987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_197_2023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_197_2087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_197_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_993 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_198_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_198_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_1964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_198_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_198_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_198_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_198_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_198_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_199_1704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_199_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_199_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_199_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_1919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_1989 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_199_2053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_199_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_199_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_200_1855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_1978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_200_2003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_200_2011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_200_2019 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_200_2083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_200_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_200_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1085 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1093 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_201_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_201_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_201_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_201_1932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_201_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_201_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_1992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_201_2056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_1489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_202_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_202_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_202_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_202_2046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_202_2110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_202_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_203_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_203_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_203_1945 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_203_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_1982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_203_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_203_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_203_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_204_1518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_204_1780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_204_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_1892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_204_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_2006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_204_2020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_204_2084 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_204_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_1569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_205_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_205_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_205_1953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_205_1967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_205_1988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_205_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_205_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_987 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1042 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_206_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_206_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_1994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_206_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_206_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_206_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_206_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_206_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_940 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1031 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_207_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_207_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_207_1900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_1985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_207_2049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_207_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_207_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_207_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1081 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_208_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_1915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_208_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_208_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_208_2063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_208_2095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_208_2111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_208_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_978 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1016 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_1973 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_209_1983 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_209_1991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_209_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_209_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_209_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_209_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_209_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1021 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_1257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_210_1535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_1702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_1968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_1972 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_210_2009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_210_2073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_210_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_210_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_210_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_210_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_1271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_1402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_1710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_211_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_1911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_211_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_211_2013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_211_2077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_211_2109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_211_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_211_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_953 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1017 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1049 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1080 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1096 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_212_1887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_212_1935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_212_1949 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_1951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_2000 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_212_2007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_212_2071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_212_2103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_212_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1011 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_1456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_213_1807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_1933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_213_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_1999 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_213_2010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_213_2074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_213_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_213_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_213_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_943 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_986 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_996 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1076 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1078 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_1210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_1301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_1407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_1432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_214_1711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_1802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_214_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_1936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_1952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_214_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_214_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_1980 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_214_2044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_214_2108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_214_2116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_215_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_997 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1003 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_1485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_1548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_1699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_215_1798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_215_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_1917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_1921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_1971 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_215_2035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_215_2099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_215_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_215_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1075 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1077 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_216_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_1299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_216_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_1891 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_1966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_1977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_216_2041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_216_2105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_216_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_216_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_216_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_965 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_967 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_998 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1054 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1062 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1074 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_1342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_1840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_217_1876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_1890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_1912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_217_1958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_217_2002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_217_2066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_217_2098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_217_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_217_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_1002 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1030 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1056 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_1475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_1515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_218_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_218_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_218_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_218_1889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_1925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_218_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_218_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_218_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_959 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1039 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1041 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_1400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_1673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_1705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_1767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_219_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_1847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_219_1863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_219_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_219_1934 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_219_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_219_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_219_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_936 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_966 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_975 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1094 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_220_1858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_220_1882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_220_1902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_220_1946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_220_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_220_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_220_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_873 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_964 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1037 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_1047 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1063 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_1231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_1406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_221_1731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_221_1861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_1865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_221_2005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_221_2069 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_221_2101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_221_2117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_221_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1025 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1035 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1053 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1071 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_1129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_1621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_222_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_222_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_222_1947 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_222_1955 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_222_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_222_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_222_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_991 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_1104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_1416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_1529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_1572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_223_1693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_223_1811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_223_1843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_1895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_1969 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_223_2033 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_223_2097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_223_2113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_223_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1010 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1073 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_1089 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_224_1662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_224_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_224_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_224_1907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_1918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_224_1950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_224_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_224_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_914 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_992 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1046 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1050 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1095 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_225_1597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_225_1836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_1852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_225_1864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_225_1874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_225_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_1984 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_225_2048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_225_2112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_951 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1005 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1007 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1051 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1055 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1057 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_226_1885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_226_1893 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_226_1897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_1909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_226_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_226_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_226_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_226_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_968 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_985 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_1001 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1009 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1013 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_1079 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1087 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_1230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_227_1304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_1774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_1778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_227_1790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_1962 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_227_2026 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_227_2090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_227_2106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_227_2114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_227_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_939 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1014 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1018 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1020 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_1083 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_1099 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_1238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_1280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_1497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_1636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_1691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_228_1707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_228_1801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_228_1832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_1906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_228_1938 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_228_1954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_228_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_228_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_976 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1065 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1067 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_1086 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_1227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_1533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_1696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_1721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_1753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_1795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_229_1803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_1853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_1857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_229_1995 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_229_2059 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_229_2091 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_229_2107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_229_2115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_229_2119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_988 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_1006 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1022 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1097 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_1105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_1148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_1248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_1324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_1437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_1561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_1618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_230_1658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_230_1674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_1684 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_230_1792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_230_1948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_230_1956 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_230_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_230_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_946 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_950 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_952 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_1015 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_1023 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1027 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1029 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_1142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_1150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_1337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_1452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_231_1536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_1645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_1713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_231_1773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_231_1777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_231_1779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_1944 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_231_2008 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_231_2072 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_231_2104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_954 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_958 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_982 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_990 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_1024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_1040 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_1048 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_1090 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1098 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_1241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_232_1336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_1344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_1473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_1562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_1638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_232_1651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_232_1771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_232_1941 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_232_1957 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_232_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_232_2088 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_935 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_937 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_961 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_977 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_994 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_1058 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1066 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_1102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_1110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_1124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_233_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_233_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_1609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_1625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_1635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_1692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_1708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_233_1715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_1725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_1748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_233_1762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_1974 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_233_2038 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_233_2102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_233_2118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_948 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1012 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_1044 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_1060 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1070 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_1168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_1192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_1206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_1214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_1218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_1245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_1258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_1274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_1278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_1334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_234_1350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_1368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_234_1384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_234_1390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_234_1422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_1586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_1764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_1910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_234_1942 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_1960 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_234_2024 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_234_2088 ();
 assign alert_major_o = net250;
endmodule
